* NGSPICE file created from sky130_fd_sc_hd__a2bb2o_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__a2bb2o_1 VGND VPWR B1 A1_N A2_N X B2 VNB VPB
X0 a_226_47.t0 A2_N.t0 a_226_297.t0 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1 a_489_413.t0 B1.t0 VPWR.t1 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 a_226_297.t1 A1_N.t0 VPWR.t3 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3 VPWR.t2 B2.t0 a_489_413.t1 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 a_489_413.t2 a_226_47.t3 a_76_199.t2 VPB.t5 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 a_76_199.t1 a_226_47.t4 VGND.t4 VNB.t5 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 VGND.t1 B1.t1 a_556_47.t0 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7 a_556_47.t1 B2.t1 a_76_199.t0 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 VGND.t0 A2_N.t1 a_226_47.t1 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9 a_226_47.t2 A1_N.t1 VGND.t2 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10 VPWR.t0 a_76_199.t3 X.t0 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 VGND.t3 a_76_199.t4 X.t1 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
R0 A2_N.n0 A2_N.t1 206.188
R1 A2_N.n0 A2_N.t0 142.34
R2 A2_N A2_N.n0 78.427
R3 a_226_297.t0 a_226_297.t1 98.5
R4 a_226_47.t0 a_226_47.n2 417.937
R5 a_226_47.n0 a_226_47.t3 286.316
R6 a_226_47.n2 a_226_47.n1 180.216
R7 a_226_47.n0 a_226_47.t4 131.097
R8 a_226_47.n2 a_226_47.n0 76
R9 a_226_47.n1 a_226_47.t1 38.571
R10 a_226_47.n1 a_226_47.t2 38.571
R11 VPB.t2 VPB.t5 565.264
R12 VPB.t1 VPB.t4 346.261
R13 VPB.t3 VPB.t0 248.598
R14 VPB.t5 VPB.t3 248.598
R15 VPB.t4 VPB.t2 213.084
R16 VPB VPB.t1 189.408
R17 B1.n0 B1.t0 327.055
R18 B1.n0 B1.t1 239.766
R19 B1.n1 B1.n0 76
R20 B1.n1 B1 14.03
R21 B1 B1.n1 2.707
R22 VPWR.n2 VPWR.n1 316.665
R23 VPWR.n2 VPWR.n0 312.522
R24 VPWR.n0 VPWR.t3 143.059
R25 VPWR.n1 VPWR.t1 63.321
R26 VPWR.n1 VPWR.t2 63.321
R27 VPWR.n0 VPWR.t0 25.61
R28 VPWR VPWR.n2 9.426
R29 a_489_413.t0 a_489_413.n0 746.507
R30 a_489_413.n0 a_489_413.t1 63.321
R31 a_489_413.n0 a_489_413.t2 63.321
R32 A1_N.n0 A1_N.t1 206.188
R33 A1_N.n0 A1_N.t0 148.348
R34 A1_N.n1 A1_N.n0 76
R35 A1_N.n1 A1_N 11.054
R36 A1_N A1_N.n1 2.133
R37 B2.n0 B2.t1 305.801
R38 B2.n0 B2.t0 235.108
R39 B2 B2.n0 82.186
R40 a_76_199.n1 a_76_199.t2 355.821
R41 a_76_199.n1 a_76_199.n0 242.523
R42 a_76_199.n0 a_76_199.t3 241.534
R43 a_76_199.n2 a_76_199.n1 228.027
R44 a_76_199.n0 a_76_199.t4 169.234
R45 a_76_199.t0 a_76_199.n2 38.571
R46 a_76_199.n2 a_76_199.t1 38.571
R47 VGND.n2 VGND.t1 148.528
R48 VGND.n1 VGND.n0 105.746
R49 VGND.n4 VGND.n3 92.5
R50 VGND.n8 VGND.n7 92.5
R51 VGND.n0 VGND.t2 85.714
R52 VGND.n3 VGND.t4 38.571
R53 VGND.n7 VGND.t0 38.571
R54 VGND.n0 VGND.t3 25.934
R55 VGND VGND.n13 9.338
R56 VGND.n6 VGND.n5 4.65
R57 VGND.n10 VGND.n9 4.65
R58 VGND.n12 VGND.n11 4.65
R59 VGND.n13 VGND.n1 3.232
R60 VGND.n9 VGND.n8 1.684
R61 VGND.n13 VGND.n12 0.838
R62 VGND.n6 VGND.n2 0.242
R63 VGND.n10 VGND.n6 0.119
R64 VGND.n12 VGND.n10 0.119
R65 VGND.n5 VGND.n4 0.112
R66 VNB VNB.t4 6053.91
R67 VNB.t0 VNB.t5 5241.18
R68 VNB.t4 VNB.t2 3041.18
R69 VNB.t3 VNB.t1 2717.65
R70 VNB.t5 VNB.t3 2717.65
R71 VNB.t2 VNB.t0 2717.65
R72 a_556_47.t0 a_556_47.t1 77.142
R73 X.t0 X 463.13
R74 X.n1 X.t0 462.98
R75 X.n0 X.t1 117.423
R76 X.n1 X.n0 76.173
R77 X.n0 X 6.646
R78 X X.n1 1.23
C0 B2 B1 0.20fF
C1 A1_N A2_N 0.14fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__a2bb2o_2.ext - technology: sky130A

.subckt sky130_fd_sc_hd__a2bb2o_2 VGND VPWR B1 A1_N A2_N X B2 VNB VPB
X0 VPWR.t1 a_82_21.t3 X.t3 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_646_47.t0 B2.t0 a_82_21.t2 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 a_574_369.t2 a_313_47.t3 a_82_21.t0 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X3 a_574_369.t1 B1.t0 VPWR.t3 VPB.t5 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X4 VGND.t1 a_82_21.t4 X.t1 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 VPWR.t4 B2.t1 a_574_369.t0 VPB.t6 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X6 X.t0 a_82_21.t5 VGND.t0 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 X.t2 a_82_21.t6 VPWR.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 a_313_47.t1 A2_N.t0 a_313_297.t1 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X9 a_313_47.t0 A1_N.t0 VGND.t2 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10 a_313_297.t0 A1_N.t1 VPWR.t2 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X11 VGND.t3 A2_N.t1 a_313_47.t2 VNB.t6 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12 a_82_21.t1 a_313_47.t4 VGND.t5 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13 VGND.t4 B1.t1 a_646_47.t1 VNB.t5 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
R0 a_82_21.t0 a_82_21.n3 334.054
R1 a_82_21.n3 a_82_21.n1 250.279
R2 a_82_21.n3 a_82_21.n2 225.997
R3 a_82_21.n1 a_82_21.t3 212.079
R4 a_82_21.n0 a_82_21.t6 212.079
R5 a_82_21.n1 a_82_21.t4 139.779
R6 a_82_21.n0 a_82_21.t5 139.779
R7 a_82_21.n1 a_82_21.n0 61.345
R8 a_82_21.n2 a_82_21.t2 38.571
R9 a_82_21.n2 a_82_21.t1 38.571
R10 X.n0 X 296.515
R11 X.n3 X.n0 292.5
R12 X.n2 X.n1 92.5
R13 X.n3 X.n2 78.18
R14 X.n0 X.t3 26.595
R15 X.n0 X.t2 26.595
R16 X.n1 X.t1 24.923
R17 X.n1 X.t0 24.923
R18 X.n2 X 6.776
R19 X X.n3 1.254
R20 VPWR.n3 VPWR.n2 455.765
R21 VPWR.n4 VPWR.n1 316.039
R22 VPWR.n0 VPWR.t0 161.95
R23 VPWR.n2 VPWR.t2 93.882
R24 VPWR.n1 VPWR.t3 41.554
R25 VPWR.n1 VPWR.t4 41.554
R26 VPWR.n2 VPWR.t1 29.055
R27 VPWR VPWR.n7 7.905
R28 VPWR.n7 VPWR.n6 4.769
R29 VPWR.n6 VPWR.n5 4.65
R30 VPWR.n4 VPWR.n3 3.992
R31 VPWR.n7 VPWR.n0 3.011
R32 VPWR.n6 VPWR.n4 0.138
R33 VPB.t3 VPB.t2 559.345
R34 VPB.t1 VPB.t4 346.261
R35 VPB.t2 VPB.t6 269.314
R36 VPB.t6 VPB.t5 248.598
R37 VPB.t0 VPB.t1 248.598
R38 VPB.t4 VPB.t3 213.084
R39 VPB VPB.t0 213.084
R40 B2.n0 B2.t0 305.801
R41 B2.n0 B2.t1 199.761
R42 B2 B2.n0 82.186
R43 a_646_47.t0 a_646_47.t1 77.142
R44 VNB VNB.t0 6247.32
R45 VNB.t6 VNB.t4 5338.23
R46 VNB.t1 VNB.t2 3041.18
R47 VNB.t3 VNB.t5 2717.65
R48 VNB.t4 VNB.t3 2717.65
R49 VNB.t2 VNB.t6 2717.65
R50 VNB.t0 VNB.t1 2030.77
R51 a_313_47.t1 a_313_47.n2 390.9
R52 a_313_47.n0 a_313_47.t3 257.84
R53 a_313_47.n2 a_313_47.n1 187.746
R54 a_313_47.n0 a_313_47.t4 138.016
R55 a_313_47.n2 a_313_47.n0 76
R56 a_313_47.n1 a_313_47.t2 38.571
R57 a_313_47.n1 a_313_47.t0 38.571
R58 a_574_369.n0 a_574_369.t1 726.225
R59 a_574_369.n0 a_574_369.t2 52.328
R60 a_574_369.t0 a_574_369.n0 41.554
R61 B1.n0 B1.t0 292.321
R62 B1.n0 B1.t1 241.429
R63 B1.n1 B1.n0 76
R64 B1.n1 B1 14.03
R65 B1 B1.n1 2.707
R66 VGND.n3 VGND.t4 148.697
R67 VGND.n0 VGND.t0 113.165
R68 VGND.n11 VGND.n10 105.746
R69 VGND.n2 VGND.n1 92.5
R70 VGND.n5 VGND.n4 92.5
R71 VGND.n10 VGND.t2 85.714
R72 VGND.n1 VGND.t5 38.571
R73 VGND.n4 VGND.t3 38.571
R74 VGND.n10 VGND.t1 25.934
R75 VGND VGND.n15 7.905
R76 VGND.n15 VGND.n14 4.769
R77 VGND.n7 VGND.n6 4.65
R78 VGND.n9 VGND.n8 4.65
R79 VGND.n12 VGND.n11 4.65
R80 VGND.n14 VGND.n13 4.65
R81 VGND.n3 VGND.n2 4.114
R82 VGND.n15 VGND.n0 3.011
R83 VGND.n6 VGND.n5 1.122
R84 VGND.n7 VGND.n3 0.152
R85 VGND.n9 VGND.n7 0.119
R86 VGND.n12 VGND.n9 0.119
R87 VGND.n14 VGND.n12 0.119
R88 A2_N.n0 A2_N.t1 206.188
R89 A2_N.n0 A2_N.t0 177.686
R90 A2_N A2_N.n0 78.427
R91 a_313_297.t0 a_313_297.t1 64.64
R92 A1_N.n0 A1_N.t0 206.188
R93 A1_N.n0 A1_N.t1 183.694
R94 A1_N.n1 A1_N.n0 76
R95 A1_N.n1 A1_N 11.054
R96 A1_N A1_N.n1 2.133
C0 X VGND 0.18fF
C1 B2 B1 0.19fF
C2 A1_N A2_N 0.14fF
C3 VGND VPWR 0.11fF
C4 X VPWR 0.20fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__a2bb2o_4.ext - technology: sky130A

.subckt sky130_fd_sc_hd__a2bb2o_4 B1 B2 X A1_N A2_N VGND VPWR VNB VPB
X0 VGND.t1 a_415_21.t6 a_193_47.t2 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 a_415_21.t0 A2_N.t0 a_717_297.t1 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 a_717_297.t2 A1_N.t0 VPWR.t8 VPB.t8 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 VGND.t6 A2_N.t1 a_415_21.t1 VNB.t7 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 a_193_47.t3 a_415_21.t7 a_27_297.t1 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 a_27_297.t5 B1.t0 VPWR.t9 VPB.t13 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 VPWR.t3 a_193_47.t6 X.t7 VPB.t7 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 X.t3 a_193_47.t7 VGND.t3 VNB.t6 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 VPWR.t4 B2.t0 a_27_297.t2 VPB.t10 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 X.t6 a_193_47.t8 VPWR.t2 VPB.t6 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 a_415_21.t4 A1_N.t1 VGND.t8 VNB.t9 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 a_415_21.t2 A2_N.t2 VGND.t7 VNB.t8 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 X.t2 a_193_47.t9 VGND.t2 VNB.t5 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 a_27_297.t3 B2.t1 VPWR.t5 VPB.t11 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14 a_193_47.t5 B2.t2 a_109_47.t1 VNB.t11 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X15 VGND.t10 B1.t1 a_109_47.t3 VNB.t12 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X16 VGND.t5 a_193_47.t10 X.t1 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X17 VGND.t9 A1_N.t2 a_415_21.t5 VNB.t10 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X18 VGND.t4 a_193_47.t11 X.t0 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X19 a_109_47.t0 B2.t3 a_193_47.t4 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X20 a_193_47.t1 a_415_21.t8 VGND.t0 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X21 VPWR.t1 a_193_47.t12 X.t5 VPB.t5 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X22 a_27_297.t0 a_415_21.t9 a_193_47.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X23 X.t4 a_193_47.t13 VPWR.t0 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X24 VPWR.t7 A1_N.t3 a_717_297.t3 VPB.t9 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X25 VPWR.t6 B1.t2 a_27_297.t4 VPB.t12 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X26 a_717_297.t0 A2_N.t3 a_415_21.t3 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X27 a_109_47.t2 B1.t3 VGND.t11 VNB.t13 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
R0 a_415_21.n6 a_415_21.n5 398.141
R1 a_415_21.n1 a_415_21.t9 212.079
R2 a_415_21.n0 a_415_21.t7 212.079
R3 a_415_21.n1 a_415_21.t6 139.779
R4 a_415_21.n0 a_415_21.t8 139.779
R5 a_415_21.n5 a_415_21.n1 119.848
R6 a_415_21.n4 a_415_21.n2 88.89
R7 a_415_21.n1 a_415_21.n0 61.345
R8 a_415_21.n4 a_415_21.n3 52.624
R9 a_415_21.n5 a_415_21.n4 52.397
R10 a_415_21.n6 a_415_21.t3 26.595
R11 a_415_21.t0 a_415_21.n6 26.595
R12 a_415_21.n2 a_415_21.t5 24.923
R13 a_415_21.n2 a_415_21.t2 24.923
R14 a_415_21.n3 a_415_21.t1 24.923
R15 a_415_21.n3 a_415_21.t4 24.923
R16 a_193_47.n0 a_193_47.t6 212.079
R17 a_193_47.n2 a_193_47.t8 212.079
R18 a_193_47.n5 a_193_47.t12 212.079
R19 a_193_47.n6 a_193_47.t13 212.079
R20 a_193_47.n11 a_193_47.n9 170.516
R21 a_193_47.n13 a_193_47.n12 152.016
R22 a_193_47.n0 a_193_47.t11 139.779
R23 a_193_47.n2 a_193_47.t9 139.779
R24 a_193_47.n5 a_193_47.t10 139.779
R25 a_193_47.n6 a_193_47.t7 139.779
R26 a_193_47.n4 a_193_47.n1 101.6
R27 a_193_47.n4 a_193_47.n3 76
R28 a_193_47.n8 a_193_47.n7 76
R29 a_193_47.n11 a_193_47.n10 52.818
R30 a_193_47.n7 a_193_47.n6 49.66
R31 a_193_47.n12 a_193_47.n11 38.204
R32 a_193_47.n1 a_193_47.n0 35.054
R33 a_193_47.n12 a_193_47.n8 31.521
R34 a_193_47.t0 a_193_47.n13 26.595
R35 a_193_47.n13 a_193_47.t3 26.595
R36 a_193_47.n8 a_193_47.n4 25.6
R37 a_193_47.n10 a_193_47.t2 24.923
R38 a_193_47.n10 a_193_47.t1 24.923
R39 a_193_47.n9 a_193_47.t4 24.923
R40 a_193_47.n9 a_193_47.t5 24.923
R41 a_193_47.n3 a_193_47.n2 23.369
R42 a_193_47.n7 a_193_47.n5 11.684
R43 VGND.n0 VGND.t4 197.839
R44 VGND.n2 VGND.n1 115.464
R45 VGND.n14 VGND.n13 115.464
R46 VGND.n28 VGND.n27 115.464
R47 VGND.n37 VGND.t11 114.4
R48 VGND.n20 VGND.n19 92.5
R49 VGND.n22 VGND.n21 92.5
R50 VGND.n8 VGND.n7 74.837
R51 VGND.n19 VGND.t8 24.923
R52 VGND.n21 VGND.t1 24.923
R53 VGND.n1 VGND.t2 24.923
R54 VGND.n1 VGND.t5 24.923
R55 VGND.n7 VGND.t3 24.923
R56 VGND.n7 VGND.t9 24.923
R57 VGND.n13 VGND.t7 24.923
R58 VGND.n13 VGND.t6 24.923
R59 VGND.n27 VGND.t0 24.923
R60 VGND.n27 VGND.t10 24.923
R61 VGND.n15 VGND.n14 17.317
R62 VGND.n9 VGND.n8 11.294
R63 VGND.n29 VGND.n28 9.788
R64 VGND.n38 VGND.n37 6.908
R65 VGND.n23 VGND.n20 6.2
R66 VGND.n3 VGND.n2 5.27
R67 VGND.n4 VGND.n3 4.65
R68 VGND.n6 VGND.n5 4.65
R69 VGND.n10 VGND.n9 4.65
R70 VGND.n12 VGND.n11 4.65
R71 VGND.n16 VGND.n15 4.65
R72 VGND.n18 VGND.n17 4.65
R73 VGND.n24 VGND.n23 4.65
R74 VGND.n26 VGND.n25 4.65
R75 VGND.n30 VGND.n29 4.65
R76 VGND.n32 VGND.n31 4.65
R77 VGND.n34 VGND.n33 4.65
R78 VGND.n36 VGND.n35 4.65
R79 VGND.n23 VGND.n22 4.2
R80 VGND.n4 VGND.n0 0.657
R81 VGND.n6 VGND.n4 0.119
R82 VGND.n10 VGND.n6 0.119
R83 VGND.n12 VGND.n10 0.119
R84 VGND.n16 VGND.n12 0.119
R85 VGND.n18 VGND.n16 0.119
R86 VGND.n24 VGND.n18 0.119
R87 VGND.n26 VGND.n24 0.119
R88 VGND.n30 VGND.n26 0.119
R89 VGND.n32 VGND.n30 0.119
R90 VGND.n34 VGND.n32 0.119
R91 VGND.n36 VGND.n34 0.119
R92 VGND.n38 VGND.n36 0.119
R93 VGND VGND.n38 0.02
R94 VNB VNB.t13 6053.91
R95 VNB.t1 VNB.t9 4545.05
R96 VNB.t5 VNB.t3 2030.77
R97 VNB.t4 VNB.t5 2030.77
R98 VNB.t6 VNB.t4 2030.77
R99 VNB.t10 VNB.t6 2030.77
R100 VNB.t8 VNB.t10 2030.77
R101 VNB.t7 VNB.t8 2030.77
R102 VNB.t9 VNB.t7 2030.77
R103 VNB.t0 VNB.t1 2030.77
R104 VNB.t12 VNB.t0 2030.77
R105 VNB.t2 VNB.t12 2030.77
R106 VNB.t11 VNB.t2 2030.77
R107 VNB.t13 VNB.t11 2030.77
R108 A2_N.n0 A2_N.t3 212.079
R109 A2_N.n1 A2_N.t0 212.079
R110 A2_N.n0 A2_N.t2 139.779
R111 A2_N.n1 A2_N.t1 139.779
R112 A2_N A2_N.n2 94.88
R113 A2_N.n2 A2_N.n1 31.403
R114 A2_N.n2 A2_N.n0 29.942
R115 a_717_297.n1 a_717_297.n0 496.344
R116 a_717_297.n0 a_717_297.t3 26.595
R117 a_717_297.n0 a_717_297.t0 26.595
R118 a_717_297.t1 a_717_297.n1 26.595
R119 a_717_297.n1 a_717_297.t2 26.595
R120 VPB.t0 VPB.t8 556.386
R121 VPB.t6 VPB.t7 248.598
R122 VPB.t5 VPB.t6 248.598
R123 VPB.t4 VPB.t5 248.598
R124 VPB.t9 VPB.t4 248.598
R125 VPB.t2 VPB.t9 248.598
R126 VPB.t3 VPB.t2 248.598
R127 VPB.t8 VPB.t3 248.598
R128 VPB.t1 VPB.t0 248.598
R129 VPB.t13 VPB.t1 248.598
R130 VPB.t10 VPB.t13 248.598
R131 VPB.t11 VPB.t10 248.598
R132 VPB.t12 VPB.t11 248.598
R133 VPB VPB.t12 189.408
R134 A1_N.n0 A1_N.t3 241.534
R135 A1_N.n2 A1_N.t0 236.179
R136 A1_N.n0 A1_N.t2 169.234
R137 A1_N.n2 A1_N.t1 163.879
R138 A1_N.n3 A1_N.n1 107.272
R139 A1_N.n3 A1_N.n2 76
R140 A1_N.n1 A1_N.n0 76
R141  A1_N.n3 2.133
R142 A1_N.n1 A1_N 1.955
R143 VPWR.n13 VPWR.t8 580.936
R144 VPWR.n23 VPWR.n22 314.004
R145 VPWR.n28 VPWR.n27 314.004
R146 VPWR.n1 VPWR.n0 312.468
R147 VPWR.n2 VPWR.t3 200.67
R148 VPWR.n6 VPWR.n5 171.981
R149 VPWR.n0 VPWR.t2 26.595
R150 VPWR.n0 VPWR.t1 26.595
R151 VPWR.n5 VPWR.t0 26.595
R152 VPWR.n5 VPWR.t7 26.595
R153 VPWR.n22 VPWR.t9 26.595
R154 VPWR.n22 VPWR.t4 26.595
R155 VPWR.n27 VPWR.t5 26.595
R156 VPWR.n27 VPWR.t6 26.595
R157 VPWR.n4 VPWR.n3 4.65
R158 VPWR.n8 VPWR.n7 4.65
R159 VPWR.n10 VPWR.n9 4.65
R160 VPWR.n12 VPWR.n11 4.65
R161 VPWR.n15 VPWR.n14 4.65
R162 VPWR.n17 VPWR.n16 4.65
R163 VPWR.n19 VPWR.n18 4.65
R164 VPWR.n21 VPWR.n20 4.65
R165 VPWR.n24 VPWR.n23 4.65
R166 VPWR.n26 VPWR.n25 4.65
R167 VPWR.n29 VPWR.n28 3.996
R168 VPWR.n2 VPWR.n1 3.784
R169 VPWR.n7 VPWR.n6 1.882
R170 VPWR.n14 VPWR.n13 1.882
R171 VPWR.n4 VPWR.n2 0.233
R172 VPWR.n29 VPWR.n26 0.136
R173 VPWR VPWR.n29 0.123
R174 VPWR.n8 VPWR.n4 0.119
R175 VPWR.n10 VPWR.n8 0.119
R176 VPWR.n12 VPWR.n10 0.119
R177 VPWR.n15 VPWR.n12 0.119
R178 VPWR.n17 VPWR.n15 0.119
R179 VPWR.n19 VPWR.n17 0.119
R180 VPWR.n21 VPWR.n19 0.119
R181 VPWR.n24 VPWR.n21 0.119
R182 VPWR.n26 VPWR.n24 0.119
R183 a_27_297.n2 a_27_297.t0 597.009
R184 a_27_297.n1 a_27_297.t4 226.103
R185 a_27_297.n1 a_27_297.n0 155.085
R186 a_27_297.n3 a_27_297.n2 94.349
R187 a_27_297.n2 a_27_297.n1 53.101
R188 a_27_297.n0 a_27_297.t2 26.595
R189 a_27_297.n0 a_27_297.t3 26.595
R190 a_27_297.t1 a_27_297.n3 26.595
R191 a_27_297.n3 a_27_297.t5 26.595
R192 B1.n1 B1.t2 241.534
R193 B1.n0 B1.t0 241.534
R194 B1.n2 B1.n0 181.933
R195 B1.n1 B1.t3 169.234
R196 B1.n0 B1.t1 169.234
R197 B1.n2 B1.n1 76
R198 B1 B1.n2 6.162
R199 X.n2 X.n0 203.821
R200 X.n2 X.n1 98.532
R201 X.n5 X.n3 88.89
R202 X.n5 X.n4 52.624
R203 X X.n2 29.267
R204 X.n1 X.t7 26.595
R205 X.n1 X.t6 26.595
R206 X.n0 X.t5 26.595
R207 X.n0 X.t4 26.595
R208  X.n5 26.551
R209 X.n3 X.t1 24.923
R210 X.n3 X.t3 24.923
R211 X.n4 X.t0 24.923
R212 X.n4 X.t2 24.923
R213  X 14.038
R214 B2.n0 B2.t0 212.079
R215 B2.n1 B2.t1 212.079
R216 B2.n0 B2.t3 139.779
R217 B2.n1 B2.t2 139.779
R218 B2 B2.n2 77.303
R219 B2.n2 B2.n0 30.672
R220 B2.n2 B2.n1 30.672
R221 a_109_47.n1 a_109_47.n0 187.937
R222 a_109_47.n0 a_109_47.t3 24.923
R223 a_109_47.n0 a_109_47.t0 24.923
R224 a_109_47.t1 a_109_47.n1 24.923
R225 a_109_47.n1 a_109_47.t2 24.923
C0 VPWR VPB 0.15fF
C1 VPWR X 0.52fF
C2 A1_N A2_N 0.35fF
C3 X VGND 0.47fF
C4 B1 B2 0.31fF
C5 VPWR VGND 0.12fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__a2bb2oi_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__a2bb2oi_1 A1_N Y VGND VPWR B2 B1 A2_N VNB VPB
X0 a_109_47.t2 A2_N.t0 a_109_297.t1 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_397_297.t0 B1.t0 VPWR.t1 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 VPWR.t2 B2.t0 a_397_297.t1 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 VGND.t2 A2_N.t1 a_109_47.t1 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 a_397_297.t2 a_109_47.t3 Y.t0 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 a_481_47.t1 B2.t1 Y.t2 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 Y.t1 a_109_47.t4 VGND.t3 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 VGND.t1 B1.t1 a_481_47.t0 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 a_109_297.t0 A1_N.t0 VPWR.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 a_109_47.t0 A1_N.t1 VGND.t0 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
R0 A2_N.n0 A2_N.t0 241.534
R1 A2_N.n0 A2_N.t1 169.234
R2 A2_N A2_N.n0 84.694
R3 a_109_297.t0 a_109_297.t1 41.37
R4 a_109_47.n0 a_109_47.t3 212.079
R5 a_109_47.n2 a_109_47.n1 186.24
R6 a_109_47.t2 a_109_47.n2 178.687
R7 a_109_47.n0 a_109_47.t4 139.779
R8 a_109_47.n2 a_109_47.n0 136.615
R9 a_109_47.n1 a_109_47.t1 24.923
R10 a_109_47.n1 a_109_47.t0 24.923
R11 VPB.t1 VPB.t3 639.252
R12 VPB.t2 VPB.t4 248.598
R13 VPB.t3 VPB.t2 248.598
R14 VPB.t0 VPB.t1 213.084
R15 VPB VPB.t0 192.367
R16 B1.n0 B1.t0 236.549
R17 B1.n0 B1.t1 164.249
R18 B1 B1.n0 78.427
R19 VPWR.n1 VPWR.n0 315.012
R20 VPWR.n1 VPWR.t0 195.077
R21 VPWR.n0 VPWR.t1 26.595
R22 VPWR.n0 VPWR.t2 26.595
R23 VPWR VPWR.n1 0.044
R24 a_397_297.t0 a_397_297.n0 545.75
R25 a_397_297.n0 a_397_297.t1 26.595
R26 a_397_297.n0 a_397_297.t2 26.595
R27 B2.n0 B2.t0 241.534
R28 B2.n0 B2.t1 169.234
R29 B2.n1 B2.n0 76
R30 B2.n1 B2 9.994
R31 B2 B2.n1 1.928
R32 VGND.n2 VGND.t1 107.701
R33 VGND.n9 VGND.t0 103.506
R34 VGND.n1 VGND.n0 92.5
R35 VGND.n4 VGND.n3 92.5
R36 VGND.n0 VGND.t3 72.923
R37 VGND.n3 VGND.t2 24.923
R38 VGND.n2 VGND.n1 8.18
R39 VGND.n10 VGND.n9 4.65
R40 VGND.n6 VGND.n5 4.65
R41 VGND.n8 VGND.n7 4.65
R42 VGND.n5 VGND.n4 1.113
R43 VGND.n6 VGND.n2 0.142
R44 VGND.n8 VGND.n6 0.119
R45 VGND.n10 VGND.n8 0.119
R46 VGND VGND.n10 0.022
R47 VNB VNB.t0 6078.09
R48 VNB.t2 VNB.t3 4931.87
R49 VNB.t4 VNB.t1 2030.77
R50 VNB.t3 VNB.t4 2030.77
R51 VNB.t0 VNB.t2 2030.77
R52 Y.n0 Y.t0 177.026
R53 Y.n3 Y.n1 99.746
R54 Y.n3 Y.n2 92.5
R55 Y.n2 Y.t2 24.923
R56 Y.n2 Y.t1 24.923
R57 Y.n1 Y 6.023
R58 Y Y.n3 4.018
R59 Y.n1 Y.n0 3.304
R60 Y.n0 Y 2.615
R61 a_481_47.t0 a_481_47.t1 49.846
R62 A1_N.n0 A1_N.t0 241.534
R63 A1_N.n0 A1_N.t1 169.234
R64 A1_N.n1 A1_N.n0 76
R65 A1_N.n1 A1_N 9.859
R66 A1_N A1_N.n1 1.902
C0 VGND Y 0.12fF
C1 B2 B1 0.16fF
C2 A1_N A2_N 0.10fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__a2bb2oi_2.ext - technology: sky130A

.subckt sky130_fd_sc_hd__a2bb2oi_2 A2_N A1_N Y B2 B1 VGND VPWR VNB VPB
X0 a_54_297.t2 B1.t0 VPWR.t2 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_442_21.t4 A1_N.t0 VGND.t7 VNB.t8 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 VPWR.t0 B2.t0 a_54_297.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 a_442_21.t0 A2_N.t0 VGND.t4 VNB.t5 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 Y.t5 B2.t1 a_136_47.t3 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 VPWR.t3 A1_N.t1 a_662_297.t1 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 a_54_297.t5 B2.t2 VPWR.t5 VPB.t8 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 a_136_47.t1 B1.t1 VGND.t1 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 VGND.t6 A1_N.t2 a_442_21.t3 VNB.t7 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 VGND.t5 A2_N.t1 a_442_21.t1 VNB.t6 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 a_136_47.t2 B2.t3 Y.t4 VNB.t9 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 Y.t1 a_442_21.t6 VGND.t2 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 VPWR.t1 B1.t2 a_54_297.t1 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13 a_662_297.t3 A2_N.t2 a_442_21.t2 VPB.t5 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14 VGND.t0 B1.t3 a_136_47.t0 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X15 VGND.t3 a_442_21.t7 Y.t0 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X16 a_442_21.t5 A2_N.t3 a_662_297.t2 VPB.t9 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17 a_662_297.t0 A1_N.t3 VPWR.t4 VPB.t7 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X18 a_54_297.t3 a_442_21.t8 Y.t3 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X19 Y.t2 a_442_21.t9 a_54_297.t4 VPB.t6 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
R0 B1.n2 B1.t2 241.534
R1 B1.n0 B1.t0 241.534
R2 B1.n2 B1.t1 169.234
R3 B1.n0 B1.t3 169.234
R4 B1.n1 B1.n0 164.892
R5 B1.n3 B1.n2 76
R6 B1.n3 B1 9.481
R7 B1.n1  7.905
R8  B1.n1 2.488
R9  B1.n3 1.422
R10 VPWR.n3 VPWR.n2 318.066
R11 VPWR.n1 VPWR.n0 314.004
R12 VPWR.n7 VPWR.n6 314.004
R13 VPWR.n2 VPWR.t4 26.595
R14 VPWR.n2 VPWR.t3 26.595
R15 VPWR.n0 VPWR.t2 26.595
R16 VPWR.n0 VPWR.t0 26.595
R17 VPWR.n6 VPWR.t5 26.595
R18 VPWR.n6 VPWR.t1 26.595
R19 VPWR.n5 VPWR.n4 4.65
R20 VPWR.n8 VPWR.n7 4.147
R21 VPWR.n3 VPWR.n1 3.927
R22 VPWR.n5 VPWR.n3 0.14
R23 VPWR.n8 VPWR.n5 0.132
R24 VPWR VPWR.n8 0.129
R25 a_54_297.n2 a_54_297.t3 238.141
R26 a_54_297.n1 a_54_297.t1 226.103
R27 a_54_297.n1 a_54_297.n0 155.085
R28 a_54_297.n3 a_54_297.n2 142.024
R29 a_54_297.n2 a_54_297.n1 57.484
R30 a_54_297.n0 a_54_297.t0 26.595
R31 a_54_297.n0 a_54_297.t5 26.595
R32 a_54_297.n3 a_54_297.t4 26.595
R33 a_54_297.t2 a_54_297.n3 26.595
R34 VPB.t3 VPB.t4 556.386
R35 VPB VPB.t1 272.274
R36 VPB.t9 VPB.t5 248.598
R37 VPB.t7 VPB.t9 248.598
R38 VPB.t4 VPB.t7 248.598
R39 VPB.t6 VPB.t3 248.598
R40 VPB.t2 VPB.t6 248.598
R41 VPB.t0 VPB.t2 248.598
R42 VPB.t8 VPB.t0 248.598
R43 VPB.t1 VPB.t8 248.598
R44 A1_N.n0 A1_N.t3 212.079
R45 A1_N.n1 A1_N.t1 212.079
R46 A1_N.n0 A1_N.t2 139.779
R47 A1_N.n1 A1_N.t0 139.779
R48 A1_N A1_N.n2 76.786
R49 A1_N.n2 A1_N.n0 32.133
R50 A1_N.n2 A1_N.n1 29.212
R51 VGND.n2 VGND.t5 122.033
R52 VGND.n1 VGND.n0 115.464
R53 VGND.n16 VGND.n15 115.464
R54 VGND.n25 VGND.t1 114.4
R55 VGND.n6 VGND.n5 92.5
R56 VGND.n10 VGND.n9 92.5
R57 VGND.n5 VGND.t7 24.923
R58 VGND.n9 VGND.t3 24.923
R59 VGND.n0 VGND.t4 24.923
R60 VGND.n0 VGND.t6 24.923
R61 VGND.n15 VGND.t2 24.923
R62 VGND.n15 VGND.t0 24.923
R63 VGND.n26 VGND.n25 17.073
R64 VGND.n2 VGND.n1 11.091
R65 VGND.n4 VGND.n3 4.65
R66 VGND.n8 VGND.n7 4.65
R67 VGND.n12 VGND.n11 4.65
R68 VGND.n14 VGND.n13 4.65
R69 VGND.n18 VGND.n17 4.65
R70 VGND.n20 VGND.n19 4.65
R71 VGND.n22 VGND.n21 4.65
R72 VGND.n24 VGND.n23 4.65
R73 VGND.n11 VGND.n10 1.5
R74 VGND.n17 VGND.n16 0.376
R75 VGND.n4 VGND.n2 0.334
R76 VGND.n7 VGND.n6 0.3
R77 VGND.n8 VGND.n4 0.119
R78 VGND.n12 VGND.n8 0.119
R79 VGND.n14 VGND.n12 0.119
R80 VGND.n18 VGND.n14 0.119
R81 VGND.n20 VGND.n18 0.119
R82 VGND.n22 VGND.n20 0.119
R83 VGND.n24 VGND.n22 0.119
R84 VGND.n26 VGND.n24 0.119
R85 VGND VGND.n26 0.022
R86 a_442_21.n3 a_442_21.n0 286.978
R87 a_442_21.n2 a_442_21.t8 212.079
R88 a_442_21.n1 a_442_21.t9 212.079
R89 a_442_21.n2 a_442_21.t7 139.779
R90 a_442_21.n1 a_442_21.t6 139.779
R91 a_442_21.n3 a_442_21.n2 106.672
R92 a_442_21.n5 a_442_21.n4 88.89
R93 a_442_21.n2 a_442_21.n1 61.345
R94 a_442_21.n5 a_442_21.n3 60.635
R95 a_442_21.n6 a_442_21.n5 52.624
R96 a_442_21.n0 a_442_21.t2 26.595
R97 a_442_21.n0 a_442_21.t5 26.595
R98 a_442_21.n4 a_442_21.t1 24.923
R99 a_442_21.n4 a_442_21.t0 24.923
R100 a_442_21.n6 a_442_21.t3 24.923
R101 a_442_21.t4 a_442_21.n6 24.923
R102 VNB VNB.t2 6730.83
R103 VNB.t3 VNB.t8 4545.05
R104 VNB.t5 VNB.t6 2030.77
R105 VNB.t7 VNB.t5 2030.77
R106 VNB.t8 VNB.t7 2030.77
R107 VNB.t4 VNB.t3 2030.77
R108 VNB.t1 VNB.t4 2030.77
R109 VNB.t9 VNB.t1 2030.77
R110 VNB.t0 VNB.t9 2030.77
R111 VNB.t2 VNB.t0 2030.77
R112 B2.n0 B2.t0 212.079
R113 B2.n1 B2.t2 212.079
R114 B2.n0 B2.t3 139.779
R115 B2.n1 B2.t1 139.779
R116 B2 B2.n2 86.88
R117 B2.n2 B2.n0 30.672
R118 B2.n2 B2.n1 30.672
R119 A2_N.n0 A2_N.t2 212.079
R120 A2_N.n1 A2_N.t3 212.079
R121 A2_N.n0 A2_N.t1 139.779
R122 A2_N.n1 A2_N.t0 139.779
R123 A2_N A2_N.n2 79.84
R124 A2_N.n2 A2_N.n1 32.133
R125 A2_N.n2 A2_N.n0 29.212
R126 a_136_47.n1 a_136_47.n0 187.937
R127 a_136_47.n0 a_136_47.t0 24.923
R128 a_136_47.n0 a_136_47.t2 24.923
R129 a_136_47.n1 a_136_47.t3 24.923
R130 a_136_47.t1 a_136_47.n1 24.923
R131 Y.n3 Y.n1 166.756
R132 Y Y.n0 158.134
R133 Y.n3 Y.n2 52.624
R134 Y.n0 Y.t3 26.595
R135 Y.n0 Y.t2 26.595
R136 Y.n2 Y.t0 24.923
R137 Y.n2 Y.t1 24.923
R138 Y.n1 Y.t4 24.923
R139 Y.n1 Y.t5 24.923
R140  Y 15.006
R141  Y.n3 12.317
R142 a_662_297.t1 a_662_297.n1 236.185
R143 a_662_297.n1 a_662_297.t3 194.328
R144 a_662_297.n1 a_662_297.n0 142.024
R145 a_662_297.n0 a_662_297.t2 26.595
R146 a_662_297.n0 a_662_297.t0 26.595
C0 Y VGND 0.22fF
C1 VPWR VPB 0.11fF
C2 B1 B2 0.30fF
C3 Y B1 0.11fF
C4 VGND VPWR 0.12fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__a2bb2oi_4.ext - technology: sky130A

.subckt sky130_fd_sc_hd__a2bb2oi_4 Y A2_N B2 A1_N B1 VGND VPWR VNB VPB
X0 Y.t8 B2.t0 a_109_47.t4 VNB.t13 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 VGND.t7 B1.t0 a_109_47.t7 VNB.t19 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 VGND.t8 a_751_21.t12 Y.t2 VNB.t5 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 a_751_21.t5 A2_N.t0 a_1139_297.t7 VPB.t15 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 a_1139_297.t0 A1_N.t0 VPWR.t7 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 VPWR.t11 B2.t1 a_27_297.t7 VPB.t11 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 VGND.t12 A2_N.t1 a_751_21.t6 VNB.t9 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 a_27_297.t6 B2.t2 VPWR.t10 VPB.t10 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 VPWR.t6 A1_N.t1 a_1139_297.t1 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 Y.t3 a_751_21.t13 VGND.t9 VNB.t6 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 a_1139_297.t2 A1_N.t2 VPWR.t5 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 VPWR.t0 B1.t1 a_27_297.t3 VPB.t7 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 a_27_297.t11 a_751_21.t14 Y.t4 VPB.t19 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13 Y.t9 a_751_21.t15 a_27_297.t10 VPB.t18 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14 VPWR.t4 A1_N.t3 a_1139_297.t3 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 a_751_21.t0 A1_N.t4 VGND.t0 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X16 a_27_297.t2 B1.t2 VPWR.t3 VPB.t6 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17 a_27_297.t9 a_751_21.t16 Y.t10 VPB.t17 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X18 VGND.t6 B1.t3 a_109_47.t5 VNB.t17 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X19 Y.t7 B2.t3 a_109_47.t3 VNB.t12 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X20 Y.t11 a_751_21.t17 a_27_297.t8 VPB.t16 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X21 a_1139_297.t6 A2_N.t2 a_751_21.t7 VPB.t14 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X22 a_751_21.t2 A2_N.t3 a_1139_297.t5 VPB.t13 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X23 a_27_297.t1 B1.t4 VPWR.t2 VPB.t5 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X24 VGND.t1 A1_N.t5 a_751_21.t1 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X25 VGND.t13 A1_N.t6 a_751_21.t8 VNB.t14 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X26 a_109_47.t6 B1.t5 VGND.t5 VNB.t18 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X27 VGND.t10 A2_N.t4 a_751_21.t3 VNB.t7 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X28 a_109_47.t2 B2.t4 Y.t6 VNB.t11 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X29 VPWR.t9 B2.t5 a_27_297.t5 VPB.t9 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X30 a_109_47.t1 B2.t6 Y.t5 VNB.t10 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X31 Y.t0 a_751_21.t18 VGND.t2 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X32 a_27_297.t4 B2.t7 VPWR.t8 VPB.t8 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X33 a_751_21.t9 A1_N.t7 VGND.t14 VNB.t15 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X34 a_751_21.t4 A2_N.t5 VGND.t11 VNB.t8 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X35 VPWR.t1 B1.t6 a_27_297.t0 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X36 a_1139_297.t4 A2_N.t6 a_751_21.t10 VPB.t12 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X37 a_109_47.t0 B1.t7 VGND.t4 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X38 VGND.t3 a_751_21.t19 Y.t1 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X39 a_751_21.t11 A2_N.t7 VGND.t15 VNB.t16 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
R0 B2.n1 B2.t7 212.079
R1 B2.n0 B2.t5 212.079
R2 B2.n3 B2.t1 212.079
R3 B2.n6 B2.t2 212.079
R4 B2.n1 B2.t0 139.779
R5 B2.n0 B2.t6 139.779
R6 B2.n3 B2.t4 139.779
R7 B2.n6 B2.t3 139.779
R8 B2 B2.n7 82.4
R9 B2.n5 B2.n4 76
R10 B2.n5 B2.n2 55.015
R11 B2.n2 B2.n0 33.414
R12 B2.n7 B2.n6 23.369
R13 B2.n2 B2.n1 16.893
R14 B2 B2.n5 15.36
R15 B2.n4 B2.n3 11.684
R16 a_109_47.n2 a_109_47.n0 141.372
R17 a_109_47.n5 a_109_47.n4 101.197
R18 a_109_47.n2 a_109_47.n1 92.5
R19 a_109_47.n4 a_109_47.n2 53.163
R20 a_109_47.n4 a_109_47.n3 42.273
R21 a_109_47.n3 a_109_47.t3 24.923
R22 a_109_47.n3 a_109_47.t6 24.923
R23 a_109_47.n1 a_109_47.t4 24.923
R24 a_109_47.n1 a_109_47.t2 24.923
R25 a_109_47.n0 a_109_47.t7 24.923
R26 a_109_47.n0 a_109_47.t1 24.923
R27 a_109_47.n5 a_109_47.t5 24.923
R28 a_109_47.t0 a_109_47.n5 24.923
R29 Y.n8 Y.n7 155.853
R30 Y.n11 Y.n10 146.391
R31 Y.n5 Y.n4 133.853
R32 Y.n5 Y.n3 92.5
R33 Y.n2 Y.n1 89.029
R34 Y.n6 Y.n5 69.961
R35 Y.n2 Y.n0 52.512
R36 Y.n8 Y.n6 45.929
R37 Y.n9 Y.n8 37.12
R38 Y.n10 Y.t4 26.595
R39 Y.n10 Y.t9 26.595
R40 Y.n7 Y.t10 26.595
R41 Y.n7 Y.t11 26.595
R42 Y.n3 Y.t5 24.923
R43 Y.n3 Y.t8 24.923
R44 Y.n4 Y.t6 24.923
R45 Y.n4 Y.t7 24.923
R46 Y.n1 Y.t1 24.923
R47 Y.n1 Y.t3 24.923
R48 Y.n0 Y.t2 24.923
R49 Y.n0 Y.t0 24.923
R50 Y.n11 Y.n9 10.753
R51 Y.n6 Y.n2 5.883
R52  Y.n11 4.805
R53 Y.n9 Y 4.072
R54 VNB VNB.t4 6053.91
R55 VNB.t3 VNB.t0 4545.05
R56 VNB.t16 VNB.t9 2030.77
R57 VNB.t7 VNB.t16 2030.77
R58 VNB.t8 VNB.t7 2030.77
R59 VNB.t14 VNB.t8 2030.77
R60 VNB.t15 VNB.t14 2030.77
R61 VNB.t1 VNB.t15 2030.77
R62 VNB.t0 VNB.t1 2030.77
R63 VNB.t6 VNB.t3 2030.77
R64 VNB.t5 VNB.t6 2030.77
R65 VNB.t2 VNB.t5 2030.77
R66 VNB.t19 VNB.t2 2030.77
R67 VNB.t10 VNB.t19 2030.77
R68 VNB.t13 VNB.t10 2030.77
R69 VNB.t11 VNB.t13 2030.77
R70 VNB.t12 VNB.t11 2030.77
R71 VNB.t18 VNB.t12 2030.77
R72 VNB.t17 VNB.t18 2030.77
R73 VNB.t4 VNB.t17 2030.77
R74 B1.n3 B1.n0 250.368
R75 B1.n0 B1.t4 241.534
R76 B1.n1 B1.t1 212.079
R77 B1.n4 B1.t2 212.079
R78 B1.n7 B1.t6 212.079
R79 B1.n0 B1.t0 169.234
R80 B1.n1 B1.t5 139.779
R81 B1.n4 B1.t3 139.779
R82 B1.n7 B1.t7 139.779
R83 B1.n3 B1.n2 76
R84 B1.n6 B1.n5 76
R85 B1.n9 B1.n8 76
R86 B1 B1.n9 24.685
R87 B1.n6 B1.n3 20.723
R88 B1.n9 B1.n6 20.723
R89 B1.n8 B1.n7 12.415
R90 B1.n2 B1.n1 10.954
R91 B1.n5 B1.n4 0.73
R92 VGND.n2 VGND.t12 204.569
R93 VGND.n1 VGND.n0 115.464
R94 VGND.n6 VGND.n5 115.464
R95 VGND.n12 VGND.n11 115.464
R96 VGND.n28 VGND.n27 115.464
R97 VGND.n34 VGND.n33 115.464
R98 VGND.n46 VGND.n45 115.464
R99 VGND.n51 VGND.t4 114.4
R100 VGND.n18 VGND.n17 92.5
R101 VGND.n22 VGND.n21 92.5
R102 VGND.n17 VGND.t0 24.923
R103 VGND.n21 VGND.t3 24.923
R104 VGND.n0 VGND.t15 24.923
R105 VGND.n0 VGND.t10 24.923
R106 VGND.n5 VGND.t11 24.923
R107 VGND.n5 VGND.t13 24.923
R108 VGND.n11 VGND.t14 24.923
R109 VGND.n11 VGND.t1 24.923
R110 VGND.n27 VGND.t9 24.923
R111 VGND.n27 VGND.t8 24.923
R112 VGND.n33 VGND.t2 24.923
R113 VGND.n33 VGND.t7 24.923
R114 VGND.n45 VGND.t5 24.923
R115 VGND.n45 VGND.t6 24.923
R116 VGND.n2 VGND.n1 16.676
R117 VGND.n35 VGND.n34 12.8
R118 VGND.n52 VGND.n51 6.908
R119 VGND.n7 VGND.n6 6.776
R120 VGND.n29 VGND.n28 6.776
R121 VGND.n4 VGND.n3 4.65
R122 VGND.n8 VGND.n7 4.65
R123 VGND.n10 VGND.n9 4.65
R124 VGND.n14 VGND.n13 4.65
R125 VGND.n16 VGND.n15 4.65
R126 VGND.n20 VGND.n19 4.65
R127 VGND.n24 VGND.n23 4.65
R128 VGND.n26 VGND.n25 4.65
R129 VGND.n30 VGND.n29 4.65
R130 VGND.n32 VGND.n31 4.65
R131 VGND.n36 VGND.n35 4.65
R132 VGND.n38 VGND.n37 4.65
R133 VGND.n40 VGND.n39 4.65
R134 VGND.n42 VGND.n41 4.65
R135 VGND.n44 VGND.n43 4.65
R136 VGND.n48 VGND.n47 4.65
R137 VGND.n50 VGND.n49 4.65
R138 VGND.n47 VGND.n46 3.764
R139 VGND.n19 VGND.n18 1.4
R140 VGND.n13 VGND.n12 0.752
R141 VGND.n4 VGND.n2 0.398
R142 VGND.n23 VGND.n22 0.2
R143 VGND.n8 VGND.n4 0.119
R144 VGND.n10 VGND.n8 0.119
R145 VGND.n14 VGND.n10 0.119
R146 VGND.n16 VGND.n14 0.119
R147 VGND.n20 VGND.n16 0.119
R148 VGND.n24 VGND.n20 0.119
R149 VGND.n26 VGND.n24 0.119
R150 VGND.n30 VGND.n26 0.119
R151 VGND.n32 VGND.n30 0.119
R152 VGND.n36 VGND.n32 0.119
R153 VGND.n38 VGND.n36 0.119
R154 VGND.n40 VGND.n38 0.119
R155 VGND.n42 VGND.n40 0.119
R156 VGND.n44 VGND.n42 0.119
R157 VGND.n48 VGND.n44 0.119
R158 VGND.n50 VGND.n48 0.119
R159 VGND.n52 VGND.n50 0.119
R160 VGND VGND.n52 0.02
R161 a_751_21.n5 a_751_21.t14 212.079
R162 a_751_21.n1 a_751_21.t15 212.079
R163 a_751_21.n3 a_751_21.t16 212.079
R164 a_751_21.n2 a_751_21.t17 212.079
R165 a_751_21.n16 a_751_21.n0 198.996
R166 a_751_21.n17 a_751_21.n16 154.572
R167 a_751_21.n5 a_751_21.t19 139.779
R168 a_751_21.n1 a_751_21.t13 139.779
R169 a_751_21.n3 a_751_21.t12 139.779
R170 a_751_21.n2 a_751_21.t18 139.779
R171 a_751_21.n9 a_751_21.n7 98.074
R172 a_751_21.n7 a_751_21.n6 76
R173 a_751_21.n16 a_751_21.n15 72.475
R174 a_751_21.n3 a_751_21.n2 61.345
R175 a_751_21.n7 a_751_21.n4 59.577
R176 a_751_21.n9 a_751_21.n8 52.624
R177 a_751_21.n11 a_751_21.n10 52.624
R178 a_751_21.n13 a_751_21.n12 52.624
R179 a_751_21.n15 a_751_21.n14 52.624
R180 a_751_21.n11 a_751_21.n9 36.266
R181 a_751_21.n13 a_751_21.n11 36.266
R182 a_751_21.n15 a_751_21.n13 36.266
R183 a_751_21.n0 a_751_21.t10 26.595
R184 a_751_21.n0 a_751_21.t5 26.595
R185 a_751_21.n17 a_751_21.t7 26.595
R186 a_751_21.t2 a_751_21.n17 26.595
R187 a_751_21.n4 a_751_21.n1 26.101
R188 a_751_21.n14 a_751_21.t6 24.923
R189 a_751_21.n14 a_751_21.t11 24.923
R190 a_751_21.n8 a_751_21.t1 24.923
R191 a_751_21.n8 a_751_21.t0 24.923
R192 a_751_21.n10 a_751_21.t8 24.923
R193 a_751_21.n10 a_751_21.t9 24.923
R194 a_751_21.n12 a_751_21.t3 24.923
R195 a_751_21.n12 a_751_21.t4 24.923
R196 a_751_21.n4 a_751_21.n3 24.392
R197 a_751_21.n6 a_751_21.n5 21.178
R198 A2_N.n0 A2_N.t2 212.079
R199 A2_N.n2 A2_N.t3 212.079
R200 A2_N.n5 A2_N.t6 212.079
R201 A2_N.n8 A2_N.t0 212.079
R202 A2_N.n0 A2_N.t1 139.779
R203 A2_N.n2 A2_N.t7 139.779
R204 A2_N.n5 A2_N.t4 139.779
R205 A2_N.n8 A2_N.t5 139.779
R206 A2_N.n4 A2_N.n1 97.76
R207 A2_N A2_N.n9 85.92
R208 A2_N.n4 A2_N.n3 76
R209 A2_N.n7 A2_N.n6 76
R210 A2_N.n7 A2_N.n4 21.76
R211 A2_N.n9 A2_N.n8 18.257
R212 A2_N.n1 A2_N.n0 16.796
R213 A2_N A2_N.n7 11.84
R214 A2_N.n6 A2_N.n5 6.572
R215 A2_N.n3 A2_N.n2 5.112
R216 a_1139_297.n5 a_1139_297.n0 292.5
R217 a_1139_297.t6 a_1139_297.n5 228.355
R218 a_1139_297.n3 a_1139_297.t3 177.181
R219 a_1139_297.n3 a_1139_297.n2 111.291
R220 a_1139_297.n4 a_1139_297.n1 90.234
R221 a_1139_297.n5 a_1139_297.n4 67.338
R222 a_1139_297.n4 a_1139_297.n3 65.327
R223 a_1139_297.n0 a_1139_297.t5 26.595
R224 a_1139_297.n0 a_1139_297.t4 26.595
R225 a_1139_297.n1 a_1139_297.t7 26.595
R226 a_1139_297.n1 a_1139_297.t0 26.595
R227 a_1139_297.n2 a_1139_297.t1 26.595
R228 a_1139_297.n2 a_1139_297.t2 26.595
R229 VPB.t19 VPB.t3 556.386
R230 VPB.t13 VPB.t14 248.598
R231 VPB.t12 VPB.t13 248.598
R232 VPB.t15 VPB.t12 248.598
R233 VPB.t0 VPB.t15 248.598
R234 VPB.t1 VPB.t0 248.598
R235 VPB.t2 VPB.t1 248.598
R236 VPB.t3 VPB.t2 248.598
R237 VPB.t18 VPB.t19 248.598
R238 VPB.t17 VPB.t18 248.598
R239 VPB.t16 VPB.t17 248.598
R240 VPB.t5 VPB.t16 248.598
R241 VPB.t9 VPB.t5 248.598
R242 VPB.t8 VPB.t9 248.598
R243 VPB.t11 VPB.t8 248.598
R244 VPB.t10 VPB.t11 248.598
R245 VPB.t7 VPB.t10 248.598
R246 VPB.t6 VPB.t7 248.598
R247 VPB.t4 VPB.t6 248.598
R248 VPB VPB.t4 189.408
R249 A1_N.n0 A1_N.t0 212.079
R250 A1_N.n2 A1_N.t1 212.079
R251 A1_N.n7 A1_N.t2 212.079
R252 A1_N.n5 A1_N.t3 212.079
R253 A1_N.n0 A1_N.t6 139.779
R254 A1_N.n2 A1_N.t7 139.779
R255 A1_N.n7 A1_N.t5 139.779
R256 A1_N.n5 A1_N.t4 139.779
R257 A1_N.n9 A1_N.n6 97.76
R258 A1_N.n4 A1_N.n1 97.76
R259 A1_N.n4 A1_N.n3 76
R260 A1_N.n9 A1_N.n8 76
R261 A1_N.n1 A1_N.n0 19.718
R262 A1_N.n6 A1_N.n5 15.336
R263 A1_N A1_N.n4 13.12
R264 A1_N A1_N.n9 8.64
R265 A1_N.n3 A1_N.n2 8.033
R266 A1_N.n8 A1_N.n7 3.651
R267 VPWR.n17 VPWR.n16 314.004
R268 VPWR.n21 VPWR.n20 314.004
R269 VPWR.n27 VPWR.n26 314.004
R270 VPWR.n1 VPWR.n0 176.855
R271 VPWR.n32 VPWR.n31 176.855
R272 VPWR.n3 VPWR.n2 175.589
R273 VPWR.n2 VPWR.t7 26.595
R274 VPWR.n2 VPWR.t6 26.595
R275 VPWR.n0 VPWR.t5 26.595
R276 VPWR.n0 VPWR.t4 26.595
R277 VPWR.n16 VPWR.t2 26.595
R278 VPWR.n16 VPWR.t9 26.595
R279 VPWR.n20 VPWR.t8 26.595
R280 VPWR.n20 VPWR.t11 26.595
R281 VPWR.n26 VPWR.t10 26.595
R282 VPWR.n26 VPWR.t0 26.595
R283 VPWR.n31 VPWR.t3 26.595
R284 VPWR.n31 VPWR.t1 26.595
R285 VPWR.n18 VPWR.n17 6.4
R286 VPWR.n5 VPWR.n4 4.65
R287 VPWR.n7 VPWR.n6 4.65
R288 VPWR.n9 VPWR.n8 4.65
R289 VPWR.n11 VPWR.n10 4.65
R290 VPWR.n13 VPWR.n12 4.65
R291 VPWR.n15 VPWR.n14 4.65
R292 VPWR.n19 VPWR.n18 4.65
R293 VPWR.n23 VPWR.n22 4.65
R294 VPWR.n25 VPWR.n24 4.65
R295 VPWR.n28 VPWR.n27 4.65
R296 VPWR.n30 VPWR.n29 4.65
R297 VPWR.n33 VPWR.n32 4.05
R298 VPWR.n3 VPWR.n1 3.856
R299 VPWR.n22 VPWR.n21 3.388
R300 VPWR.n5 VPWR.n3 0.232
R301 VPWR.n33 VPWR.n30 0.134
R302 VPWR VPWR.n33 0.124
R303 VPWR.n7 VPWR.n5 0.119
R304 VPWR.n9 VPWR.n7 0.119
R305 VPWR.n11 VPWR.n9 0.119
R306 VPWR.n13 VPWR.n11 0.119
R307 VPWR.n15 VPWR.n13 0.119
R308 VPWR.n19 VPWR.n15 0.119
R309 VPWR.n23 VPWR.n19 0.119
R310 VPWR.n25 VPWR.n23 0.119
R311 VPWR.n28 VPWR.n25 0.119
R312 VPWR.n30 VPWR.n28 0.119
R313 a_27_297.n8 a_27_297.t0 189.54
R314 a_27_297.n1 a_27_297.t11 175.231
R315 a_27_297.n1 a_27_297.n0 154.914
R316 a_27_297.n5 a_27_297.n4 154.573
R317 a_27_297.n7 a_27_297.n6 154.573
R318 a_27_297.n3 a_27_297.n2 142.024
R319 a_27_297.n9 a_27_297.n8 98.233
R320 a_27_297.n3 a_27_297.n1 56.972
R321 a_27_297.n5 a_27_297.n3 56.972
R322 a_27_297.n8 a_27_297.n7 49.833
R323 a_27_297.n7 a_27_297.n5 44.423
R324 a_27_297.n2 a_27_297.t8 26.595
R325 a_27_297.n2 a_27_297.t1 26.595
R326 a_27_297.n0 a_27_297.t10 26.595
R327 a_27_297.n0 a_27_297.t9 26.595
R328 a_27_297.n4 a_27_297.t5 26.595
R329 a_27_297.n4 a_27_297.t4 26.595
R330 a_27_297.n6 a_27_297.t7 26.595
R331 a_27_297.n6 a_27_297.t6 26.595
R332 a_27_297.t3 a_27_297.n9 26.595
R333 a_27_297.n9 a_27_297.t2 26.595
C0 Y VGND 0.42fF
C1 B2 B1 0.53fF
C2 B2 Y 0.24fF
C3 VPWR VGND 0.20fF
C4 Y B1 0.14fF
C5 VPWR VPB 0.18fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__a21bo_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__a21bo_1 X A1 B1_N A2 VGND VPWR VNB VPB
X0 a_298_297.t2 a_27_413.t2 a_215_297.t2 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_215_297.t1 a_27_413.t3 VGND.t3 VNB sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 a_298_297.t0 A2.t0 VPWR.t1 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 X.t1 a_215_297.t3 VGND.t0 VNB sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 VPWR.t2 B1_N.t0 a_27_413.t0 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 X.t0 a_215_297.t4 VPWR.t0 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 a_382_47.t0 A1.t0 a_215_297.t0 VNB sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 VGND.t2 B1_N.t1 a_27_413.t1 VNB sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 VPWR.t3 A1.t1 a_298_297.t1 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 VGND.t1 A2.t1 a_382_47.t1 VNB sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
R0 a_27_413.t0 a_27_413.n1 403.045
R1 a_27_413.n1 a_27_413.n0 238.63
R2 a_27_413.n0 a_27_413.t3 200.833
R3 a_27_413.n0 a_27_413.t2 192.799
R4 a_27_413.n1 a_27_413.t1 182.643
R5 a_215_297.n0 a_215_297.t4 231.242
R6 a_215_297.n2 a_215_297.n0 168.397
R7 a_215_297.t2 a_215_297.n2 166.42
R8 a_215_297.n0 a_215_297.t3 158.942
R9 a_215_297.n2 a_215_297.n1 48.65
R10 a_215_297.n1 a_215_297.t0 24.923
R11 a_215_297.n1 a_215_297.t1 24.923
R12 a_298_297.t0 a_298_297.n0 384.249
R13 a_298_297.n0 a_298_297.t1 26.595
R14 a_298_297.n0 a_298_297.t2 26.595
R15 VPB.t0 VPB.t1 559.345
R16 VPB.t2 VPB.t4 559.345
R17 VPB.t3 VPB.t0 254.517
R18 VPB.t4 VPB.t3 248.598
R19 VPB VPB.t2 192.367
R20 VGND.n3 VGND.n2 92.5
R21 VGND.n5 VGND.n4 92.5
R22 VGND.n1 VGND.n0 70.811
R23 VGND.n0 VGND.t2 67.309
R24 VGND.n0 VGND.t3 42.065
R25 VGND.n2 VGND.t0 41.538
R26 VGND.n4 VGND.t1 40.615
R27 VGND.n7 VGND.n3 6.102
R28 VGND.n7 VGND.n6 4.65
R29 VGND.n9 VGND.n8 4.65
R30 VGND.n11 VGND.n10 4.65
R31 VGND.n12 VGND.n1 3.86
R32 VGND.n6 VGND.n5 0.711
R33 VGND VGND.n12 0.239
R34 VGND.n12 VGND.n11 0.141
R35 VGND.n9 VGND.n7 0.119
R36 VGND.n11 VGND.n9 0.119
R37 A2.n0 A2.t0 231.014
R38 A2.n0 A2.t1 158.714
R39 A2.n1 A2.n0 76
R40 A2.n1 A2 14.03
R41 A2 A2.n1 2.707
R42 VPWR.n7 VPWR.t2 369.718
R43 VPWR.n1 VPWR.n0 311.118
R44 VPWR.n2 VPWR.t0 152.846
R45 VPWR.n0 VPWR.t1 27.58
R46 VPWR.n0 VPWR.t3 27.58
R47 VPWR.n4 VPWR.n3 4.65
R48 VPWR.n6 VPWR.n5 4.65
R49 VPWR.n8 VPWR.n7 3.932
R50 VPWR.n2 VPWR.n1 3.878
R51 VPWR.n4 VPWR.n2 0.226
R52 VPWR.n8 VPWR.n6 0.137
R53 VPWR VPWR.n8 0.123
R54 VPWR.n6 VPWR.n4 0.119
R55 X.n0 X.t0 207.034
R56 X.n1 X.t1 117.423
R57 X.n1 X 8.914
R58 X X.n0 8.176
R59 X.n0 X 7.11
R60 X X.n1 6.628
R61 B1_N.n1 B1_N.t1 299.91
R62 B1_N.n0 B1_N.t0 199.761
R63 B1_N.n0 B1_N 79.06
R64 B1_N.n2 B1_N.n1 76
R65 B1_N.n1 B1_N.n0 60.696
R66 B1_N.n2 B1_N 15.86
R67 B1_N B1_N.n2 3.06
R68 A1.n0 A1.t1 241.534
R69 A1.n0 A1.t0 169.234
R70 A1.n1 A1.n0 76
R71 A1.n1 A1 8.583
R72 A1 A1.n1 1.656
R73 a_382_47.t0 a_382_47.t1 51.692
C0 A2 A1 0.15fF
C1 X VPWR 0.13fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__a21bo_2.ext - technology: sky130A

.subckt sky130_fd_sc_hd__a21bo_2 B1_N A2 X A1 VGND VPWR VNB VPB
X0 VPWR.t0 A1.t0 a_485_297.t1 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_485_297.t0 a_297_93.t2 a_79_21.t1 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 a_297_93.t0 B1_N.t0 VGND.t2 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3 a_581_47.t0 A1.t1 a_79_21.t0 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 VGND.t1 a_79_21.t3 X.t3 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 a_79_21.t2 a_297_93.t3 VGND.t4 VNB.t5 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 VGND.t3 A2.t0 a_581_47.t1 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 VPWR.t3 a_79_21.t4 X.t1 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 a_297_93.t1 B1_N.t1 VPWR.t1 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9 X.t0 a_79_21.t5 VPWR.t4 VPB.t5 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 a_485_297.t2 A2.t1 VPWR.t2 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 X.t2 a_79_21.t6 VGND.t0 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
R0 A1.n0 A1.t0 241.534
R1 A1.n0 A1.t1 169.234
R2 A1 A1.n0 84.79
R3 a_485_297.n0 a_485_297.t2 369.376
R4 a_485_297.n0 a_485_297.t1 26.595
R5 a_485_297.t0 a_485_297.n0 26.595
R6 VPWR.n6 VPWR.t4 575.999
R7 VPWR.n2 VPWR.n1 390.244
R8 VPWR.n3 VPWR.n0 317.98
R9 VPWR.n1 VPWR.t1 103.19
R10 VPWR.n1 VPWR.t3 27.293
R11 VPWR.n0 VPWR.t2 26.595
R12 VPWR.n0 VPWR.t0 26.595
R13 VPWR.n5 VPWR.n4 4.65
R14 VPWR.n7 VPWR.n6 4.65
R15 VPWR.n3 VPWR.n2 3.825
R16 VPWR.n5 VPWR.n3 0.144
R17 VPWR.n7 VPWR.n5 0.119
R18 VPWR VPWR.n7 0.02
R19 VPB.t2 VPB.t0 556.386
R20 VPB.t4 VPB.t2 301.869
R21 VPB.t5 VPB.t4 254.517
R22 VPB.t1 VPB.t3 248.598
R23 VPB.t0 VPB.t1 248.598
R24 VPB VPB.t5 189.408
R25 a_297_93.n1 a_297_93.t1 389.585
R26 a_297_93.n0 a_297_93.t2 229
R27 a_297_93.t0 a_297_93.n1 160.318
R28 a_297_93.n0 a_297_93.t3 155.607
R29 a_297_93.n1 a_297_93.n0 76
R30 a_79_21.n1 a_79_21.t4 221.719
R31 a_79_21.n2 a_79_21.t5 221.719
R32 a_79_21.n4 a_79_21.n0 189.6
R33 a_79_21.n4 a_79_21.n3 186.715
R34 a_79_21.t1 a_79_21.n4 170.634
R35 a_79_21.n1 a_79_21.t3 149.419
R36 a_79_21.n2 a_79_21.t6 149.419
R37 a_79_21.n3 a_79_21.n2 47.307
R38 a_79_21.n0 a_79_21.t0 33.23
R39 a_79_21.n3 a_79_21.n1 29.455
R40 a_79_21.n0 a_79_21.t2 27.692
R41 B1_N.n0 B1_N.t1 148.348
R42 B1_N.n0 B1_N.t0 132.281
R43 B1_N B1_N.n0 92.33
R44 VGND.n1 VGND.t3 208.413
R45 VGND.n9 VGND.t0 194.65
R46 VGND.n0 VGND.t4 190.315
R47 VGND.n5 VGND.n4 74.159
R48 VGND.n4 VGND.t2 62.857
R49 VGND.n4 VGND.t1 25.846
R50 VGND.n10 VGND.n9 4.65
R51 VGND.n3 VGND.n2 4.65
R52 VGND.n6 VGND.n5 4.65
R53 VGND.n8 VGND.n7 4.65
R54 VGND.n1 VGND.n0 3.775
R55 VGND.n3 VGND.n1 0.159
R56 VGND.n6 VGND.n3 0.119
R57 VGND.n8 VGND.n6 0.119
R58 VGND.n10 VGND.n8 0.119
R59 VGND VGND.n10 0.02
R60 VNB VNB.t0 6053.91
R61 VNB.t3 VNB.t5 4545.05
R62 VNB.t1 VNB.t3 2465.93
R63 VNB.t5 VNB.t2 2320.88
R64 VNB.t0 VNB.t1 2079.12
R65 VNB.t2 VNB.t4 1740.66
R66 a_581_47.t0 a_581_47.t1 38.769
R67 X X.n0 174.098
R68 X X.n1 117.013
R69 X.n0 X.t1 27.58
R70 X.n0 X.t0 27.58
R71 X.n1 X.t3 25.846
R72 X.n1 X.t2 25.846
R73 A2.n0 A2.t1 233.287
R74 A2.n0 A2.t0 160.987
R75 A2 A2.n0 78.427
C0 A2 A1 0.17fF
C1 X VGND 0.19fF
C2 X VPWR 0.13fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__a21bo_4.ext - technology: sky130A

.subckt sky130_fd_sc_hd__a21bo_4 B1_N A2 A1 X VGND VPWR VNB VPB
X0 a_1021_47.t1 A1.t0 a_205_21.t5 VNB.t10 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 X.t7 a_205_21.t6 VPWR.t4 VPB.t8 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 VPWR.t3 a_205_21.t7 X.t6 VPB.t7 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 X.t3 a_205_21.t8 VGND.t7 VNB.t7 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 VGND.t2 A2.t0 a_1021_47.t0 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 VGND.t8 a_42_47.t2 a_205_21.t3 VNB.t8 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 a_861_47.t0 A2.t1 VGND.t3 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 a_205_21.t4 A1.t1 a_861_47.t1 VNB.t9 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 X.t5 a_205_21.t9 VPWR.t6 VPB.t6 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 a_603_297.t5 A1.t2 VPWR.t8 VPB.t10 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 VGND.t1 B1_N.t0 a_42_47.t0 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 VPWR.t2 A2.t2 a_603_297.t3 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 a_603_297.t1 a_42_47.t3 a_205_21.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13 VPWR.t5 a_205_21.t10 X.t4 VPB.t5 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14 a_205_21.t1 a_42_47.t4 a_603_297.t0 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 VGND.t6 a_205_21.t11 X.t2 VNB.t6 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X16 VPWR.t0 B1_N.t1 a_42_47.t1 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17 VGND.t5 a_205_21.t12 X.t1 VNB.t5 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X18 VPWR.t7 A1.t3 a_603_297.t4 VPB.t9 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X19 a_603_297.t2 A2.t3 VPWR.t1 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X20 a_205_21.t2 a_42_47.t5 VGND.t0 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X21 X.t0 a_205_21.t13 VGND.t4 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
R0 A1.n0 A1.t3 212.079
R1 A1.n1 A1.t2 212.079
R2 A1.n0 A1.t0 139.779
R3 A1.n1 A1.t1 139.779
R4 A1 A1.n2 77.928
R5 A1.n2 A1.n0 35.054
R6 A1.n2 A1.n1 26.29
R7 a_205_21.n13 a_205_21.n12 357.252
R8 a_205_21.n2 a_205_21.t10 212.079
R9 a_205_21.n6 a_205_21.t9 212.079
R10 a_205_21.n4 a_205_21.t7 212.079
R11 a_205_21.n3 a_205_21.t6 212.079
R12 a_205_21.n11 a_205_21.n1 179.262
R13 a_205_21.n2 a_205_21.t11 139.779
R14 a_205_21.n6 a_205_21.t13 139.779
R15 a_205_21.n4 a_205_21.t12 139.779
R16 a_205_21.n3 a_205_21.t8 139.779
R17 a_205_21.n12 a_205_21.n0 92.5
R18 a_205_21.n8 a_205_21.n5 89.187
R19 a_205_21.n10 a_205_21.n9 85.843
R20 a_205_21.n9 a_205_21.n2 84.033
R21 a_205_21.n8 a_205_21.n7 76
R22 a_205_21.n4 a_205_21.n3 62.806
R23 a_205_21.n5 a_205_21.n4 34.324
R24 a_205_21.t0 a_205_21.n13 26.595
R25 a_205_21.n13 a_205_21.t1 26.595
R26 a_205_21.n0 a_205_21.t3 24.923
R27 a_205_21.n0 a_205_21.t2 24.923
R28 a_205_21.n1 a_205_21.t5 24.923
R29 a_205_21.n1 a_205_21.t4 24.923
R30 a_205_21.n7 a_205_21.n6 21.178
R31 a_205_21.n9 a_205_21.n8 13.187
R32 a_205_21.n11 a_205_21.n10 4.141
R33 a_205_21.n12 a_205_21.n11 0.376
R34 a_1021_47.t0 a_1021_47.t1 49.846
R35 VNB VNB.t1 7045.12
R36 VNB.t6 VNB.t0 4641.76
R37 VNB.t8 VNB.t3 2224.18
R38 VNB.t4 VNB.t6 2079.12
R39 VNB.t5 VNB.t4 2079.12
R40 VNB.t7 VNB.t5 2079.12
R41 VNB.t1 VNB.t7 2079.12
R42 VNB.t10 VNB.t2 2030.77
R43 VNB.t9 VNB.t10 2030.77
R44 VNB.t0 VNB.t8 2030.77
R45 VNB.t3 VNB.t9 1837.36
R46 VPWR.n10 VPWR.t5 570.094
R47 VPWR.n3 VPWR.n2 309.949
R48 VPWR.n1 VPWR.n0 306.463
R49 VPWR.n15 VPWR.n14 306.463
R50 VPWR.n20 VPWR.n19 306.463
R51 VPWR.n14 VPWR.t6 27.58
R52 VPWR.n14 VPWR.t3 27.58
R53 VPWR.n19 VPWR.t4 27.58
R54 VPWR.n19 VPWR.t0 27.58
R55 VPWR.n2 VPWR.t1 26.595
R56 VPWR.n2 VPWR.t7 26.595
R57 VPWR.n0 VPWR.t8 26.595
R58 VPWR.n0 VPWR.t2 26.595
R59 VPWR.n21 VPWR.n20 6.405
R60 VPWR.n5 VPWR.n4 4.65
R61 VPWR.n7 VPWR.n6 4.65
R62 VPWR.n9 VPWR.n8 4.65
R63 VPWR.n11 VPWR.n10 4.65
R64 VPWR.n13 VPWR.n12 4.65
R65 VPWR.n16 VPWR.n15 4.65
R66 VPWR.n18 VPWR.n17 4.65
R67 VPWR.n3 VPWR.n1 3.759
R68 VPWR.n5 VPWR.n3 0.254
R69 VPWR.n21 VPWR.n18 0.132
R70 VPWR VPWR.n21 0.129
R71 VPWR.n7 VPWR.n5 0.119
R72 VPWR.n9 VPWR.n7 0.119
R73 VPWR.n11 VPWR.n9 0.119
R74 VPWR.n13 VPWR.n11 0.119
R75 VPWR.n16 VPWR.n13 0.119
R76 VPWR.n18 VPWR.n16 0.119
R77 X.n2 X.n0 357.252
R78 X.n2 X.n1 292.5
R79 X.n5 X.n3 157.252
R80 X.n5 X.n4 92.5
R81 X X.n5 46.601
R82 X.n1 X.t6 27.58
R83 X.n1 X.t7 27.58
R84 X.n0 X.t4 27.58
R85 X.n0 X.t5 27.58
R86 X.n4 X.t1 25.846
R87 X.n4 X.t3 25.846
R88 X.n3 X.t2 25.846
R89 X.n3 X.t0 25.846
R90 X X.n2 18.823
R91 VPB.t5 VPB.t1 568.224
R92 VPB VPB.t2 310.747
R93 VPB.t6 VPB.t5 254.517
R94 VPB.t7 VPB.t6 254.517
R95 VPB.t8 VPB.t7 254.517
R96 VPB.t2 VPB.t8 254.517
R97 VPB.t9 VPB.t3 248.598
R98 VPB.t10 VPB.t9 248.598
R99 VPB.t4 VPB.t10 248.598
R100 VPB.t0 VPB.t4 248.598
R101 VPB.t1 VPB.t0 248.598
R102 VGND.n2 VGND.t2 110.996
R103 VGND.n1 VGND.n0 106.463
R104 VGND.n16 VGND.n15 106.463
R105 VGND.n21 VGND.n20 106.052
R106 VGND.n6 VGND.n5 92.5
R107 VGND.n10 VGND.n9 92.5
R108 VGND.n9 VGND.t6 46.153
R109 VGND.n0 VGND.t8 32.307
R110 VGND.n5 VGND.t0 28.615
R111 VGND.n15 VGND.t4 25.846
R112 VGND.n15 VGND.t5 25.846
R113 VGND.n20 VGND.t7 25.846
R114 VGND.n20 VGND.t1 25.846
R115 VGND.n0 VGND.t3 24.923
R116 VGND.n22 VGND.n21 5.652
R117 VGND.n4 VGND.n3 4.65
R118 VGND.n8 VGND.n7 4.65
R119 VGND.n12 VGND.n11 4.65
R120 VGND.n14 VGND.n13 4.65
R121 VGND.n17 VGND.n16 4.65
R122 VGND.n19 VGND.n18 4.65
R123 VGND.n11 VGND.n10 4.467
R124 VGND.n2 VGND.n1 3.675
R125 VGND.n7 VGND.n6 3.139
R126 VGND.n4 VGND.n2 0.148
R127 VGND.n22 VGND.n19 0.132
R128 VGND VGND.n22 0.129
R129 VGND.n8 VGND.n4 0.119
R130 VGND.n12 VGND.n8 0.119
R131 VGND.n14 VGND.n12 0.119
R132 VGND.n17 VGND.n14 0.119
R133 VGND.n19 VGND.n17 0.119
R134 A2.n1 A2.t2 241.534
R135 A2.n0 A2.t3 241.534
R136 A2 A2.n1 172.619
R137 A2.n1 A2.t1 169.234
R138 A2.n0 A2.t0 169.234
R139 A2 A2.n0 98.835
R140 a_42_47.n2 a_42_47.n1 380.114
R141 a_42_47.n0 a_42_47.t3 212.079
R142 a_42_47.n1 a_42_47.t4 212.079
R143 a_42_47.t1 a_42_47.n2 176.523
R144 a_42_47.n2 a_42_47.t0 152.144
R145 a_42_47.n0 a_42_47.t2 139.779
R146 a_42_47.n1 a_42_47.t5 139.779
R147 a_42_47.n1 a_42_47.n0 61.345
R148 a_861_47.t0 a_861_47.t1 42.461
R149 a_603_297.n1 a_603_297.n0 292.5
R150 a_603_297.n2 a_603_297.t0 253.49
R151 a_603_297.n1 a_603_297.t2 234.435
R152 a_603_297.n3 a_603_297.n2 152.575
R153 a_603_297.n2 a_603_297.n1 58.146
R154 a_603_297.n0 a_603_297.t4 26.595
R155 a_603_297.n0 a_603_297.t5 26.595
R156 a_603_297.n3 a_603_297.t3 26.595
R157 a_603_297.t1 a_603_297.n3 26.595
R158 B1_N.n0 B1_N.t1 241.534
R159 B1_N.n0 B1_N.t0 169.234
R160 B1_N B1_N.n0 77.248
C0 A2 A1 0.27fF
C1 VGND X 0.14fF
C2 VGND VPWR 0.13fF
C3 VPB VPWR 0.12fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__a21boi_0.ext - technology: sky130A

.subckt sky130_fd_sc_hd__a21boi_0 B1_N Y A1 A2 VPWR VGND VNB VPB
X0 a_300_369.t0 A2.t0 VPWR.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1 a_400_47.t1 A1.t0 Y.t0 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 VGND.t0 A2.t1 a_400_47.t0 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3 VGND.t1 B1_N.t0 a_27_47.t0 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 VPWR.t1 B1_N.t1 a_27_47.t1 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 Y.t2 a_27_47.t2 VGND.t2 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 a_300_369.t1 a_27_47.t3 Y.t1 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X7 VPWR.t2 A1.t1 a_300_369.t2 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
R0 A2.n0 A2.t0 276.256
R1 A2.n0 A2.t1 141.134
R2 A2 A2.n0 40.391
R3 VPWR.n1 VPWR.t1 377.867
R4 VPWR.n1 VPWR.n0 322.024
R5 VPWR.n0 VPWR.t0 43.093
R6 VPWR.n0 VPWR.t2 43.093
R7 VPWR VPWR.n1 0.151
R8 a_300_369.t0 a_300_369.n0 405.117
R9 a_300_369.n0 a_300_369.t2 43.093
R10 a_300_369.n0 a_300_369.t1 43.093
R11 VPB.t1 VPB.t2 562.305
R12 VPB.t3 VPB.t0 254.517
R13 VPB.t2 VPB.t3 254.517
R14 VPB VPB.t1 195.327
R15 A1.n0 A1.t1 284.634
R16 A1.n0 A1.t0 155.914
R17 A1 A1.n0 35.334
R18 Y Y.t1 337.726
R19 Y Y.n0 161.011
R20 Y.n0 Y.t0 111.428
R21 Y.n0 Y.t2 40
R22 a_400_47.t0 a_400_47.t1 60
R23 VNB VNB.t2 6502.94
R24 VNB.t2 VNB.t3 4982.35
R25 VNB.t3 VNB.t1 4400
R26 VNB.t1 VNB.t0 2329.41
R27 VGND.n2 VGND.t0 153.373
R28 VGND.n1 VGND.n0 92.5
R29 VGND.n4 VGND.n3 92.5
R30 VGND.n0 VGND.t2 40
R31 VGND.n3 VGND.t1 40
R32 VGND.n2 VGND.n1 6.624
R33 VGND.n5 VGND.n4 4.036
R34 VGND.n5 VGND.n2 0.158
R35 VGND VGND.n5 0.126
R36 B1_N.n0 B1_N.t0 301.399
R37 B1_N.n0 B1_N.t1 162.31
R38 B1_N B1_N.n0 32.706
R39 a_27_47.n1 a_27_47.t1 440.237
R40 a_27_47.n0 a_27_47.t2 291.232
R41 a_27_47.n0 a_27_47.t3 229.621
R42 a_27_47.t0 a_27_47.n1 153.159
R43 a_27_47.n1 a_27_47.n0 112.075
C0 A1 Y 0.13fF
C1 A1 A2 0.22fF
C2 VGND Y 0.13fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__a21boi_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__a21boi_1 Y A1 B1_N A2 VPWR VGND VNB VPB
X0 a_300_297.t1 a_27_413.t2 Y.t1 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 VGND.t2 A2.t0 a_384_47.t1 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 VPWR.t1 B1_N.t0 a_27_413.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3 Y.t2 a_27_413.t3 VGND.t1 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 VPWR.t0 A1.t0 a_300_297.t0 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 a_384_47.t0 A1.t1 Y.t0 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 VGND.t0 B1_N.t1 a_27_413.t1 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7 a_300_297.t2 A2.t1 VPWR.t2 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
R0 a_27_413.t0 a_27_413.n1 403.417
R1 a_27_413.n0 a_27_413.t2 233.769
R2 a_27_413.n0 a_27_413.t3 200.833
R3 a_27_413.n1 a_27_413.n0 200.07
R4 a_27_413.n1 a_27_413.t1 176.821
R5 Y.n1 Y.n0 146.535
R6 Y.n3 Y.n2 92.5
R7 Y.n2 Y.t0 40.615
R8 Y.n2 Y.t2 40.615
R9 Y.n4 Y.n3 30.509
R10 Y.n0 Y.t1 27.58
R11 Y Y.n1 10.115
R12 Y.n5 Y 7.175
R13 Y.n4 Y 6.186
R14 Y Y.n5 6.012
R15 Y.n3 Y 4.018
R16 Y Y.n4 3.878
R17 Y.n1 Y 3.012
R18 a_300_297.n0 a_300_297.t2 418.863
R19 a_300_297.t0 a_300_297.n0 27.58
R20 a_300_297.n0 a_300_297.t1 27.58
R21 VPB.t0 VPB.t2 562.305
R22 VPB.t1 VPB.t3 254.517
R23 VPB.t2 VPB.t1 254.517
R24 VPB VPB.t0 195.327
R25 A2.n0 A2.t1 231.014
R26 A2.n0 A2.t0 158.714
R27 A2 A2.n0 78.427
R28 a_384_47.t0 a_384_47.t1 51.692
R29 VGND.n1 VGND.t2 106.963
R30 VGND.n1 VGND.n0 74.206
R31 VGND.n0 VGND.t0 57.778
R32 VGND.n0 VGND.t1 25.706
R33 VGND VGND.n1 0.259
R34 VNB VNB.t0 11776.5
R35 VNB.t2 VNB.t1 2852.75
R36 VNB.t0 VNB.t2 2327.87
R37 VNB.t1 VNB.t3 2079.12
R38 B1_N.n1 B1_N.t1 283.844
R39 B1_N.n0 B1_N.t0 201.368
R40 B1_N B1_N.n0 79.06
R41 B1_N.n2 B1_N.n1 76
R42 B1_N B1_N.n2 15.86
R43 B1_N.n2 B1_N 3.06
R44 VPWR.n1 VPWR.t1 376.315
R45 VPWR.n1 VPWR.n0 167.203
R46 VPWR.n0 VPWR.t2 27.58
R47 VPWR.n0 VPWR.t0 27.58
R48 VPWR VPWR.n1 0.152
R49 A1.n0 A1.t0 241.534
R50 A1.n0 A1.t1 169.234
R51 A1 A1.n0 80.754
C0 Y VGND 0.18fF
C1 A2 A1 0.11fF
C2 VGND A1 0.10fF
C3 Y A1 0.11fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__a21boi_2.ext - technology: sky130A

.subckt sky130_fd_sc_hd__a21boi_2 VPWR VGND B1_N A2 A1 Y VNB VPB
X0 Y.t5 a_61_47.t2 VGND.t3 VNB.t5 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 VPWR.t1 A2.t0 a_217_297.t1 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 a_217_297.t5 a_61_47.t3 Y.t3 VPB.t5 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 a_479_47.t0 A2.t1 VGND.t0 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 a_217_297.t0 A2.t2 VPWR.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 Y.t2 a_61_47.t4 a_217_297.t4 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 VPWR.t2 A1.t0 a_217_297.t2 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 a_61_47.t0 B1_N.t0 VPWR.t4 VPB.t6 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 VGND.t1 A2.t3 a_637_47.t0 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 VGND.t2 a_61_47.t5 Y.t4 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 Y.t1 A1.t1 a_479_47.t1 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 VGND.t4 B1_N.t1 a_61_47.t1 VNB.t6 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12 a_217_297.t3 A1.t2 VPWR.t3 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13 a_637_47.t1 A1.t3 Y.t0 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
R0 a_61_47.t0 a_61_47.n2 403.704
R1 a_61_47.n0 a_61_47.t3 218.506
R2 a_61_47.n1 a_61_47.t4 218.506
R3 a_61_47.n2 a_61_47.t1 200.092
R4 a_61_47.n0 a_61_47.t5 146.206
R5 a_61_47.n1 a_61_47.t2 146.206
R6 a_61_47.n2 a_61_47.n1 137.371
R7 a_61_47.n1 a_61_47.n0 69.806
R8 VGND.n3 VGND.n2 106.463
R9 VGND.n4 VGND.t1 95.237
R10 VGND.n0 VGND.t4 72.197
R11 VGND.n1 VGND.n0 70.646
R12 VGND.n0 VGND.t3 44.307
R13 VGND.n2 VGND.t2 35.076
R14 VGND.n2 VGND.t0 25.846
R15 VGND.n6 VGND.n5 4.65
R16 VGND.n7 VGND.n1 3.936
R17 VGND.n4 VGND.n3 3.868
R18 VGND VGND.n7 0.239
R19 VGND.n6 VGND.n4 0.143
R20 VGND.n7 VGND.n6 0.139
R21 Y.n2 Y.n1 207.378
R22 Y.n3 Y.n0 125.375
R23 Y Y.n4 92.82
R24 Y.n1 Y.t3 26.595
R25 Y.n1 Y.t2 26.595
R26 Y.n0 Y.t0 25.846
R27 Y.n0 Y.t1 25.846
R28 Y.n4 Y.t4 24.923
R29 Y.n4 Y.t5 24.923
R30 Y Y.n3 17.6
R31 Y.n3 Y.n2 3.84
R32 VNB VNB.t6 7821.6
R33 VNB.t6 VNB.t5 3536.66
R34 VNB.t4 VNB.t2 2320.88
R35 VNB.t0 VNB.t3 2079.12
R36 VNB.t1 VNB.t0 2079.12
R37 VNB.t5 VNB.t4 2030.77
R38 VNB.t2 VNB.t1 1740.66
R39 A2.n0 A2.t0 241.534
R40 A2.n1 A2.t2 239.684
R41 A2.n0 A2.t1 169.234
R42 A2.n1 A2.t3 167.384
R43 A2 A2.n0 167.183
R44 A2 A2.n1 88.578
R45 a_217_297.t4 a_217_297.n3 224.548
R46 a_217_297.n1 a_217_297.t0 217.093
R47 a_217_297.n1 a_217_297.n0 149.831
R48 a_217_297.n3 a_217_297.n2 143.026
R49 a_217_297.n3 a_217_297.n1 58.704
R50 a_217_297.n0 a_217_297.t2 27.58
R51 a_217_297.n0 a_217_297.t3 27.58
R52 a_217_297.n2 a_217_297.t1 26.595
R53 a_217_297.n2 a_217_297.t5 26.595
R54 VPWR.n12 VPWR.t4 379.693
R55 VPWR.n2 VPWR.n1 313.205
R56 VPWR.n3 VPWR.n0 309.862
R57 VPWR.n0 VPWR.t0 27.58
R58 VPWR.n0 VPWR.t2 27.58
R59 VPWR.n1 VPWR.t3 26.595
R60 VPWR.n1 VPWR.t1 26.595
R61 VPWR.n3 VPWR.n2 8.554
R62 VPWR.n5 VPWR.n4 4.65
R63 VPWR.n7 VPWR.n6 4.65
R64 VPWR.n9 VPWR.n8 4.65
R65 VPWR.n11 VPWR.n10 4.65
R66 VPWR.n13 VPWR.n12 4.65
R67 VPWR.n5 VPWR.n3 0.231
R68 VPWR.n7 VPWR.n5 0.119
R69 VPWR.n9 VPWR.n7 0.119
R70 VPWR.n11 VPWR.n9 0.119
R71 VPWR.n13 VPWR.n11 0.119
R72 VPWR VPWR.n13 0.02
R73 VPB.t6 VPB.t4 559.345
R74 VPB.t2 VPB.t0 254.517
R75 VPB.t3 VPB.t2 254.517
R76 VPB.t1 VPB.t3 248.598
R77 VPB.t5 VPB.t1 248.598
R78 VPB.t4 VPB.t5 248.598
R79 VPB VPB.t6 192.367
R80 a_479_47.t0 a_479_47.t1 38.769
R81 A1.n0 A1.t0 212.079
R82 A1.n1 A1.t2 212.079
R83 A1.n0 A1.t3 139.779
R84 A1.n1 A1.t1 139.779
R85 A1 A1.n2 31.749
R86 A1.n2 A1.n1 28.034
R87 A1.n2 A1.n0 23.293
R88 B1_N.n0 B1_N.t0 253.682
R89 B1_N.n0 B1_N.t1 165.237
R90 B1_N B1_N.n0 39.598
R91 a_637_47.t0 a_637_47.t1 51.692
C0 A1 A2 0.36fF
C1 VGND Y 0.30fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__a21boi_4.ext - technology: sky130A

.subckt sky130_fd_sc_hd__a21boi_4 Y A1 B1_N A2 VGND VPWR VNB VPB
X0 a_223_297.t5 A2.t0 VPWR.t5 VPB.t5 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 Y.t3 A1.t0 a_658_47.t0 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 VPWR.t8 B1_N.t0 a_27_47.t0 VPB.t8 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 a_223_297.t6 A1.t1 VPWR.t6 VPB.t6 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 Y.t4 a_27_47.t2 VGND.t8 VNB.t5 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 VGND.t4 A2.t1 a_658_47.t7 VNB.t9 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 a_223_297.t10 a_27_47.t3 Y.t9 VPB.t11 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 Y.t10 a_27_47.t4 VGND.t7 VNB.t12 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 VPWR.t4 A2.t2 a_223_297.t4 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 a_658_47.t6 A2.t3 VGND.t3 VNB.t8 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 VPWR.t7 A1.t2 a_223_297.t7 VPB.t7 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 a_223_297.t0 A1.t3 VPWR.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 a_658_47.t5 A2.t4 VGND.t2 VNB.t7 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 Y.t11 a_27_47.t5 a_223_297.t11 VPB.t12 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14 a_223_297.t3 A2.t5 VPWR.t3 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 VPWR.t2 A2.t6 a_223_297.t2 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16 VPWR.t1 A1.t4 a_223_297.t1 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17 a_658_47.t3 A1.t5 Y.t2 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X18 VGND.t0 B1_N.t1 a_27_47.t1 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X19 a_223_297.t8 a_27_47.t6 Y.t5 VPB.t9 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X20 a_658_47.t2 A1.t6 Y.t1 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X21 VGND.t1 A2.t7 a_658_47.t4 VNB.t6 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X22 VGND.t6 a_27_47.t7 Y.t6 VNB.t10 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X23 VGND.t5 a_27_47.t8 Y.t7 VNB.t11 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X24 Y.t0 A1.t7 a_658_47.t1 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X25 Y.t8 a_27_47.t9 a_223_297.t9 VPB.t10 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
R0 A2.n3 A2.t6 236.179
R1 A2.n0 A2.t5 212.079
R2 A2.n5 A2.t2 212.079
R3 A2.n1 A2.t0 212.079
R4 A2.n4 A2.n3 204.185
R5 A2.n3 A2.t3 163.879
R6 A2.n0 A2.t1 139.779
R7 A2.n5 A2.t4 139.779
R8 A2.n1 A2.t7 139.779
R9 A2 A2.n0 88.013
R10 A2.n4 A2.n2 76
R11 A2.n7 A2.n6 76
R12 A2.n2 A2.n1 35.054
R13 A2.n6 A2.n5 21.909
R14 A2.n7 A2.n4 6.907
R15 A2 A2.n7 3.657
R16 VPWR.n24 VPWR.t8 575.112
R17 VPWR.n3 VPWR.n2 310.653
R18 VPWR.n1 VPWR.n0 306.463
R19 VPWR.n7 VPWR.n6 306.463
R20 VPWR.n12 VPWR.n11 306.463
R21 VPWR.n11 VPWR.t2 29.55
R22 VPWR.n2 VPWR.t3 27.58
R23 VPWR.n2 VPWR.t4 27.58
R24 VPWR.n0 VPWR.t5 27.58
R25 VPWR.n0 VPWR.t1 27.58
R26 VPWR.n6 VPWR.t0 27.58
R27 VPWR.n6 VPWR.t7 27.58
R28 VPWR.n11 VPWR.t6 27.58
R29 VPWR.n5 VPWR.n4 4.65
R30 VPWR.n8 VPWR.n7 4.65
R31 VPWR.n10 VPWR.n9 4.65
R32 VPWR.n13 VPWR.n12 4.65
R33 VPWR.n15 VPWR.n14 4.65
R34 VPWR.n17 VPWR.n16 4.65
R35 VPWR.n19 VPWR.n18 4.65
R36 VPWR.n21 VPWR.n20 4.65
R37 VPWR.n23 VPWR.n22 4.65
R38 VPWR.n25 VPWR.n24 4.084
R39 VPWR.n3 VPWR.n1 3.915
R40 VPWR.n5 VPWR.n3 0.328
R41 VPWR.n25 VPWR.n23 0.134
R42 VPWR VPWR.n25 0.127
R43 VPWR.n8 VPWR.n5 0.119
R44 VPWR.n10 VPWR.n8 0.119
R45 VPWR.n13 VPWR.n10 0.119
R46 VPWR.n15 VPWR.n13 0.119
R47 VPWR.n17 VPWR.n15 0.119
R48 VPWR.n19 VPWR.n17 0.119
R49 VPWR.n21 VPWR.n19 0.119
R50 VPWR.n23 VPWR.n21 0.119
R51 a_223_297.n9 a_223_297.n8 306.366
R52 a_223_297.n4 a_223_297.n3 292.5
R53 a_223_297.n5 a_223_297.n2 292.5
R54 a_223_297.n6 a_223_297.n1 292.5
R55 a_223_297.n8 a_223_297.t3 220.788
R56 a_223_297.n4 a_223_297.t11 219.988
R57 a_223_297.n7 a_223_297.n0 149.462
R58 a_223_297.n6 a_223_297.n5 54.785
R59 a_223_297.n7 a_223_297.n6 47.86
R60 a_223_297.n8 a_223_297.n7 47.582
R61 a_223_297.n5 a_223_297.n4 43.815
R62 a_223_297.n2 a_223_297.t10 33.49
R63 a_223_297.n0 a_223_297.t1 27.58
R64 a_223_297.n0 a_223_297.t0 27.58
R65 a_223_297.n1 a_223_297.t7 27.58
R66 a_223_297.n1 a_223_297.t6 27.58
R67 a_223_297.n2 a_223_297.t2 27.58
R68 a_223_297.n3 a_223_297.t9 27.58
R69 a_223_297.n3 a_223_297.t8 27.58
R70 a_223_297.n9 a_223_297.t4 27.58
R71 a_223_297.t5 a_223_297.n9 27.58
R72 VPB.t8 VPB.t12 562.305
R73 VPB.t11 VPB.t2 272.274
R74 VPB.t2 VPB.t6 260.436
R75 VPB.t4 VPB.t3 254.517
R76 VPB.t5 VPB.t4 254.517
R77 VPB.t1 VPB.t5 254.517
R78 VPB.t0 VPB.t1 254.517
R79 VPB.t7 VPB.t0 254.517
R80 VPB.t6 VPB.t7 254.517
R81 VPB.t10 VPB.t11 254.517
R82 VPB.t9 VPB.t10 254.517
R83 VPB.t12 VPB.t9 254.517
R84 VPB VPB.t8 213.084
R85 A1.n0 A1.t4 221.719
R86 A1.n7 A1.t3 221.719
R87 A1.n4 A1.t2 221.719
R88 A1.n2 A1.t1 221.719
R89 A1.n0 A1.t5 138.173
R90 A1.n7 A1.t7 138.173
R91 A1.n4 A1.t6 138.173
R92 A1.n2 A1.t0 138.173
R93 A1.n6 A1.n3 93.763
R94 A1 A1.n1 78.612
R95 A1.n9 A1.n8 76
R96 A1.n6 A1.n5 76
R97 A1.n1 A1.n0 22.124
R98 A1.n3 A1.n2 20.544
R99 A1.n9 A1.n6 17.763
R100 A1 A1.n9 15.151
R101 A1.n8 A1.n7 7.901
R102 A1.n5 A1.n4 6.321
R103 a_658_47.n5 a_658_47.n4 136.532
R104 a_658_47.n2 a_658_47.n0 105.66
R105 a_658_47.n4 a_658_47.n3 92.5
R106 a_658_47.n4 a_658_47.n2 46.468
R107 a_658_47.n2 a_658_47.n1 42.865
R108 a_658_47.n3 a_658_47.t1 25.846
R109 a_658_47.n3 a_658_47.t2 25.846
R110 a_658_47.n1 a_658_47.t4 25.846
R111 a_658_47.n1 a_658_47.t3 25.846
R112 a_658_47.n0 a_658_47.t7 25.846
R113 a_658_47.n0 a_658_47.t5 25.846
R114 a_658_47.t0 a_658_47.n5 25.846
R115 a_658_47.n5 a_658_47.t6 25.846
R116 Y Y.n9 314.544
R117 Y.n8 Y.n7 292.5
R118 Y.n2 Y.n0 142.536
R119 Y.n5 Y.n4 141.921
R120 Y.n6 Y.n2 93.191
R121 Y.n2 Y.n1 92.5
R122 Y.n6 Y.n5 53.04
R123 Y.n5 Y.n3 49.316
R124 Y.n9 Y.t5 27.58
R125 Y.n9 Y.t11 27.58
R126 Y.n7 Y.t9 27.58
R127 Y.n7 Y.t8 27.58
R128 Y.n3 Y.t6 25.846
R129 Y.n3 Y.t4 25.846
R130 Y.n4 Y.t7 25.846
R131 Y.n4 Y.t10 25.846
R132 Y.n0 Y.t2 25.846
R133 Y.n0 Y.t0 25.846
R134 Y.n1 Y.t1 25.846
R135 Y.n1 Y.t3 25.846
R136 Y.n8 Y.n6 24.481
R137 Y Y.n8 2.417
R138 VNB VNB.t0 6827.54
R139 VNB.t10 VNB.t8 3723.08
R140 VNB.t0 VNB.t12 2562.64
R141 VNB.t7 VNB.t9 2079.12
R142 VNB.t6 VNB.t7 2079.12
R143 VNB.t3 VNB.t6 2079.12
R144 VNB.t1 VNB.t3 2079.12
R145 VNB.t2 VNB.t1 2079.12
R146 VNB.t4 VNB.t2 2079.12
R147 VNB.t8 VNB.t4 2079.12
R148 VNB.t5 VNB.t10 2079.12
R149 VNB.t11 VNB.t5 2079.12
R150 VNB.t12 VNB.t11 2079.12
R151 B1_N.n0 B1_N.t0 241.534
R152 B1_N.n0 B1_N.t1 169.234
R153 B1_N B1_N.n0 85.955
R154 a_27_47.n0 a_27_47.t3 255.897
R155 a_27_47.t0 a_27_47.n13 242.708
R156 a_27_47.n1 a_27_47.t9 212.079
R157 a_27_47.n4 a_27_47.t6 212.079
R158 a_27_47.n8 a_27_47.t5 212.079
R159 a_27_47.n11 a_27_47.t4 148.542
R160 a_27_47.n13 a_27_47.t1 140.638
R161 a_27_47.n7 a_27_47.t8 139.779
R162 a_27_47.n3 a_27_47.t2 139.779
R163 a_27_47.n0 a_27_47.t7 139.779
R164 a_27_47.n6 a_27_47.n2 90.038
R165 a_27_47.n12 a_27_47.n11 76
R166 a_27_47.n6 a_27_47.n5 76
R167 a_27_47.n10 a_27_47.n9 76
R168 a_27_47.n1 a_27_47.n0 18.987
R169 a_27_47.n5 a_27_47.n3 17.527
R170 a_27_47.n9 a_27_47.n8 14.606
R171 a_27_47.n10 a_27_47.n6 14.038
R172 a_27_47.n12 a_27_47.n10 14.038
R173 a_27_47.n2 a_27_47.n1 11.684
R174 a_27_47.n13 a_27_47.n12 10.529
R175 a_27_47.n9 a_27_47.n7 4.381
R176 a_27_47.n5 a_27_47.n4 1.46
R177 VGND.n1 VGND.n0 119.447
R178 VGND.n2 VGND.t4 113.262
R179 VGND.n24 VGND.n23 106.463
R180 VGND.n14 VGND.n13 92.5
R181 VGND.n18 VGND.n17 92.5
R182 VGND.n30 VGND.n29 92.5
R183 VGND.n29 VGND.t0 36.923
R184 VGND.n29 VGND.t7 33.23
R185 VGND.n13 VGND.t3 25.846
R186 VGND.n17 VGND.t6 25.846
R187 VGND.n0 VGND.t2 25.846
R188 VGND.n0 VGND.t1 25.846
R189 VGND.n23 VGND.t8 25.846
R190 VGND.n23 VGND.t5 25.846
R191 VGND.n31 VGND.n30 10.752
R192 VGND.n2 VGND.n1 9.586
R193 VGND.n4 VGND.n3 4.65
R194 VGND.n6 VGND.n5 4.65
R195 VGND.n8 VGND.n7 4.65
R196 VGND.n10 VGND.n9 4.65
R197 VGND.n12 VGND.n11 4.65
R198 VGND.n16 VGND.n15 4.65
R199 VGND.n20 VGND.n19 4.65
R200 VGND.n22 VGND.n21 4.65
R201 VGND.n26 VGND.n25 4.65
R202 VGND.n28 VGND.n27 4.65
R203 VGND.n19 VGND.n18 2.727
R204 VGND.n25 VGND.n24 1.882
R205 VGND.n4 VGND.n2 0.33
R206 VGND.n15 VGND.n14 0.209
R207 VGND.n31 VGND.n28 0.132
R208 VGND VGND.n31 0.129
R209 VGND.n6 VGND.n4 0.119
R210 VGND.n8 VGND.n6 0.119
R211 VGND.n10 VGND.n8 0.119
R212 VGND.n12 VGND.n10 0.119
R213 VGND.n16 VGND.n12 0.119
R214 VGND.n20 VGND.n16 0.119
R215 VGND.n22 VGND.n20 0.119
R216 VGND.n26 VGND.n22 0.119
R217 VGND.n28 VGND.n26 0.119
C0 VPB VPWR 0.13fF
C1 Y A2 0.20fF
C2 A2 A1 0.55fF
C3 Y VGND 0.41fF
C4 VGND VPWR 0.15fF
C5 Y A1 0.24fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__a21o_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__a21o_1 A2 A1 B1 X VPWR VGND VNB VPB
X0 a_81_21.t1 B1.t0 VGND.t2 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 a_299_297.t2 B1.t1 a_81_21.t2 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 VPWR.t2 a_81_21.t3 X.t0 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 VPWR.t0 A1.t0 a_299_297.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 VGND.t0 a_81_21.t4 X.t1 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 VGND.t1 A2.t0 a_384_47.t1 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 a_299_297.t1 A2.t1 VPWR.t1 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 a_384_47.t0 A1.t1 a_81_21.t0 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
R0 B1.n0 B1.t1 230.791
R1 B1.n0 B1.t0 158.491
R2 B1 B1.n0 81.78
R3 VGND.n2 VGND.t1 145.987
R4 VGND.n1 VGND.n0 92.5
R5 VGND.n4 VGND.n3 92.5
R6 VGND.n0 VGND.t2 41.538
R7 VGND.n3 VGND.t0 41.538
R8 VGND.n5 VGND.n4 6.232
R9 VGND.n2 VGND.n1 4.744
R10 VGND.n5 VGND.n2 0.16
R11 VGND VGND.n5 0.127
R12 a_81_21.t2 a_81_21.n2 261.964
R13 a_81_21.n0 a_81_21.t3 230.791
R14 a_81_21.n2 a_81_21.n1 159.216
R15 a_81_21.n0 a_81_21.t4 158.491
R16 a_81_21.n2 a_81_21.n0 76
R17 a_81_21.n1 a_81_21.t0 25.846
R18 a_81_21.n1 a_81_21.t1 24.923
R19 VNB VNB.t2 6126.44
R20 VNB.t2 VNB.t3 4545.05
R21 VNB.t0 VNB.t1 2079.12
R22 VNB.t3 VNB.t0 2054.95
R23 a_299_297.n0 a_299_297.t1 426.358
R24 a_299_297.t0 a_299_297.n0 27.58
R25 a_299_297.n0 a_299_297.t2 26.595
R26 VPB.t2 VPB.t3 556.386
R27 VPB.t0 VPB.t1 254.517
R28 VPB.t3 VPB.t0 251.557
R29 VPB VPB.t2 198.286
R30 X.t0 X 467.164
R31 X.n0 X.t0 455.403
R32 X.n1 X.t1 117.423
R33 X X.n0 16
R34 X X.n1 10.092
R35 X.n1 X 6.646
R36 X.n0 X 0.738
R37 VPWR.n1 VPWR.t2 193.678
R38 VPWR.n1 VPWR.n0 167.199
R39 VPWR.n0 VPWR.t1 27.58
R40 VPWR.n0 VPWR.t0 27.58
R41 VPWR VPWR.n1 0.153
R42 A1.n0 A1.t0 241.534
R43 A1.n0 A1.t1 169.234
R44 A1 A1.n0 81.78
R45 A2.n0 A2.t1 231.014
R46 A2.n0 A2.t0 158.714
R47 A2 A2.n0 78.346
R48 a_384_47.t0 a_384_47.t1 51.692
C0 A1 VGND 0.10fF
C1 VPWR X 0.11fF
C2 A2 A1 0.10fF
C3 B1 A1 0.11fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__a21o_2.ext - technology: sky130A

.subckt sky130_fd_sc_hd__a21o_2 X B1 A1 A2 VGND VPWR VNB VPB
X0 VPWR.t2 a_80_199.t3 X.t3 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 X.t2 a_80_199.t4 VPWR.t1 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 VGND.t2 a_80_199.t5 X.t1 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 a_386_297.t1 A2.t0 VPWR.t3 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 X.t0 a_80_199.t6 VGND.t1 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 a_80_199.t2 B1.t0 VGND.t3 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 a_386_297.t2 B1.t1 a_80_199.t1 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 a_458_47.t0 A1.t0 a_80_199.t0 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 VPWR.t0 A1.t1 a_386_297.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 VGND.t0 A2.t1 a_458_47.t1 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
R0 a_80_199.n0 a_80_199.t4 324.545
R1 a_80_199.n2 a_80_199.t3 231.014
R2 a_80_199.t1 a_80_199.n4 215.323
R3 a_80_199.n4 a_80_199.n3 168.079
R4 a_80_199.n1 a_80_199.t5 148.386
R5 a_80_199.n0 a_80_199.t6 139.779
R6 a_80_199.n4 a_80_199.n2 76
R7 a_80_199.n3 a_80_199.t0 66.461
R8 a_80_199.n1 a_80_199.n0 59.446
R9 a_80_199.n3 a_80_199.t2 25.846
R10 a_80_199.n2 a_80_199.n1 10.328
R11 X.n2 X.n0 183.423
R12 X.n2 X.n1 144.587
R13 X.n1 X.t3 27.58
R14 X.n1 X.t2 27.58
R15 X.n0 X.t1 25.846
R16 X.n0 X.t0 25.846
R17 X X.n2 8.253
R18 VPWR.n1 VPWR.t2 571.144
R19 VPWR.n2 VPWR.n0 310.984
R20 VPWR.n5 VPWR.t1 195.868
R21 VPWR.n0 VPWR.t0 31.52
R22 VPWR.n0 VPWR.t3 30.535
R23 VPWR.n4 VPWR.n3 4.65
R24 VPWR.n6 VPWR.n5 4.65
R25 VPWR.n2 VPWR.n1 3.975
R26 VPWR.n4 VPWR.n2 0.147
R27 VPWR.n6 VPWR.n4 0.119
R28 VPWR VPWR.n6 0.02
R29 VPB.t3 VPB.t1 562.305
R30 VPB.t0 VPB.t4 275.233
R31 VPB.t1 VPB.t0 254.517
R32 VPB.t2 VPB.t3 254.517
R33 VPB VPB.t2 192.367
R34 VGND.n2 VGND.t0 193.072
R35 VGND.n5 VGND.t1 188.748
R36 VGND.n1 VGND.n0 106.463
R37 VGND.n0 VGND.t3 36.923
R38 VGND.n0 VGND.t2 25.846
R39 VGND.n6 VGND.n5 7.285
R40 VGND.n4 VGND.n3 4.65
R41 VGND.n2 VGND.n1 3.568
R42 VGND.n4 VGND.n2 0.152
R43 VGND.n6 VGND.n4 0.119
R44 VGND VGND.n6 0.02
R45 VNB VNB.t2 6940.96
R46 VNB.t4 VNB.t0 3142.86
R47 VNB.t0 VNB.t1 2562.64
R48 VNB.t3 VNB.t4 2369.23
R49 VNB.t2 VNB.t3 2079.12
R50 A2.n0 A2.t0 236.659
R51 A2.n0 A2.t1 183.826
R52 A2 A2.n0 78.234
R53 a_386_297.n0 a_386_297.t1 372.278
R54 a_386_297.t0 a_386_297.n0 27.58
R55 a_386_297.n0 a_386_297.t2 27.58
R56 B1.n0 B1.t1 230.154
R57 B1.n0 B1.t0 157.854
R58 B1 B1.n0 79.855
R59 A1.n0 A1.t1 236.932
R60 A1.n0 A1.t0 164.632
R61 A1 A1.n0 89.305
R62 a_458_47.t0 a_458_47.t1 70.153
C0 A1 A2 0.14fF
C1 X VPWR 0.17fF
C2 X VGND 0.11fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__a21o_4.ext - technology: sky130A

.subckt sky130_fd_sc_hd__a21o_4 A2 A1 X B1 VGND VPWR VNB VPB
X0 VGND.t3 B1.t0 a_84_21.t4 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 a_741_47.t0 A2.t0 VGND.t0 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 a_84_21.t5 A1.t0 a_741_47.t1 VNB.t9 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 VGND.t1 A2.t1 a_901_47.t0 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 VPWR.t7 a_84_21.t6 X.t7 VPB.t9 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 VPWR.t1 A2.t2 a_483_297.t1 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 a_483_297.t5 B1.t1 a_84_21.t3 VPB.t5 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 X.t3 a_84_21.t7 VGND.t4 VNB.t8 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 a_84_21.t2 B1.t2 a_483_297.t4 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 VGND.t7 a_84_21.t8 X.t2 VNB.t7 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 VPWR.t6 a_84_21.t9 X.t6 VPB.t8 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 a_483_297.t0 A2.t3 VPWR.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 VPWR.t3 A1.t1 a_483_297.t3 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13 VGND.t6 a_84_21.t10 X.t1 VNB.t6 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14 X.t5 a_84_21.t11 VPWR.t5 VPB.t7 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 a_84_21.t1 B1.t3 VGND.t2 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X16 a_483_297.t2 A1.t2 VPWR.t2 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17 X.t0 a_84_21.t12 VGND.t5 VNB.t5 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X18 a_901_47.t1 A1.t3 a_84_21.t0 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X19 X.t4 a_84_21.t13 VPWR.t4 VPB.t6 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
R0 B1.n0 B1.t1 212.079
R1 B1.n1 B1.t2 212.079
R2 B1.n0 B1.t0 139.779
R3 B1.n1 B1.t3 139.779
R4 B1 B1.n1 98.73
R5 B1.n1 B1.n0 61.345
R6 a_84_21.n13 a_84_21.n12 217.135
R7 a_84_21.n2 a_84_21.t6 212.079
R8 a_84_21.n6 a_84_21.t13 212.079
R9 a_84_21.n4 a_84_21.t9 212.079
R10 a_84_21.n3 a_84_21.t11 212.079
R11 a_84_21.n11 a_84_21.n1 179.262
R12 a_84_21.n2 a_84_21.t8 139.779
R13 a_84_21.n6 a_84_21.t12 139.779
R14 a_84_21.n4 a_84_21.t10 139.779
R15 a_84_21.n3 a_84_21.t7 139.779
R16 a_84_21.n12 a_84_21.n0 92.5
R17 a_84_21.n8 a_84_21.n5 89.187
R18 a_84_21.n9 a_84_21.n2 84.033
R19 a_84_21.n10 a_84_21.n9 83.518
R20 a_84_21.n8 a_84_21.n7 76
R21 a_84_21.n4 a_84_21.n3 62.806
R22 a_84_21.n5 a_84_21.n4 34.324
R23 a_84_21.n13 a_84_21.t3 26.595
R24 a_84_21.t2 a_84_21.n13 26.595
R25 a_84_21.n0 a_84_21.t4 24.923
R26 a_84_21.n0 a_84_21.t1 24.923
R27 a_84_21.n1 a_84_21.t0 24.923
R28 a_84_21.n1 a_84_21.t5 24.923
R29 a_84_21.n7 a_84_21.n6 21.178
R30 a_84_21.n9 a_84_21.n8 13.187
R31 a_84_21.n11 a_84_21.n10 4.141
R32 a_84_21.n12 a_84_21.n11 0.376
R33 VGND.n20 VGND.t4 190.262
R34 VGND.n2 VGND.t1 112.546
R35 VGND.n1 VGND.n0 106.463
R36 VGND.n16 VGND.n15 106.463
R37 VGND.n6 VGND.n5 92.5
R38 VGND.n10 VGND.n9 92.5
R39 VGND.n9 VGND.t7 46.153
R40 VGND.n0 VGND.t3 32.307
R41 VGND.n5 VGND.t2 28.615
R42 VGND.n15 VGND.t5 25.846
R43 VGND.n15 VGND.t6 25.846
R44 VGND.n0 VGND.t0 24.923
R45 VGND.n21 VGND.n20 4.65
R46 VGND.n4 VGND.n3 4.65
R47 VGND.n8 VGND.n7 4.65
R48 VGND.n12 VGND.n11 4.65
R49 VGND.n14 VGND.n13 4.65
R50 VGND.n17 VGND.n16 4.65
R51 VGND.n19 VGND.n18 4.65
R52 VGND.n2 VGND.n1 3.981
R53 VGND.n11 VGND.n10 0.966
R54 VGND.n7 VGND.n6 0.241
R55 VGND.n4 VGND.n2 0.141
R56 VGND.n8 VGND.n4 0.119
R57 VGND.n12 VGND.n8 0.119
R58 VGND.n14 VGND.n12 0.119
R59 VGND.n17 VGND.n14 0.119
R60 VGND.n19 VGND.n17 0.119
R61 VGND.n21 VGND.n19 0.119
R62 VGND VGND.n21 0.022
R63 VNB VNB.t8 6198.96
R64 VNB.t7 VNB.t3 4665.93
R65 VNB.t4 VNB.t1 2224.18
R66 VNB.t5 VNB.t7 2079.12
R67 VNB.t6 VNB.t5 2079.12
R68 VNB.t8 VNB.t6 2079.12
R69 VNB.t0 VNB.t2 2030.77
R70 VNB.t9 VNB.t0 2030.77
R71 VNB.t3 VNB.t4 2030.77
R72 VNB.t1 VNB.t9 1837.36
R73 A2.n1 A2.t3 241.534
R74 A2.n0 A2.t2 241.534
R75 A2 A2.n0 178.976
R76 A2.n1 A2.t1 169.234
R77 A2.n0 A2.t0 169.234
R78 A2 A2.n1 90.592
R79 a_741_47.t0 a_741_47.t1 42.461
R80 A1.n0 A1.t1 212.079
R81 A1.n1 A1.t2 212.079
R82 A1.n0 A1.t3 139.779
R83 A1.n1 A1.t0 139.779
R84 A1 A1.n2 81.554
R85 A1.n2 A1.n0 35.054
R86 A1.n2 A1.n1 26.29
R87 a_901_47.t0 a_901_47.t1 49.846
R88 X.n2 X.n0 208.95
R89 X.n5 X.n3 157.252
R90 X.n2 X.n1 151.074
R91 X.n5 X.n4 92.5
R92 X.n1 X.t6 27.58
R93 X.n1 X.t5 27.58
R94 X.n0 X.t7 27.58
R95 X.n0 X.t4 27.58
R96 X.n4 X.t1 25.846
R97 X.n4 X.t3 25.846
R98 X.n3 X.t2 25.846
R99 X.n3 X.t0 25.846
R100 X X.n5 25.684
R101 X.n6 X.n2 24.47
R102 X X.n6 18.07
R103 X.n6 X 3.694
R104 VPWR.n3 VPWR.n0 310.449
R105 VPWR.n2 VPWR.n1 306.463
R106 VPWR.n19 VPWR.t5 191.018
R107 VPWR.n15 VPWR.n14 163.438
R108 VPWR.n10 VPWR.t7 152.677
R109 VPWR.n14 VPWR.t4 27.58
R110 VPWR.n14 VPWR.t6 27.58
R111 VPWR.n1 VPWR.t2 26.595
R112 VPWR.n1 VPWR.t1 26.595
R113 VPWR.n0 VPWR.t0 26.595
R114 VPWR.n0 VPWR.t3 26.595
R115 VPWR.n5 VPWR.n4 4.65
R116 VPWR.n7 VPWR.n6 4.65
R117 VPWR.n9 VPWR.n8 4.65
R118 VPWR.n11 VPWR.n10 4.65
R119 VPWR.n13 VPWR.n12 4.65
R120 VPWR.n16 VPWR.n15 4.65
R121 VPWR.n18 VPWR.n17 4.65
R122 VPWR.n20 VPWR.n19 4.65
R123 VPWR.n3 VPWR.n2 3.895
R124 VPWR.n5 VPWR.n3 0.317
R125 VPWR.n7 VPWR.n5 0.119
R126 VPWR.n9 VPWR.n7 0.119
R127 VPWR.n11 VPWR.n9 0.119
R128 VPWR.n13 VPWR.n11 0.119
R129 VPWR.n16 VPWR.n13 0.119
R130 VPWR.n18 VPWR.n16 0.119
R131 VPWR.n20 VPWR.n18 0.119
R132 VPWR VPWR.n20 0.022
R133 VPB.t9 VPB.t4 571.183
R134 VPB.t6 VPB.t9 254.517
R135 VPB.t8 VPB.t6 254.517
R136 VPB.t7 VPB.t8 254.517
R137 VPB.t3 VPB.t0 248.598
R138 VPB.t2 VPB.t3 248.598
R139 VPB.t1 VPB.t2 248.598
R140 VPB.t5 VPB.t1 248.598
R141 VPB.t4 VPB.t5 248.598
R142 VPB VPB.t7 207.165
R143 a_483_297.n2 a_483_297.t4 268.803
R144 a_483_297.n1 a_483_297.t0 215.302
R145 a_483_297.n1 a_483_297.n0 151.337
R146 a_483_297.n3 a_483_297.n2 149.708
R147 a_483_297.n2 a_483_297.n1 61.216
R148 a_483_297.n0 a_483_297.t3 26.595
R149 a_483_297.n0 a_483_297.t2 26.595
R150 a_483_297.t1 a_483_297.n3 26.595
R151 a_483_297.n3 a_483_297.t5 26.595
C0 X VGND 0.18fF
C1 VPWR VGND 0.13fF
C2 VPWR X 0.39fF
C3 A2 A1 0.30fF
C4 VPWR VPB 0.11fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__a21oi_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__a21oi_1 A1 B1 Y A2 VPWR VGND VNB VPB
X0 a_199_47.t0 A1.t0 Y.t1 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 a_113_297.t1 A2.t0 VPWR.t1 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 Y.t0 B1.t0 VGND.t0 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 VPWR.t0 A1.t1 a_113_297.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 a_113_297.t2 B1.t1 Y.t2 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 VGND.t1 A2.t1 a_199_47.t1 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
R0 A1.n0 A1.t1 241.534
R1 A1.n0 A1.t0 169.234
R2 A1 A1.n0 80.654
R3 Y.n0 Y.t2 211.964
R4 Y Y.n1 177.787
R5 Y.n1 Y.t1 25.846
R6 Y.n1 Y.t0 25.846
R7 Y Y.n0 8.226
R8 Y.n0 Y 7.354
R9 a_199_47.t0 a_199_47.t1 54.461
R10 VNB VNB.t0 6174.79
R11 VNB.t1 VNB.t2 2151.65
R12 VNB.t0 VNB.t1 2079.12
R13 A2.n0 A2.t0 231.014
R14 A2.n0 A2.t1 158.714
R15 A2 A2.n0 78.386
R16 VPWR VPWR.n0 319.958
R17 VPWR.n0 VPWR.t1 30.535
R18 VPWR.n0 VPWR.t0 27.58
R19 a_113_297.n0 a_113_297.t1 294.857
R20 a_113_297.t0 a_113_297.n0 27.58
R21 a_113_297.n0 a_113_297.t2 27.58
R22 VPB.t0 VPB.t1 263.395
R23 VPB.t2 VPB.t0 254.517
R24 VPB VPB.t2 204.205
R25 B1.n0 B1.t1 229.368
R26 B1.n0 B1.t0 157.068
R27 B1 B1.n0 78.933
R28 VGND.n0 VGND.t0 192.584
R29 VGND.n0 VGND.t1 145.199
R30 VGND VGND.n0 0.057
C0 A2 A1 0.11fF
C1 VGND A1 0.10fF
C2 Y B1 0.14fF
C3 Y A1 0.11fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__a21oi_2.ext - technology: sky130A

.subckt sky130_fd_sc_hd__a21oi_2 B1 A2 A1 Y VGND VPWR VNB VPB
X0 VGND.t2 A2.t0 a_285_47.t1 VNB.t5 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 VGND.t1 B1.t0 Y.t3 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 Y.t1 A1.t0 a_114_47.t0 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 a_114_47.t1 A2.t1 VGND.t3 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 a_27_297.t3 B1.t1 Y.t5 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 a_27_297.t1 A1.t1 VPWR.t1 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 Y.t4 B1.t2 a_27_297.t2 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 VPWR.t3 A2.t2 a_27_297.t4 VPB.t5 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 a_27_297.t5 A2.t3 VPWR.t2 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 VPWR.t0 A1.t2 a_27_297.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 a_285_47.t0 A1.t3 Y.t0 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 Y.t2 B1.t3 VGND.t0 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
R0 A2.n1 A2.t2 671.729
R1 A2.n0 A2.t3 241.534
R2 A2.n0 A2.t0 169.234
R3 A2.n1 A2.t1 167.068
R4 A2.n2 A2.n0 165.904
R5 A2.n2 A2.n1 76
R6 A2 A2.n2 5.1
R7 a_285_47.t0 a_285_47.t1 38.769
R8 VGND.n2 VGND.t1 119.005
R9 VGND.n1 VGND.n0 106.463
R10 VGND.n9 VGND.t3 91.133
R11 VGND.n0 VGND.t0 35.076
R12 VGND.n0 VGND.t2 25.846
R13 VGND.n10 VGND.n9 4.65
R14 VGND.n4 VGND.n3 4.65
R15 VGND.n6 VGND.n5 4.65
R16 VGND.n8 VGND.n7 4.65
R17 VGND.n2 VGND.n1 4.036
R18 VGND.n4 VGND.n2 0.217
R19 VGND.n6 VGND.n4 0.119
R20 VGND.n8 VGND.n6 0.119
R21 VGND.n10 VGND.n8 0.119
R22 VGND VGND.n10 0.022
R23 VNB VNB.t4 6198.96
R24 VNB.t5 VNB.t0 2320.88
R25 VNB.t2 VNB.t1 2079.12
R26 VNB.t4 VNB.t2 2054.95
R27 VNB.t0 VNB.t3 2030.77
R28 VNB.t1 VNB.t5 1740.66
R29 B1.n1 B1.t1 218.506
R30 B1.n0 B1.t2 218.506
R31 B1.n1 B1.t0 146.206
R32 B1.n0 B1.t3 146.206
R33 B1.n2 B1.n1 132.51
R34 B1.n1 B1.n0 69.806
R35 B1.n2 B1 13.265
R36 B1 B1.n2 2.56
R37 Y.n2 Y.n1 185.99
R38 Y.n3 Y.n0 124.12
R39 Y Y.n4 92.7
R40 Y.n1 Y.t5 26.595
R41 Y.n1 Y.t4 26.595
R42 Y.n0 Y.t0 25.846
R43 Y.n0 Y.t1 25.846
R44 Y.n4 Y.t3 24.923
R45 Y.n4 Y.t2 24.923
R46 Y Y.n3 11
R47 Y.n3 Y.n2 2.4
R48 A1.n0 A1.t2 212.079
R49 A1.n1 A1.t1 212.079
R50 A1.n0 A1.t3 139.779
R51 A1.n1 A1.t0 139.779
R52 A1 A1.n2 31.731
R53 A1.n2 A1.n0 28.347
R54 A1.n2 A1.n1 22.979
R55 a_114_47.t0 a_114_47.t1 50.769
R56 a_27_297.t3 a_27_297.n3 251.715
R57 a_27_297.n1 a_27_297.t4 217.093
R58 a_27_297.n1 a_27_297.n0 149.831
R59 a_27_297.n3 a_27_297.n2 143.026
R60 a_27_297.n3 a_27_297.n1 58.704
R61 a_27_297.n0 a_27_297.t0 27.58
R62 a_27_297.n0 a_27_297.t1 27.58
R63 a_27_297.n2 a_27_297.t2 26.595
R64 a_27_297.n2 a_27_297.t5 26.595
R65 VPB.t1 VPB.t0 254.517
R66 VPB.t5 VPB.t1 254.517
R67 VPB.t2 VPB.t3 248.598
R68 VPB.t4 VPB.t2 248.598
R69 VPB.t0 VPB.t4 248.598
R70 VPB VPB.t5 204.205
R71 VPWR.n2 VPWR.n0 319.729
R72 VPWR.n2 VPWR.n1 309.764
R73 VPWR.n1 VPWR.t1 27.58
R74 VPWR.n1 VPWR.t3 27.58
R75 VPWR.n0 VPWR.t2 26.595
R76 VPWR.n0 VPWR.t0 26.595
R77 VPWR VPWR.n2 0.259
C0 B1 Y 0.12fF
C1 VGND Y 0.33fF
C2 A1 A2 0.36fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__a21oi_4.ext - technology: sky130A

.subckt sky130_fd_sc_hd__a21oi_4 B1 A2 A1 Y VGND VPWR VNB VPB
X0 a_28_297.t3 B1.t0 Y.t7 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_462_47.t4 A1.t0 Y.t8 VNB.t8 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 Y.t6 B1.t1 a_28_297.t2 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 Y.t3 B1.t2 VGND.t3 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 a_462_47.t3 A1.t1 Y.t9 VNB.t7 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 a_28_297.t7 A2.t0 VPWR.t7 VPB.t7 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 a_462_47.t5 A2.t1 VGND.t5 VNB.t9 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 Y.t5 B1.t3 a_28_297.t1 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 VGND.t2 B1.t4 Y.t2 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 VGND.t1 B1.t5 Y.t1 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 Y.t10 A1.t2 a_462_47.t2 VNB.t6 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 a_28_297.t8 A1.t3 VPWR.t3 VPB.t8 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 VPWR.t6 A2.t2 a_28_297.t6 VPB.t6 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13 Y.t0 B1.t6 VGND.t0 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14 VGND.t4 A2.t3 a_462_47.t0 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X15 a_28_297.t0 B1.t7 Y.t4 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16 VPWR.t2 A1.t4 a_28_297.t9 VPB.t9 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17 a_28_297.t10 A1.t5 VPWR.t1 VPB.t10 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X18 VGND.t6 A2.t4 a_462_47.t6 VNB.t10 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X19 VPWR.t5 A2.t5 a_28_297.t4 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X20 a_28_297.t5 A2.t6 VPWR.t4 VPB.t5 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X21 Y.t11 A1.t6 a_462_47.t1 VNB.t5 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X22 a_462_47.t7 A2.t7 VGND.t7 VNB.t11 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X23 VPWR.t0 A1.t7 a_28_297.t11 VPB.t11 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
R0 B1.n0 B1.t7 212.079
R1 B1.n1 B1.t3 212.079
R2 B1.n5 B1.t0 212.079
R3 B1.n3 B1.t1 212.079
R4 B1.n0 B1.t4 139.779
R5 B1.n1 B1.t2 139.779
R6 B1.n5 B1.t5 139.779
R7 B1.n3 B1.t6 139.779
R8 B1 B1.n2 82.568
R9 B1.n7 B1.n6 76
R10 B1.n1 B1.n0 62.806
R11 B1.n7 B1.n4 54.62
R12 B1.n2 B1.n1 10.224
R13 B1.n4 B1.n3 9.126
R14 B1 B1.n7 4.884
R15 B1.n6 B1.n5 2.921
R16 Y Y.n12 316.393
R17 Y.n11 Y.n10 292.5
R18 Y.n2 Y.n0 142.536
R19 Y.n6 Y.n5 140.641
R20 Y.n9 Y.n2 93.191
R21 Y.n2 Y.n1 92.5
R22 Y.n7 Y.n3 92.5
R23 Y.n9 Y.n8 31.779
R24 Y.n12 Y.t7 27.58
R25 Y.n12 Y.t6 27.58
R26 Y.n10 Y.t4 27.58
R27 Y.n10 Y.t5 27.58
R28 Y.n0 Y.t8 25.846
R29 Y.n0 Y.t11 25.846
R30 Y.n1 Y.t9 25.846
R31 Y.n1 Y.t10 25.846
R32 Y.n5 Y.t1 25.846
R33 Y.n5 Y.t0 25.846
R34 Y.n3 Y.t2 25.846
R35 Y.n3 Y.t3 25.846
R36 Y.n11 Y.n9 25.416
R37 Y.n6 Y.n4 15.889
R38 Y.n8 Y.n7 2.56
R39 Y.n7 Y.n6 1.28
R40 Y Y.n11 0.568
R41 a_28_297.n1 a_28_297.n0 306.366
R42 a_28_297.n7 a_28_297.n6 292.5
R43 a_28_297.n9 a_28_297.n8 292.5
R44 a_28_297.n1 a_28_297.t5 220.788
R45 a_28_297.n8 a_28_297.t2 219.988
R46 a_28_297.n5 a_28_297.n4 149.462
R47 a_28_297.n3 a_28_297.n2 149.462
R48 a_28_297.n7 a_28_297.n5 54.785
R49 a_28_297.n5 a_28_297.n3 47.86
R50 a_28_297.n3 a_28_297.n1 47.582
R51 a_28_297.n8 a_28_297.n7 43.815
R52 a_28_297.n6 a_28_297.t0 33.49
R53 a_28_297.n6 a_28_297.t4 27.58
R54 a_28_297.n2 a_28_297.t11 27.58
R55 a_28_297.n2 a_28_297.t10 27.58
R56 a_28_297.n4 a_28_297.t9 27.58
R57 a_28_297.n4 a_28_297.t8 27.58
R58 a_28_297.n0 a_28_297.t6 27.58
R59 a_28_297.n0 a_28_297.t7 27.58
R60 a_28_297.n9 a_28_297.t1 27.58
R61 a_28_297.t3 a_28_297.n9 27.58
R62 VPB.t0 VPB.t4 272.274
R63 VPB.t4 VPB.t8 260.436
R64 VPB.t6 VPB.t5 254.517
R65 VPB.t7 VPB.t6 254.517
R66 VPB.t11 VPB.t7 254.517
R67 VPB.t10 VPB.t11 254.517
R68 VPB.t9 VPB.t10 254.517
R69 VPB.t8 VPB.t9 254.517
R70 VPB.t1 VPB.t0 254.517
R71 VPB.t3 VPB.t1 254.517
R72 VPB.t2 VPB.t3 254.517
R73 VPB VPB.t2 192.367
R74 A1.n0 A1.t7 221.719
R75 A1.n7 A1.t5 221.719
R76 A1.n4 A1.t4 221.719
R77 A1.n2 A1.t3 221.719
R78 A1.n0 A1.t0 138.173
R79 A1.n7 A1.t6 138.173
R80 A1.n4 A1.t1 138.173
R81 A1.n2 A1.t2 138.173
R82 A1.n6 A1.n3 93.763
R83 A1.n10 A1.n1 76
R84 A1.n9 A1.n8 76
R85 A1.n6 A1.n5 76
R86 A1.n1 A1.n0 22.124
R87 A1.n3 A1.n2 20.544
R88 A1.n10 A1.n9 17.763
R89 A1.n9 A1.n6 17.763
R90 A1.n8 A1.n7 7.901
R91 A1.n5 A1.n4 6.321
R92 A1 A1.n10 0.783
R93 a_462_47.n3 a_462_47.n2 136.532
R94 a_462_47.n4 a_462_47.n0 105.66
R95 a_462_47.n3 a_462_47.n1 92.5
R96 a_462_47.n4 a_462_47.n3 46.468
R97 a_462_47.n5 a_462_47.n4 42.865
R98 a_462_47.n2 a_462_47.t2 25.846
R99 a_462_47.n2 a_462_47.t5 25.846
R100 a_462_47.n1 a_462_47.t1 25.846
R101 a_462_47.n1 a_462_47.t3 25.846
R102 a_462_47.n0 a_462_47.t0 25.846
R103 a_462_47.n0 a_462_47.t7 25.846
R104 a_462_47.n5 a_462_47.t6 25.846
R105 a_462_47.t4 a_462_47.n5 25.846
R106 VNB VNB.t0 6078.09
R107 VNB.t2 VNB.t9 2272.53
R108 VNB.t11 VNB.t4 2079.12
R109 VNB.t10 VNB.t11 2079.12
R110 VNB.t8 VNB.t10 2079.12
R111 VNB.t5 VNB.t8 2079.12
R112 VNB.t7 VNB.t5 2079.12
R113 VNB.t6 VNB.t7 2079.12
R114 VNB.t9 VNB.t6 2079.12
R115 VNB.t3 VNB.t2 2079.12
R116 VNB.t1 VNB.t3 2079.12
R117 VNB.t0 VNB.t1 2079.12
R118 VGND.n1 VGND.n0 119.447
R119 VGND.n2 VGND.t4 113.192
R120 VGND.n14 VGND.n13 108.957
R121 VGND.n19 VGND.n18 106.463
R122 VGND.n23 VGND.t0 102.497
R123 VGND.n13 VGND.t2 33.23
R124 VGND.n0 VGND.t7 25.846
R125 VGND.n0 VGND.t6 25.846
R126 VGND.n13 VGND.t5 25.846
R127 VGND.n18 VGND.t3 25.846
R128 VGND.n18 VGND.t1 25.846
R129 VGND.n2 VGND.n1 14.011
R130 VGND.n24 VGND.n23 4.65
R131 VGND.n4 VGND.n3 4.65
R132 VGND.n6 VGND.n5 4.65
R133 VGND.n8 VGND.n7 4.65
R134 VGND.n10 VGND.n9 4.65
R135 VGND.n12 VGND.n11 4.65
R136 VGND.n15 VGND.n14 4.65
R137 VGND.n17 VGND.n16 4.65
R138 VGND.n20 VGND.n19 4.65
R139 VGND.n22 VGND.n21 4.65
R140 VGND.n4 VGND.n2 0.423
R141 VGND.n6 VGND.n4 0.119
R142 VGND.n8 VGND.n6 0.119
R143 VGND.n10 VGND.n8 0.119
R144 VGND.n12 VGND.n10 0.119
R145 VGND.n15 VGND.n12 0.119
R146 VGND.n17 VGND.n15 0.119
R147 VGND.n20 VGND.n17 0.119
R148 VGND.n22 VGND.n20 0.119
R149 VGND.n24 VGND.n22 0.119
R150 VGND VGND.n24 0.02
R151 A2.n3 A2.t5 236.179
R152 A2.n0 A2.t6 212.079
R153 A2.n5 A2.t2 212.079
R154 A2.n1 A2.t0 212.079
R155 A2.n4 A2.n3 204.185
R156 A2.n3 A2.t1 163.879
R157 A2.n0 A2.t3 139.779
R158 A2.n5 A2.t7 139.779
R159 A2.n1 A2.t4 139.779
R160 A2 A2.n0 86.693
R161 A2.n4 A2.n2 76
R162 A2.n7 A2.n6 76
R163 A2.n2 A2.n1 35.054
R164 A2.n6 A2.n5 21.909
R165 A2.n7 A2.n4 6.907
R166 A2 A2.n7 4.977
R167 VPWR.n3 VPWR.n2 310.509
R168 VPWR.n1 VPWR.n0 306.463
R169 VPWR.n7 VPWR.n6 306.463
R170 VPWR.n12 VPWR.n11 306.463
R171 VPWR.n11 VPWR.t5 29.55
R172 VPWR.n2 VPWR.t4 27.58
R173 VPWR.n2 VPWR.t6 27.58
R174 VPWR.n0 VPWR.t7 27.58
R175 VPWR.n0 VPWR.t0 27.58
R176 VPWR.n6 VPWR.t1 27.58
R177 VPWR.n6 VPWR.t2 27.58
R178 VPWR.n11 VPWR.t3 27.58
R179 VPWR.n3 VPWR.n1 6.461
R180 VPWR.n5 VPWR.n4 4.65
R181 VPWR.n8 VPWR.n7 4.65
R182 VPWR.n10 VPWR.n9 4.65
R183 VPWR.n13 VPWR.n12 3.765
R184 VPWR VPWR.n13 0.592
R185 VPWR.n5 VPWR.n3 0.441
R186 VPWR.n13 VPWR.n10 0.144
R187 VPWR.n8 VPWR.n5 0.119
R188 VPWR.n10 VPWR.n8 0.119
C0 VPWR VGND 0.13fF
C1 Y A1 0.24fF
C2 A2 A1 0.55fF
C3 VPB VPWR 0.11fF
C4 B1 Y 0.37fF
C5 Y VGND 0.36fF
C6 Y A2 0.20fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__a22o_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__a22o_1 A1 A2 X B2 B1 VPWR VGND VNB VPB
X0 VPWR.t0 A2.t0 a_109_297.t1 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_27_297.t1 B1.t0 a_109_47.t1 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 VGND.t1 A2.t1 a_373_47.t0 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 X.t1 a_27_297.t4 VPWR.t1 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 a_27_297.t2 B1.t1 a_109_297.t3 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 a_109_297.t2 A1.t0 VPWR.t2 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 a_373_47.t1 A1.t1 a_27_297.t3 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 X.t0 a_27_297.t5 VGND.t2 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 a_109_297.t0 B2.t0 a_27_297.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 a_109_47.t0 B2.t1 VGND.t0 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
R0 A2.n0 A2.t0 722.091
R1 A2.n0 A2.t1 162.961
R2 A2 A2.n0 86.281
R3 a_109_297.n1 a_109_297.n0 521.274
R4 a_109_297.n0 a_109_297.t1 34.475
R5 a_109_297.n0 a_109_297.t2 28.565
R6 a_109_297.n1 a_109_297.t3 26.595
R7 a_109_297.t0 a_109_297.n1 26.595
R8 VPWR.n1 VPWR.t2 500.492
R9 VPWR.n1 VPWR.n0 172.583
R10 VPWR.n0 VPWR.t0 34.475
R11 VPWR.n0 VPWR.t1 26.595
R12 VPWR VPWR.n1 0.445
R13 VPB.t4 VPB.t3 550.467
R14 VPB.t3 VPB.t1 278.193
R15 VPB.t1 VPB.t2 272.274
R16 VPB.t0 VPB.t4 248.598
R17 VPB VPB.t0 192.367
R18 B1.n0 B1.t1 239.503
R19 B1.n0 B1.t0 167.203
R20 B1 B1.n0 85.848
R21 a_109_47.t0 a_109_47.t1 42.461
R22 a_27_297.n3 a_27_297.t2 481.625
R23 a_27_297.n1 a_27_297.t4 233.573
R24 a_27_297.n0 a_27_297.t1 207.271
R25 a_27_297.t0 a_27_297.n3 191.658
R26 a_27_297.n0 a_27_297.t3 175.576
R27 a_27_297.n1 a_27_297.t5 161.273
R28 a_27_297.n3 a_27_297.n2 139.822
R29 a_27_297.n2 a_27_297.n0 106.151
R30 a_27_297.n2 a_27_297.n1 76.89
R31 VNB VNB.t0 6078.09
R32 VNB.t1 VNB.t3 4545.05
R33 VNB.t3 VNB.t2 2417.58
R34 VNB.t2 VNB.t4 2224.18
R35 VNB.t0 VNB.t1 1837.36
R36 a_373_47.t0 a_373_47.t1 64.615
R37 VGND.n1 VGND.n0 110.445
R38 VGND.n1 VGND.t0 102.402
R39 VGND.n0 VGND.t1 32.307
R40 VGND.n0 VGND.t2 24.923
R41 VGND VGND.n1 0.054
R42 X X.t0 255.59
R43 X.n0 X.t1 172.965
R44 X X.n0 12.564
R45 X.n0 X 4.065
R46 A1.n0 A1.t0 256.714
R47 A1.n0 A1.t1 161.273
R48 A1.n1 A1.n0 79.657
R49 A1 A1.n1 18.895
R50 A1.n1 A1 3.961
R51 B2.n0 B2.t0 241.534
R52 B2.n0 B2.t1 169.234
R53 B2 B2.n0 92.64
C0 X VPWR 0.12fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__a22o_2.ext - technology: sky130A

.subckt sky130_fd_sc_hd__a22o_2 A1 A2 X B2 B1 VPWR VGND VNB VPB
X0 VPWR.t1 a_27_297.t4 X.t3 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 VGND.t3 A2.t0 a_381_47.t1 VNB.t5 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 X.t1 a_27_297.t5 VGND.t2 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 X.t2 a_27_297.t6 VPWR.t0 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 a_27_297.t0 B1.t0 a_109_47.t1 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 a_27_297.t1 B1.t1 a_109_297.t2 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 VGND.t1 a_27_297.t7 X.t0 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 a_109_297.t1 A1.t0 VPWR.t2 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 VPWR.t3 A2.t1 a_109_297.t0 VPB.t5 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 a_381_47.t0 A1.t1 a_27_297.t2 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 a_109_297.t3 B2.t0 a_27_297.t3 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 a_109_47.t0 B2.t1 VGND.t0 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
R0 a_27_297.t1 a_27_297.n4 624.107
R1 a_27_297.n4 a_27_297.n3 213.036
R2 a_27_297.n0 a_27_297.t4 212.079
R3 a_27_297.n1 a_27_297.t6 212.079
R4 a_27_297.n2 a_27_297.t0 185.787
R5 a_27_297.n2 a_27_297.t2 157.115
R6 a_27_297.n0 a_27_297.t7 139.779
R7 a_27_297.n1 a_27_297.t5 139.779
R8 a_27_297.n4 a_27_297.t3 118.508
R9 a_27_297.n3 a_27_297.n2 109.492
R10 a_27_297.n3 a_27_297.n1 82.572
R11 a_27_297.n1 a_27_297.n0 61.345
R12 X X.n0 190.975
R13 X.n2 X.n1 146.37
R14 X.n1 X.t3 26.595
R15 X.n1 X.t2 26.595
R16 X.n0 X.t0 24.923
R17 X.n0 X.t1 24.923
R18 X X.n2 12.564
R19 X.n2 X 4.065
R20 VPWR.n5 VPWR.t2 546.316
R21 VPWR.n2 VPWR.t1 169.794
R22 VPWR.n1 VPWR.n0 165.765
R23 VPWR.n0 VPWR.t3 35.46
R24 VPWR.n0 VPWR.t0 26.595
R25 VPWR.n4 VPWR.n3 4.65
R26 VPWR.n6 VPWR.n5 3.953
R27 VPWR.n2 VPWR.n1 3.745
R28 VPWR VPWR.n6 0.359
R29 VPWR.n4 VPWR.n2 0.267
R30 VPWR.n6 VPWR.n4 0.139
R31 VPB.t0 VPB.t3 556.386
R32 VPB.t3 VPB.t5 284.112
R33 VPB.t5 VPB.t1 275.233
R34 VPB.t1 VPB.t2 248.598
R35 VPB.t4 VPB.t0 248.598
R36 VPB VPB.t4 189.408
R37 A2.n0 A2.t1 241.534
R38 A2.n0 A2.t0 169.234
R39 A2 A2.n0 91.36
R40 a_381_47.t0 a_381_47.t1 60.923
R41 VGND.n2 VGND.t1 119.449
R42 VGND.n1 VGND.n0 108.015
R43 VGND.n11 VGND.t0 99.022
R44 VGND.n0 VGND.t2 33.23
R45 VGND.n0 VGND.t3 24.923
R46 VGND.n12 VGND.n11 4.65
R47 VGND.n4 VGND.n3 4.65
R48 VGND.n6 VGND.n5 4.65
R49 VGND.n8 VGND.n7 4.65
R50 VGND.n10 VGND.n9 4.65
R51 VGND.n2 VGND.n1 3.841
R52 VGND.n4 VGND.n2 0.251
R53 VGND.n6 VGND.n4 0.119
R54 VGND.n8 VGND.n6 0.119
R55 VGND.n10 VGND.n8 0.119
R56 VGND.n12 VGND.n10 0.119
R57 VGND VGND.n12 0.02
R58 VNB VNB.t0 6053.91
R59 VNB.t1 VNB.t2 4738.46
R60 VNB.t2 VNB.t5 2320.88
R61 VNB.t5 VNB.t4 2248.35
R62 VNB.t4 VNB.t3 2030.77
R63 VNB.t0 VNB.t1 1837.36
R64 B1.n0 B1.t1 239.503
R65 B1.n0 B1.t0 167.203
R66 B1 B1.n0 85.848
R67 a_109_47.t0 a_109_47.t1 42.461
R68 a_109_297.n1 a_109_297.n0 514.222
R69 a_109_297.t0 a_109_297.n1 33.49
R70 a_109_297.n1 a_109_297.t1 31.52
R71 a_109_297.n0 a_109_297.t2 26.595
R72 a_109_297.n0 a_109_297.t3 26.595
R73 A1.n0 A1.t0 233.868
R74 A1.n0 A1.t1 161.568
R75 A1.n1 A1.n0 79.657
R76 A1 A1.n1 18.895
R77 A1.n1 A1 3.961
R78 B2.n0 B2.t0 241.534
R79 B2.n0 B2.t1 169.234
R80 B2 B2.n0 92.64
C0 X VGND 0.18fF
C1 X VPWR 0.30fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__a22o_4.ext - technology: sky130A

.subckt sky130_fd_sc_hd__a22o_4 B1 B2 X A2 A1 VGND VPWR VNB VPB
X0 a_484_297.t2 B2.t0 a_96_21.t2 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 VGND.t1 B2.t1 a_566_47.t1 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 X.t5 a_96_21.t8 VGND.t6 VNB.t7 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 VPWR.t4 a_96_21.t9 X.t7 VPB.t7 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 X.t6 a_96_21.t10 VPWR.t3 VPB.t6 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 a_96_21.t7 B1.t0 a_484_297.t7 VPB.t11 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 VPWR.t2 a_96_21.t11 X.t1 VPB.t5 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 X.t4 a_96_21.t12 VGND.t5 VNB.t6 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 VGND.t4 a_96_21.t13 X.t3 VNB.t5 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 a_484_297.t0 B1.t1 a_96_21.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 a_484_297.t4 A2.t0 VPWR.t5 VPB.t8 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 VGND.t2 A2.t1 a_918_47.t2 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 a_96_21.t1 B2.t2 a_484_297.t1 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13 a_96_21.t4 B1.t2 a_566_47.t2 VNB.t8 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14 a_484_297.t5 A1.t0 VPWR.t6 VPB.t9 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 VPWR.t0 A1.t1 a_484_297.t3 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16 a_96_21.t6 A1.t2 a_918_47.t3 VNB.t10 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X17 VPWR.t7 A2.t2 a_484_297.t6 VPB.t10 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X18 a_566_47.t0 B2.t3 VGND.t0 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X19 a_918_47.t0 A1.t3 a_96_21.t3 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X20 a_566_47.t3 B1.t3 a_96_21.t5 VNB.t9 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X21 a_918_47.t1 A2.t3 VGND.t7 VNB.t11 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X22 X.t0 a_96_21.t14 VPWR.t1 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X23 VGND.t3 a_96_21.t15 X.t2 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
R0 B2.n1 B2.t2 241.534
R1 B2.n0 B2.t0 241.534
R2 B2.n1 B2.t3 169.234
R3 B2.n0 B2.t1 169.234
R4 B2.n2 B2.n0 162.479
R5 B2.n2 B2.n1 76
R6 B2 B2.n2 6.874
R7 a_96_21.n16 a_96_21.n0 346.333
R8 a_96_21.n17 a_96_21.n16 292.5
R9 a_96_21.n14 a_96_21.n12 213.809
R10 a_96_21.n9 a_96_21.t9 212.079
R11 a_96_21.n6 a_96_21.t10 212.079
R12 a_96_21.n3 a_96_21.t11 212.079
R13 a_96_21.n1 a_96_21.t14 212.079
R14 a_96_21.n9 a_96_21.t13 139.779
R15 a_96_21.n6 a_96_21.t8 139.779
R16 a_96_21.n3 a_96_21.t15 139.779
R17 a_96_21.n1 a_96_21.t12 139.779
R18 a_96_21.n5 a_96_21.n2 97.76
R19 a_96_21.n15 a_96_21.n14 96.493
R20 a_96_21.n14 a_96_21.n13 92.5
R21 a_96_21.n16 a_96_21.n15 77.591
R22 a_96_21.n8 a_96_21.n7 76
R23 a_96_21.n5 a_96_21.n4 76
R24 a_96_21.n11 a_96_21.n10 76
R25 a_96_21.n0 a_96_21.t2 26.595
R26 a_96_21.n0 a_96_21.t7 26.595
R27 a_96_21.t0 a_96_21.n17 26.595
R28 a_96_21.n17 a_96_21.t1 26.595
R29 a_96_21.n13 a_96_21.t5 24.923
R30 a_96_21.n13 a_96_21.t4 24.923
R31 a_96_21.n12 a_96_21.t3 24.923
R32 a_96_21.n12 a_96_21.t6 24.923
R33 a_96_21.n2 a_96_21.n1 21.909
R34 a_96_21.n11 a_96_21.n8 21.76
R35 a_96_21.n8 a_96_21.n5 21.76
R36 a_96_21.n10 a_96_21.n9 13.145
R37 a_96_21.n15 a_96_21.n11 11.2
R38 a_96_21.n4 a_96_21.n3 10.224
R39 a_96_21.n7 a_96_21.n6 1.46
R40 a_484_297.n1 a_484_297.t1 585.006
R41 a_484_297.n1 a_484_297.n0 292.5
R42 a_484_297.n3 a_484_297.t4 179.392
R43 a_484_297.n3 a_484_297.n2 155.085
R44 a_484_297.n5 a_484_297.n4 143.027
R45 a_484_297.n4 a_484_297.n1 58.68
R46 a_484_297.n4 a_484_297.n3 54.362
R47 a_484_297.n5 a_484_297.t6 35.46
R48 a_484_297.t2 a_484_297.n5 33.49
R49 a_484_297.n0 a_484_297.t7 26.595
R50 a_484_297.n0 a_484_297.t0 26.595
R51 a_484_297.n2 a_484_297.t3 26.595
R52 a_484_297.n2 a_484_297.t5 26.595
R53 VPB.t7 VPB.t1 556.386
R54 VPB.t2 VPB.t10 295.95
R55 VPB.t3 VPB.t8 248.598
R56 VPB.t9 VPB.t3 248.598
R57 VPB.t10 VPB.t9 248.598
R58 VPB.t11 VPB.t2 248.598
R59 VPB.t0 VPB.t11 248.598
R60 VPB.t1 VPB.t0 248.598
R61 VPB.t6 VPB.t7 248.598
R62 VPB.t5 VPB.t6 248.598
R63 VPB.t4 VPB.t5 248.598
R64 VPB VPB.t4 242.679
R65 a_566_47.n1 a_566_47.n0 233.872
R66 a_566_47.n0 a_566_47.t1 24.923
R67 a_566_47.n0 a_566_47.t3 24.923
R68 a_566_47.n1 a_566_47.t2 24.923
R69 a_566_47.t0 a_566_47.n1 24.923
R70 VGND.n25 VGND.t5 188.321
R71 VGND.n2 VGND.t2 125.619
R72 VGND.n1 VGND.n0 115.464
R73 VGND.n20 VGND.n19 115.464
R74 VGND.n10 VGND.n9 92.5
R75 VGND.n14 VGND.n13 92.5
R76 VGND.n0 VGND.t1 33.23
R77 VGND.n0 VGND.t7 31.384
R78 VGND.n9 VGND.t0 24.923
R79 VGND.n13 VGND.t4 24.923
R80 VGND.n19 VGND.t6 24.923
R81 VGND.n19 VGND.t3 24.923
R82 VGND.n26 VGND.n25 13.308
R83 VGND.n2 VGND.n1 11.666
R84 VGND.n4 VGND.n3 4.65
R85 VGND.n6 VGND.n5 4.65
R86 VGND.n8 VGND.n7 4.65
R87 VGND.n12 VGND.n11 4.65
R88 VGND.n16 VGND.n15 4.65
R89 VGND.n18 VGND.n17 4.65
R90 VGND.n22 VGND.n21 4.65
R91 VGND.n24 VGND.n23 4.65
R92 VGND.n21 VGND.n20 2.635
R93 VGND.n15 VGND.n14 0.9
R94 VGND.n11 VGND.n10 0.3
R95 VGND.n4 VGND.n2 0.137
R96 VGND.n6 VGND.n4 0.119
R97 VGND.n8 VGND.n6 0.119
R98 VGND.n12 VGND.n8 0.119
R99 VGND.n16 VGND.n12 0.119
R100 VGND.n18 VGND.n16 0.119
R101 VGND.n22 VGND.n18 0.119
R102 VGND.n24 VGND.n22 0.119
R103 VGND.n26 VGND.n24 0.119
R104 VGND VGND.n26 0.022
R105 VNB VNB.t6 6489.08
R106 VNB.t5 VNB.t0 4545.05
R107 VNB.t1 VNB.t11 2417.58
R108 VNB.t3 VNB.t2 2030.77
R109 VNB.t10 VNB.t3 2030.77
R110 VNB.t11 VNB.t10 2030.77
R111 VNB.t9 VNB.t1 2030.77
R112 VNB.t8 VNB.t9 2030.77
R113 VNB.t0 VNB.t8 2030.77
R114 VNB.t7 VNB.t5 2030.77
R115 VNB.t4 VNB.t7 2030.77
R116 VNB.t6 VNB.t4 2030.77
R117 X.n2 X.n0 155.695
R118 X.n2 X.n1 111.273
R119 X.n5 X.n3 88.89
R120 X.n5 X.n4 52.624
R121 X X.n2 39.416
R122 X X.n5 29.379
R123 X.n0 X.t7 26.595
R124 X.n0 X.t6 26.595
R125 X.n1 X.t1 26.595
R126 X.n1 X.t0 26.595
R127 X.n3 X.t3 24.923
R128 X.n3 X.t5 24.923
R129 X.n4 X.t2 24.923
R130 X.n4 X.t4 24.923
R131 VPWR.n14 VPWR.t4 552.677
R132 VPWR.n3 VPWR.n0 319.521
R133 VPWR.n2 VPWR.n1 314.004
R134 VPWR.n23 VPWR.t1 197.04
R135 VPWR.n19 VPWR.n18 170.445
R136 VPWR.n18 VPWR.t3 26.595
R137 VPWR.n18 VPWR.t2 26.595
R138 VPWR.n1 VPWR.t6 26.595
R139 VPWR.n1 VPWR.t7 26.595
R140 VPWR.n0 VPWR.t5 26.595
R141 VPWR.n0 VPWR.t0 26.595
R142 VPWR.n5 VPWR.n4 4.65
R143 VPWR.n7 VPWR.n6 4.65
R144 VPWR.n9 VPWR.n8 4.65
R145 VPWR.n11 VPWR.n10 4.65
R146 VPWR.n13 VPWR.n12 4.65
R147 VPWR.n15 VPWR.n14 4.65
R148 VPWR.n17 VPWR.n16 4.65
R149 VPWR.n20 VPWR.n19 4.65
R150 VPWR.n22 VPWR.n21 4.65
R151 VPWR.n24 VPWR.n23 4.65
R152 VPWR.n3 VPWR.n2 3.934
R153 VPWR.n5 VPWR.n3 0.317
R154 VPWR.n7 VPWR.n5 0.119
R155 VPWR.n9 VPWR.n7 0.119
R156 VPWR.n11 VPWR.n9 0.119
R157 VPWR.n13 VPWR.n11 0.119
R158 VPWR.n15 VPWR.n13 0.119
R159 VPWR.n17 VPWR.n15 0.119
R160 VPWR.n20 VPWR.n17 0.119
R161 VPWR.n22 VPWR.n20 0.119
R162 VPWR.n24 VPWR.n22 0.119
R163 VPWR VPWR.n24 0.022
R164 B1.n0 B1.t0 212.079
R165 B1.n1 B1.t1 212.079
R166 B1.n0 B1.t3 139.779
R167 B1.n1 B1.t2 139.779
R168 B1 B1.n2 77.268
R169 B1.n2 B1.n0 30.672
R170 B1.n2 B1.n1 30.672
R171 A2.n0 A2.t0 241.534
R172 A2.n1 A2.t2 241.534
R173 A2.n2 A2.n1 184.186
R174 A2.n0 A2.t1 169.234
R175 A2.n1 A2.t3 169.234
R176 A2.n2 A2.n0 76
R177 A2 A2.n2 22.4
R178 a_918_47.n1 a_918_47.n0 187.935
R179 a_918_47.n0 a_918_47.t3 24.923
R180 a_918_47.n0 a_918_47.t1 24.923
R181 a_918_47.t2 a_918_47.n1 24.923
R182 a_918_47.n1 a_918_47.t0 24.923
R183 A1.n0 A1.t1 212.079
R184 A1.n1 A1.t0 212.079
R185 A1.n0 A1.t3 139.779
R186 A1.n1 A1.t2 139.779
R187 A1 A1.n2 81.12
R188 A1.n2 A1.n0 30.672
R189 A1.n2 A1.n1 30.672
C0 VGND X 0.43fF
C1 VGND VPWR 0.14fF
C2 VPWR X 0.52fF
C3 A2 A1 0.31fF
C4 VPWR VPB 0.13fF
C5 B2 A2 0.14fF
C6 B2 B1 0.33fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__a22oi_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__a22oi_1 B1 A1 B2 A2 Y VPWR VGND VNB VPB
X0 Y.t2 B1.t0 a_109_47.t0 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 Y.t1 B1.t1 a_109_297.t2 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 VPWR.t1 A2.t0 a_109_297.t3 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 a_109_297.t0 A1.t0 VPWR.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 a_381_47.t1 A1.t1 Y.t3 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 a_109_297.t1 B2.t0 Y.t0 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 a_109_47.t1 B2.t1 VGND.t0 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 VGND.t1 A2.t1 a_381_47.t0 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
R0 B1.n0 B1.t1 239.503
R1 B1.n0 B1.t0 167.203
R2 B1 B1.n0 83.424
R3 a_109_47.t0 a_109_47.t1 42.461
R4 Y.n2 Y.t1 624.107
R5 Y.n1 Y.n0 192.977
R6 Y.n0 Y.t2 185.787
R7 Y.n0 Y.t3 157.115
R8 Y.n2 Y.t0 118.508
R9 Y Y.n3 78.577
R10 Y.n3 Y.n2 17.467
R11 Y Y.n1 6.044
R12 Y.n1 Y 4.945
R13 Y.n3 Y 3.49
R14 VNB VNB.t2 6053.91
R15 VNB.t1 VNB.t3 4738.46
R16 VNB.t2 VNB.t1 1837.36
R17 VNB.t3 VNB.t0 1740.66
R18 a_109_297.n1 a_109_297.n0 658.685
R19 a_109_297.n0 a_109_297.t2 26.595
R20 a_109_297.n0 a_109_297.t1 26.595
R21 a_109_297.n1 a_109_297.t3 26.595
R22 a_109_297.t0 a_109_297.n1 26.595
R23 VPB.t2 VPB.t0 556.386
R24 VPB.t0 VPB.t3 248.598
R25 VPB.t1 VPB.t2 248.598
R26 VPB VPB.t1 189.408
R27 A2.n0 A2.t0 241.534
R28 A2.n0 A2.t1 169.234
R29 A2 A2.n0 85.309
R30 VPWR.n0 VPWR.t0 577.692
R31 VPWR.n0 VPWR.t1 198.264
R32 VPWR VPWR.n0 0.479
R33 A1.n0 A1.t0 232.736
R34 A1.n0 A1.t1 160.436
R35 A1 A1.n0 79.352
R36 a_381_47.t0 a_381_47.t1 38.769
R37 B2.n0 B2.t0 241.534
R38 B2.n0 B2.t1 169.234
R39 B2 B2.n0 77.564
R40  B2 9.671
R41 VGND.n0 VGND.t1 150.218
R42 VGND.n0 VGND.t0 135.458
R43 VGND VGND.n0 0.052
C0 B2 B1 0.11fF
C1 B1 Y 0.18fF
C2 Y VPWR 0.32fF
C3 B2 Y 0.12fF
C4 VGND Y 0.36fF
C5 A1 A2 0.10fF
C6 A2 Y 0.20fF
C7 A1 Y 0.14fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__a22oi_2.ext - technology: sky130A

.subckt sky130_fd_sc_hd__a22oi_2 A1 A2 B1 B2 Y VPWR VGND VNB VPB
X0 a_109_297.t2 A2.t0 VPWR.t1 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_467_47.t1 A1.t0 Y.t1 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 VPWR.t0 A2.t1 a_109_297.t1 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 a_467_47.t3 A2.t2 VGND.t1 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 Y.t5 B1.t0 a_109_297.t6 VPB.t6 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 Y.t0 A1.t1 a_467_47.t0 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 a_109_297.t7 B1.t1 Y.t6 VPB.t7 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 VGND.t0 A2.t3 a_467_47.t2 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 Y.t4 B2.t0 a_109_297.t3 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 a_27_47.t3 B2.t1 VGND.t3 VNB.t6 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 a_27_47.t1 B1.t2 Y.t7 VNB.t7 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 a_109_297.t4 A1.t2 VPWR.t2 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 VPWR.t3 A1.t3 a_109_297.t5 VPB.t5 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13 Y.t2 B1.t3 a_27_47.t0 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14 a_109_297.t0 B2.t2 Y.t3 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 VGND.t2 B2.t3 a_27_47.t2 VNB.t5 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
R0 A2.n0 A2.t0 212.079
R1 A2.n1 A2.t1 212.079
R2 A2.n0 A2.t2 139.779
R3 A2.n1 A2.t3 139.779
R4 A2.n3 A2.n2 76
R5 A2.n2 A2.n0 48.2
R6 A2 A2.n3 16
R7 A2.n3 A2 13.44
R8 A2.n2 A2.n1 13.145
R9 VPWR.n3 VPWR.n0 185.045
R10 VPWR.n2 VPWR.n1 174.594
R11 VPWR.n14 VPWR 33.261
R12 VPWR.n1 VPWR.t2 26.595
R13 VPWR.n1 VPWR.t3 26.595
R14 VPWR.n0 VPWR.t1 26.595
R15 VPWR.n0 VPWR.t0 26.595
R16 VPWR.n3 VPWR.n2 12.212
R17 VPWR VPWR.n13 6.023
R18 VPWR.n7 VPWR.n6 4.65
R19 VPWR.n9 VPWR.n8 4.65
R20 VPWR.n11 VPWR.n10 4.65
R21 VPWR.n13 VPWR.n12 4.65
R22 VPWR.n5 VPWR.n4 4.65
R23 VPWR.n5 VPWR.n3 0.344
R24 VPWR.n7 VPWR.n5 0.119
R25 VPWR.n9 VPWR.n7 0.119
R26 VPWR.n11 VPWR.n9 0.119
R27 VPWR.n12 VPWR.n11 0.119
R28 VPWR.n14 VPWR.n12 0.119
R29 VPWR VPWR.n14 0.02
R30 a_109_297.n2 a_109_297.n1 209.372
R31 a_109_297.t2 a_109_297.n5 173.017
R32 a_109_297.n2 a_109_297.n0 151.6
R33 a_109_297.n3 a_109_297.t5 116.829
R34 a_109_297.n5 a_109_297.n4 108.022
R35 a_109_297.n3 a_109_297.n2 82.855
R36 a_109_297.n5 a_109_297.n3 59.439
R37 a_109_297.n0 a_109_297.t6 26.595
R38 a_109_297.n0 a_109_297.t7 26.595
R39 a_109_297.n1 a_109_297.t3 26.595
R40 a_109_297.n1 a_109_297.t0 26.595
R41 a_109_297.n4 a_109_297.t1 26.595
R42 a_109_297.n4 a_109_297.t4 26.595
R43 VPB.t6 VPB.t5 556.386
R44 VPB.t1 VPB.t2 248.598
R45 VPB.t4 VPB.t1 248.598
R46 VPB.t5 VPB.t4 248.598
R47 VPB.t7 VPB.t6 248.598
R48 VPB.t3 VPB.t7 248.598
R49 VPB.t0 VPB.t3 248.598
R50 VPB VPB.t0 189.408
R51 A1.n0 A1.t2 212.079
R52 A1.n1 A1.t3 212.079
R53 A1.n0 A1.t0 139.779
R54 A1.n1 A1.t1 139.779
R55 A1.n2 A1.n1 84.763
R56 A1.n1 A1.n0 61.345
R57 A1 A1.n2 20.48
R58 A1.n2 A1 8.96
R59 Y.n4 Y.t3 271.198
R60 Y.n5 Y.t5 173.58
R61 Y.n4 Y.n3 152.965
R62 Y.n2 Y.n1 146.711
R63 Y.n2 Y.n0 118.852
R64 Y.n6 Y.n4 38.4
R65 Y.n3 Y.t6 26.595
R66 Y.n3 Y.t4 26.595
R67 Y.n1 Y.t1 24.923
R68 Y.n1 Y.t0 24.923
R69 Y.n0 Y.t7 24.923
R70 Y.n0 Y.t2 24.923
R71 Y.n6 Y.n5 5.031
R72 Y.n7 Y.n6 2.825
R73 Y.n5 Y 2.088
R74 Y.n7 Y 1.765
R75 Y Y.n7 1.329
R76 Y Y.n2 0.22
R77 a_467_47.n0 a_467_47.t0 205.017
R78 a_467_47.n0 a_467_47.t3 190.352
R79 a_467_47.n1 a_467_47.n0 92.5
R80 a_467_47.n1 a_467_47.t2 24.923
R81 a_467_47.t1 a_467_47.n1 24.923
R82 VNB VNB.t5 6053.91
R83 VNB.t7 VNB.t0 4545.05
R84 VNB.t3 VNB.t4 2030.77
R85 VNB.t1 VNB.t3 2030.77
R86 VNB.t0 VNB.t1 2030.77
R87 VNB.t2 VNB.t7 2030.77
R88 VNB.t6 VNB.t2 2030.77
R89 VNB.t5 VNB.t6 2030.77
R90 VGND.n3 VGND.n2 112.801
R91 VGND.n1 VGND.n0 108.015
R92 VGND.n0 VGND.t3 24.923
R93 VGND.n0 VGND.t2 24.923
R94 VGND.n2 VGND.t1 24.923
R95 VGND.n2 VGND.t0 24.923
R96 VGND.n3 VGND.n1 3.418
R97 VGND.n1 VGND 3.296
R98 VGND VGND.n3 0.142
R99 B1.n0 B1.t0 212.079
R100 B1.n1 B1.t1 212.079
R101 B1.n0 B1.t2 139.779
R102 B1.n1 B1.t3 139.779
R103 B1.n3 B1.n2 76
R104 B1.n2 B1.n0 48.2
R105 B1 B1.n3 21.12
R106 B1.n2 B1.n1 13.145
R107 B1.n3 B1 8.32
R108 B2.n0 B2.t0 212.079
R109 B2.n1 B2.t2 212.079
R110 B2.n0 B2.t1 139.779
R111 B2.n1 B2.t3 139.779
R112 B2.n2 B2.n1 84.763
R113 B2.n1 B2.n0 61.345
R114 B2 B2.n2 16.64
R115 B2.n2 B2 12.8
R116 a_27_47.t1 a_27_47.n1 205.017
R117 a_27_47.n1 a_27_47.t2 192.536
R118 a_27_47.n1 a_27_47.n0 92.5
R119 a_27_47.n0 a_27_47.t0 24.923
R120 a_27_47.n0 a_27_47.t3 24.923
C0 B1 Y 0.22fF
C1 B2 Y 0.14fF
C2 Y A1 0.10fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__a22oi_4.ext - technology: sky130A

.subckt sky130_fd_sc_hd__a22oi_4 A2 B2 A1 B1 Y VGND VPWR VNB VPB
X0 a_27_47.t3 B1.t0 Y.t7 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 a_27_47.t2 B1.t1 Y.t6 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 a_27_297.t7 A2.t0 VPWR.t3 VPB.t7 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 Y.t3 B1.t2 a_27_297.t3 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 a_27_297.t10 B2.t0 Y.t11 VPB.t10 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 VPWR.t2 A2.t1 a_27_297.t6 VPB.t6 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 a_27_297.t5 A2.t2 VPWR.t1 VPB.t5 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 Y.t14 A1.t0 a_803_47.t7 VNB.t14 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 Y.t12 B2.t1 a_27_297.t11 VPB.t11 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 VPWR.t0 A2.t3 a_27_297.t4 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 Y.t15 A1.t1 a_803_47.t6 VNB.t15 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 VGND.t3 A2.t4 a_803_47.t3 VNB.t10 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 a_27_297.t13 B2.t2 Y.t13 VPB.t13 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13 a_27_47.t6 B2.t3 VGND.t7 VNB.t12 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14 a_27_47.t7 B2.t4 VGND.t6 VNB.t13 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X15 a_803_47.t5 A1.t2 Y.t10 VNB.t9 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X16 a_27_297.t2 B1.t3 Y.t2 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17 a_803_47.t4 A1.t3 Y.t8 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X18 a_803_47.t2 A2.t5 VGND.t2 VNB.t11 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X19 a_803_47.t1 A2.t6 VGND.t1 VNB.t7 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X20 VGND.t5 B2.t5 a_27_47.t4 VNB.t5 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X21 Y.t5 B1.t4 a_27_47.t1 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X22 Y.t1 B1.t5 a_27_297.t1 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X23 a_27_297.t12 A1.t4 VPWR.t5 VPB.t12 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X24 Y.t4 B1.t6 a_27_47.t0 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X25 a_27_297.t0 B1.t7 Y.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X26 VPWR.t4 A1.t5 a_27_297.t8 VPB.t8 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X27 a_27_297.t14 A1.t6 VPWR.t6 VPB.t14 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X28 VGND.t0 A2.t7 a_803_47.t0 VNB.t8 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X29 Y.t9 B2.t6 a_27_297.t9 VPB.t9 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X30 VPWR.t7 A1.t7 a_27_297.t15 VPB.t15 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X31 VGND.t4 B2.t7 a_27_47.t5 VNB.t6 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
R0 B1.n0 B1.t3 212.079
R1 B1.n1 B1.t5 212.079
R2 B1.n4 B1.t7 212.079
R3 B1.n3 B1.t2 212.079
R4 B1.n0 B1.t1 139.779
R5 B1.n1 B1.t6 139.779
R6 B1.n4 B1.t0 139.779
R7 B1.n3 B1.t4 139.779
R8 B1 B1.n5 82.08
R9 B1.n4 B1.n3 61.345
R10 B1 B1.n2 53.159
R11 B1.n2 B1.n1 36.77
R12 B1.n5 B1.n4 35.784
R13 B1.n2 B1.n0 18.368
R14 Y.n9 Y.n7 205.672
R15 Y.n14 Y.n13 156.435
R16 Y.n12 Y.n11 154.829
R17 Y.n9 Y.n8 150.416
R18 Y.n2 Y.n0 137.3
R19 Y.n6 Y.n5 94.292
R20 Y.n4 Y.n3 92.5
R21 Y.n2 Y.n1 92.5
R22 Y.n4 Y.n2 72.533
R23 Y.n12 Y.n10 47.999
R24 Y.n6 Y.n4 40.266
R25 Y.n10 Y.n6 34.816
R26 Y.n13 Y.t13 26.595
R27 Y.n13 Y.t9 26.595
R28 Y.n8 Y.t0 26.595
R29 Y.n8 Y.t3 26.595
R30 Y.n7 Y.t2 26.595
R31 Y.n7 Y.t1 26.595
R32 Y.n11 Y.t11 26.595
R33 Y.n11 Y.t12 26.595
R34 Y.n5 Y.t7 24.923
R35 Y.n5 Y.t5 24.923
R36 Y.n0 Y.t10 24.923
R37 Y.n0 Y.t14 24.923
R38 Y.n1 Y.t8 24.923
R39 Y.n1 Y.t15 24.923
R40 Y.n3 Y.t6 24.923
R41 Y.n3 Y.t4 24.923
R42  Y.n12 23.111
R43  Y.n14 18.844
R44 Y.n14 Y 5.485
R45 Y.n10 Y.n9 2.844
R46 a_27_47.n4 a_27_47.t2 219.833
R47 a_27_47.n1 a_27_47.t5 128.218
R48 a_27_47.n5 a_27_47.n4 92.5
R49 a_27_47.n4 a_27_47.n3 53.163
R50 a_27_47.n1 a_27_47.n0 52.624
R51 a_27_47.n3 a_27_47.n1 48.574
R52 a_27_47.n3 a_27_47.n2 42.273
R53 a_27_47.n2 a_27_47.t1 24.923
R54 a_27_47.n2 a_27_47.t7 24.923
R55 a_27_47.n0 a_27_47.t4 24.923
R56 a_27_47.n0 a_27_47.t6 24.923
R57 a_27_47.n5 a_27_47.t0 24.923
R58 a_27_47.t3 a_27_47.n5 24.923
R59 VNB VNB.t6 6053.91
R60 VNB.t2 VNB.t15 4545.05
R61 VNB.t8 VNB.t7 2030.77
R62 VNB.t11 VNB.t8 2030.77
R63 VNB.t10 VNB.t11 2030.77
R64 VNB.t9 VNB.t10 2030.77
R65 VNB.t14 VNB.t9 2030.77
R66 VNB.t4 VNB.t14 2030.77
R67 VNB.t15 VNB.t4 2030.77
R68 VNB.t0 VNB.t2 2030.77
R69 VNB.t3 VNB.t0 2030.77
R70 VNB.t1 VNB.t3 2030.77
R71 VNB.t13 VNB.t1 2030.77
R72 VNB.t5 VNB.t13 2030.77
R73 VNB.t12 VNB.t5 2030.77
R74 VNB.t6 VNB.t12 2030.77
R75 A2.n0 A2.t0 212.079
R76 A2.n2 A2.t1 212.079
R77 A2.n7 A2.t2 212.079
R78 A2.n5 A2.t3 212.079
R79 A2.n0 A2.t6 139.779
R80 A2.n2 A2.t7 139.779
R81 A2.n7 A2.t5 139.779
R82 A2.n5 A2.t4 139.779
R83 A2.n9 A2.n6 96.723
R84 A2.n4 A2.n1 96.723
R85 A2.n4 A2.n3 76
R86 A2.n9 A2.n8 76
R87 A2.n1 A2.n0 21.909
R88 A2.n6 A2.n5 13.145
R89 A2 A2.n4 11.58
R90 A2.n3 A2.n2 10.224
R91 A2 A2.n9 9.142
R92 A2.n8 A2.n7 1.46
R93 VPWR.n5 VPWR.n4 175.594
R94 VPWR.n1 VPWR.n0 171.981
R95 VPWR.n3 VPWR.n2 171.981
R96 VPWR.n9 VPWR.n8 171.981
R97 VPWR.n4 VPWR.t3 26.595
R98 VPWR.n4 VPWR.t2 26.595
R99 VPWR.n2 VPWR.t1 26.595
R100 VPWR.n2 VPWR.t0 26.595
R101 VPWR.n8 VPWR.t5 26.595
R102 VPWR.n8 VPWR.t4 26.595
R103 VPWR.n0 VPWR.t6 26.595
R104 VPWR.n0 VPWR.t7 26.595
R105 VPWR.n13 VPWR.n1 9.034
R106 VPWR.n7 VPWR.n6 4.65
R107 VPWR.n10 VPWR.n9 4.65
R108 VPWR.n12 VPWR.n11 4.65
R109 VPWR.n5 VPWR.n3 3.855
R110 VPWR VPWR.n13 1.082
R111 VPWR.n7 VPWR.n5 0.232
R112 VPWR.n13 VPWR.n12 0.134
R113 VPWR.n10 VPWR.n7 0.119
R114 VPWR.n12 VPWR.n10 0.119
R115 a_27_297.n13 a_27_297.n3 193.753
R116 a_27_297.n5 a_27_297.t7 181.779
R117 a_27_297.n1 a_27_297.t9 174.73
R118 a_27_297.n14 a_27_297.n2 174.616
R119 a_27_297.n16 a_27_297.n15 154.573
R120 a_27_297.n1 a_27_297.n0 154.573
R121 a_27_297.n18 a_27_297.n17 154.572
R122 a_27_297.n12 a_27_297.n11 144.851
R123 a_27_297.n5 a_27_297.n4 110.76
R124 a_27_297.n7 a_27_297.n6 110.76
R125 a_27_297.n9 a_27_297.n8 110.76
R126 a_27_297.n10 a_27_297.n9 45.752
R127 a_27_297.n16 a_27_297.n14 45.752
R128 a_27_297.n7 a_27_297.n5 44.423
R129 a_27_297.n9 a_27_297.n7 44.423
R130 a_27_297.n17 a_27_297.n1 44.423
R131 a_27_297.n17 a_27_297.n16 44.423
R132 a_27_297.n3 a_27_297.t15 26.595
R133 a_27_297.n11 a_27_297.t2 26.595
R134 a_27_297.n4 a_27_297.t6 26.595
R135 a_27_297.n4 a_27_297.t5 26.595
R136 a_27_297.n6 a_27_297.t4 26.595
R137 a_27_297.n6 a_27_297.t12 26.595
R138 a_27_297.n8 a_27_297.t8 26.595
R139 a_27_297.n8 a_27_297.t14 26.595
R140 a_27_297.n15 a_27_297.t1 26.595
R141 a_27_297.n15 a_27_297.t0 26.595
R142 a_27_297.n0 a_27_297.t11 26.595
R143 a_27_297.n0 a_27_297.t13 26.595
R144 a_27_297.t3 a_27_297.n18 26.595
R145 a_27_297.n18 a_27_297.t10 26.595
R146 a_27_297.n13 a_27_297.n12 4.671
R147 a_27_297.n14 a_27_297.n13 3.744
R148 a_27_297.n12 a_27_297.n10 2.799
R149 VPB.t2 VPB.t15 556.386
R150 VPB.t6 VPB.t7 248.598
R151 VPB.t5 VPB.t6 248.598
R152 VPB.t4 VPB.t5 248.598
R153 VPB.t12 VPB.t4 248.598
R154 VPB.t8 VPB.t12 248.598
R155 VPB.t14 VPB.t8 248.598
R156 VPB.t15 VPB.t14 248.598
R157 VPB.t1 VPB.t2 248.598
R158 VPB.t0 VPB.t1 248.598
R159 VPB.t3 VPB.t0 248.598
R160 VPB.t10 VPB.t3 248.598
R161 VPB.t11 VPB.t10 248.598
R162 VPB.t13 VPB.t11 248.598
R163 VPB.t9 VPB.t13 248.598
R164 VPB VPB.t9 189.408
R165 B2.n0 B2.t0 212.079
R166 B2.n2 B2.t1 212.079
R167 B2.n7 B2.t2 212.079
R168 B2.n5 B2.t6 212.079
R169 B2.n0 B2.t4 139.779
R170 B2.n2 B2.t5 139.779
R171 B2.n7 B2.t3 139.779
R172 B2.n5 B2.t7 139.779
R173 B2.n9 B2.n6 97.76
R174 B2.n4 B2.n1 97.76
R175 B2.n4 B2.n3 76
R176 B2.n9 B2.n8 76
R177 B2.n6 B2.n5 21.909
R178 B2 B2.n4 14.72
R179 B2.n1 B2.n0 13.145
R180 B2.n8 B2.n7 10.224
R181 B2 B2.n9 7.04
R182 B2.n3 B2.n2 1.46
R183 A1.n0 A1.t4 212.079
R184 A1.n2 A1.t5 212.079
R185 A1.n5 A1.t6 212.079
R186 A1.n8 A1.t7 212.079
R187 A1.n0 A1.t2 139.779
R188 A1.n2 A1.t0 139.779
R189 A1.n5 A1.t3 139.779
R190 A1.n8 A1.t1 139.779
R191 A1.n4 A1.n1 96.723
R192 A1 A1.n9 96.114
R193 A1.n4 A1.n3 76
R194 A1.n7 A1.n6 76
R195 A1.n1 A1.n0 21.909
R196 A1.n7 A1.n4 20.723
R197 A1.n9 A1.n8 13.145
R198 A1.n3 A1.n2 10.224
R199 A1.n6 A1.n5 1.46
R200 A1 A1.n7 0.609
R201 a_803_47.t6 a_803_47.n5 219.833
R202 a_803_47.n1 a_803_47.t1 128.218
R203 a_803_47.n5 a_803_47.n4 92.5
R204 a_803_47.n5 a_803_47.n3 53.163
R205 a_803_47.n1 a_803_47.n0 52.624
R206 a_803_47.n3 a_803_47.n1 48.574
R207 a_803_47.n3 a_803_47.n2 42.273
R208 a_803_47.n4 a_803_47.t7 24.923
R209 a_803_47.n4 a_803_47.t4 24.923
R210 a_803_47.n2 a_803_47.t3 24.923
R211 a_803_47.n2 a_803_47.t5 24.923
R212 a_803_47.n0 a_803_47.t0 24.923
R213 a_803_47.n0 a_803_47.t2 24.923
R214 VGND.n1 VGND.n0 121.164
R215 VGND.n3 VGND.n2 115.464
R216 VGND.n25 VGND.n24 115.464
R217 VGND.n31 VGND.n30 115.464
R218 VGND.n0 VGND.t1 24.923
R219 VGND.n0 VGND.t0 24.923
R220 VGND.n2 VGND.t2 24.923
R221 VGND.n2 VGND.t3 24.923
R222 VGND.n24 VGND.t6 24.923
R223 VGND.n24 VGND.t5 24.923
R224 VGND.n30 VGND.t7 24.923
R225 VGND.n30 VGND.t4 24.923
R226 VGND.n26 VGND.n25 6.776
R227 VGND.n5 VGND.n4 4.65
R228 VGND.n7 VGND.n6 4.65
R229 VGND.n9 VGND.n8 4.65
R230 VGND.n11 VGND.n10 4.65
R231 VGND.n13 VGND.n12 4.65
R232 VGND.n15 VGND.n14 4.65
R233 VGND.n17 VGND.n16 4.65
R234 VGND.n19 VGND.n18 4.65
R235 VGND.n21 VGND.n20 4.65
R236 VGND.n23 VGND.n22 4.65
R237 VGND.n27 VGND.n26 4.65
R238 VGND.n29 VGND.n28 4.65
R239 VGND.n33 VGND.n32 4.65
R240 VGND.n4 VGND.n3 2.258
R241 VGND.n5 VGND.n1 0.978
R242 VGND.n32 VGND.n31 0.752
R243 VGND.n7 VGND.n5 0.119
R244 VGND.n9 VGND.n7 0.119
R245 VGND.n11 VGND.n9 0.119
R246 VGND.n13 VGND.n11 0.119
R247 VGND.n15 VGND.n13 0.119
R248 VGND.n17 VGND.n15 0.119
R249 VGND.n19 VGND.n17 0.119
R250 VGND.n21 VGND.n19 0.119
R251 VGND.n23 VGND.n21 0.119
R252 VGND.n27 VGND.n23 0.119
R253 VGND.n29 VGND.n27 0.119
R254 VGND.n33 VGND.n29 0.119
R255 VGND.n34 VGND.n33 0.119
R256 VGND VGND.n34 0.02
C0 VPWR VGND 0.16fF
C1 VPB VPWR 0.15fF
C2 B2 Y 0.25fF
C3 A1 Y 0.21fF
C4 B1 Y 0.43fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__a31o_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__a31o_1 A2 B1 A1 A3 X VGND VPWR VNB VPB
X0 VPWR.t3 a_80_21.t3 X.t1 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_209_297.t3 A3.t0 VPWR.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 a_303_47.t0 A2.t0 a_209_47.t0 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 a_209_47.t1 A3.t1 VGND.t2 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 VGND.t1 a_80_21.t4 X.t0 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 VGND.t0 B1.t0 a_80_21.t0 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 a_80_21.t2 A1.t0 a_303_47.t1 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 VPWR.t2 A2.t1 a_209_297.t2 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 a_80_21.t1 B1.t1 a_209_297.t1 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 a_209_297.t0 A1.t1 VPWR.t1 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
R0 a_80_21.t1 a_80_21.n2 321.583
R1 a_80_21.n0 a_80_21.t3 240.999
R2 a_80_21.n2 a_80_21.n0 193.117
R3 a_80_21.n0 a_80_21.t4 168.699
R4 a_80_21.n2 a_80_21.n1 49.328
R5 a_80_21.n1 a_80_21.t0 34.153
R6 a_80_21.n1 a_80_21.t2 26.769
R7 X.n2 X.n1 292.5
R8 X.n3 X.n2 147.104
R9 X.n0 X.t0 82.289
R10 X.n1 X.n0 63.654
R11 X.n2 X.t1 27.58
R12 X.n3 X 10.71
R13 X.n0 X 5.727
R14 X.n1 X 4.848
R15 X X.n3 2.439
R16 VPWR.n2 VPWR.n0 314.275
R17 VPWR.n2 VPWR.n1 129.562
R18 VPWR.n1 VPWR.t0 34.475
R19 VPWR.n1 VPWR.t3 33.49
R20 VPWR.n0 VPWR.t1 32.505
R21 VPWR.n0 VPWR.t2 32.505
R22 VPWR VPWR.n2 0.208
R23 VPB.t4 VPB.t0 292.99
R24 VPB.t1 VPB.t2 284.112
R25 VPB.t3 VPB.t1 284.112
R26 VPB.t0 VPB.t3 278.193
R27 VPB VPB.t4 192.367
R28 A3.n0 A3.t0 241.534
R29 A3.n0 A3.t1 169.234
R30 A3.n1 A3.n0 76
R31 A3.n1 A3 14.068
R32 A3 A3.n1 2.308
R33 a_209_297.n1 a_209_297.n0 360.435
R34 a_209_297.n0 a_209_297.t2 32.505
R35 a_209_297.n1 a_209_297.t1 32.505
R36 a_209_297.t0 a_209_297.n1 32.505
R37 a_209_297.n0 a_209_297.t3 30.535
R38 A2.n0 A2.t1 241.534
R39 A2.n0 A2.t0 169.234
R40 A2.n1 A2.n0 76
R41 A2.n1 A2 12.8
R42 A2 A2.n1 2.47
R43 a_209_47.t0 a_209_47.t1 59.076
R44 a_303_47.t0 a_303_47.t1 60.923
R45 VNB VNB.t2 6078.09
R46 VNB.t2 VNB.t3 2393.41
R47 VNB.t4 VNB.t0 2320.88
R48 VNB.t1 VNB.t4 2320.88
R49 VNB.t3 VNB.t1 2272.53
R50 VGND.n1 VGND.t0 142.283
R51 VGND.n1 VGND.n0 111.392
R52 VGND.n0 VGND.t1 38.769
R53 VGND.n0 VGND.t2 24.923
R54 VGND VGND.n1 0.149
R55 B1.n0 B1.t1 241.534
R56 B1.n0 B1.t0 169.234
R57 B1.n1 B1.n0 76
R58 B1.n1 B1 14.889
R59 B1 B1.n1 2.873
R60 A1.n0 A1.t1 241.534
R61 A1.n0 A1.t0 169.234
R62 A1.n1 A1.n0 76
R63 A1.n1 A1 13.766
R64 A1 A1.n1 2.656
C0 X VPWR 0.20fF
C1 A3 A2 0.13fF
C2 A2 A1 0.15fF
C3 A1 B1 0.14fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__a31o_2.ext - technology: sky130A

.subckt sky130_fd_sc_hd__a31o_2 X B1 A3 A1 A2 VGND VPWR VNB VPB
X0 VPWR.t4 A2.t0 a_277_297.t2 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_277_297.t0 A1.t0 VPWR.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 a_79_21.t2 B1.t0 a_277_297.t3 VPB.t5 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 a_277_297.t1 A3.t0 VPWR.t3 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 VPWR.t1 a_79_21.t3 X.t1 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 VGND.t2 a_79_21.t4 X.t3 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 a_361_47.t0 A2.t1 a_277_47.t1 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 a_277_47.t0 A3.t1 VGND.t0 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 VGND.t3 B1.t1 a_79_21.t1 VNB.t5 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 a_79_21.t0 A1.t1 a_361_47.t1 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 X.t0 a_79_21.t5 VPWR.t2 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 X.t2 a_79_21.t6 VGND.t1 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
R0 A2.n0 A2.t0 241.534
R1 A2.n0 A2.t1 169.234
R2 A2 A2.n0 123.647
R3 a_277_297.n1 a_277_297.n0 355.918
R4 a_277_297.t0 a_277_297.n1 38.415
R5 a_277_297.n0 a_277_297.t2 26.595
R6 a_277_297.n0 a_277_297.t1 26.595
R7 a_277_297.n1 a_277_297.t3 26.595
R8 VPWR.n6 VPWR.t2 580.936
R9 VPWR.n3 VPWR.n0 313.809
R10 VPWR.n2 VPWR.n1 169.933
R11 VPWR.n0 VPWR.t4 34.475
R12 VPWR.n0 VPWR.t0 30.535
R13 VPWR.n1 VPWR.t3 26.595
R14 VPWR.n1 VPWR.t1 26.595
R15 VPWR.n5 VPWR.n4 4.65
R16 VPWR.n7 VPWR.n6 4.65
R17 VPWR.n3 VPWR.n2 4.011
R18 VPWR.n5 VPWR.n3 0.225
R19 VPWR.n7 VPWR.n5 0.119
R20 VPWR VPWR.n7 0.02
R21 VPB.t0 VPB.t5 284.112
R22 VPB.t4 VPB.t0 284.112
R23 VPB.t3 VPB.t4 248.598
R24 VPB.t1 VPB.t3 248.598
R25 VPB.t2 VPB.t1 248.598
R26 VPB VPB.t2 189.408
R27 A1.n0 A1.t0 241.534
R28 A1.n0 A1.t1 169.234
R29 A1 A1.n0 126.929
R30 B1.n0 B1.t0 227.985
R31 B1.n0 B1.t1 155.685
R32 B1 B1.n0 79.61
R33 a_79_21.n4 a_79_21.n3 247.201
R34 a_79_21.t2 a_79_21.n4 238.609
R35 a_79_21.n1 a_79_21.t3 212.079
R36 a_79_21.n2 a_79_21.t5 212.079
R37 a_79_21.n4 a_79_21.n0 171.137
R38 a_79_21.n1 a_79_21.t4 139.779
R39 a_79_21.n2 a_79_21.t6 139.779
R40 a_79_21.n0 a_79_21.t0 47.076
R41 a_79_21.n3 a_79_21.n2 36.515
R42 a_79_21.n0 a_79_21.t1 24.923
R43 a_79_21.n3 a_79_21.n1 24.83
R44 A3.n0 A3.t0 241.534
R45 A3.n0 A3.t1 169.234
R46 A3.n1 A3.n0 81.624
R47 A3.n1 A3 14.36
R48 A3 A3.n1 3.684
R49 X X.n1 346.71
R50 X.n2 X.n0 139.934
R51 X.n1 X.t1 26.595
R52 X.n1 X.t0 26.595
R53 X.n0 X.t3 24.923
R54 X.n0 X.t2 24.923
R55 X.n2 X 15.309
R56 X X.n2 1.756
R57 VGND.n5 VGND.t1 194.65
R58 VGND.n2 VGND.t3 190.492
R59 VGND.n1 VGND.n0 107.239
R60 VGND.n0 VGND.t0 24.923
R61 VGND.n0 VGND.t2 24.923
R62 VGND.n6 VGND.n5 4.65
R63 VGND.n4 VGND.n3 4.65
R64 VGND.n2 VGND.n1 3.983
R65 VGND.n4 VGND.n2 0.139
R66 VGND.n6 VGND.n4 0.119
R67 VGND VGND.n6 0.02
R68 VNB VNB.t1 6053.91
R69 VNB.t4 VNB.t5 2610.99
R70 VNB.t3 VNB.t4 2320.88
R71 VNB.t0 VNB.t3 2030.77
R72 VNB.t2 VNB.t0 2030.77
R73 VNB.t1 VNB.t2 2030.77
R74 a_277_47.t0 a_277_47.t1 49.846
R75 a_361_47.t0 a_361_47.t1 60.923
C0 VPWR X 0.23fF
C1 A2 A1 0.15fF
C2 VGND X 0.15fF
C3 A3 A2 0.11fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__a31o_4.ext - technology: sky130A

.subckt sky130_fd_sc_hd__a31o_4 B1 A2 A3 A1 X VGND VPWR VNB VPB
X0 VPWR.t5 a_277_47.t6 X.t3 VPB.t7 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 X.t2 a_277_47.t7 VPWR.t4 VPB.t6 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 X.t1 a_277_47.t8 VPWR.t3 VPB.t5 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 VPWR.t8 A2.t0 a_27_297.t7 VPB.t10 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 a_27_297.t2 A3.t0 VPWR.t0 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 a_277_47.t0 B1.t0 a_27_297.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 a_27_297.t4 A1.t0 VPWR.t6 VPB.t8 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 VGND.t5 a_277_47.t9 X.t7 VNB.t5 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 VPWR.t7 A1.t1 a_27_297.t5 VPB.t9 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 VGND.t4 a_277_47.t10 X.t6 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 a_27_297.t6 A2.t1 VPWR.t9 VPB.t11 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 a_193_47.t0 A2.t2 a_109_47.t1 VNB.t9 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 a_361_47.t1 A1.t2 a_277_47.t4 VNB.t11 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 X.t5 a_277_47.t11 VGND.t3 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14 VGND.t0 A3.t1 a_445_47.t0 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X15 X.t4 a_277_47.t12 VGND.t2 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X16 a_277_47.t3 A1.t3 a_193_47.t1 VNB.t10 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X17 a_445_47.t1 A2.t3 a_361_47.t0 VNB.t8 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X18 VGND.t7 B1.t1 a_277_47.t1 VNB.t7 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X19 a_27_297.t1 B1.t2 a_277_47.t2 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X20 VPWR.t1 A3.t2 a_27_297.t3 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X21 VPWR.t2 a_277_47.t13 X.t0 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X22 a_109_47.t0 A3.t3 VGND.t1 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X23 a_277_47.t5 B1.t3 VGND.t6 VNB.t6 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
R0 a_277_47.n13 a_277_47.n11 225.769
R1 a_277_47.n1 a_277_47.t13 212.079
R2 a_277_47.n0 a_277_47.t7 212.079
R3 a_277_47.n5 a_277_47.t6 212.079
R4 a_277_47.n8 a_277_47.t8 212.079
R5 a_277_47.n15 a_277_47.n14 153.52
R6 a_277_47.n1 a_277_47.t9 139.779
R7 a_277_47.n0 a_277_47.t11 139.779
R8 a_277_47.n5 a_277_47.t10 139.779
R9 a_277_47.n8 a_277_47.t12 139.779
R10 a_277_47.n14 a_277_47.n10 78.886
R11 a_277_47.n10 a_277_47.n9 76
R12 a_277_47.n4 a_277_47.n3 76
R13 a_277_47.n7 a_277_47.n6 76
R14 a_277_47.n13 a_277_47.n12 55.724
R15 a_277_47.n4 a_277_47.n2 50.937
R16 a_277_47.n14 a_277_47.n13 48.432
R17 a_277_47.n2 a_277_47.n0 40.579
R18 a_277_47.n15 a_277_47.t2 26.595
R19 a_277_47.t0 a_277_47.n15 26.595
R20 a_277_47.n12 a_277_47.t1 24.923
R21 a_277_47.n12 a_277_47.t5 24.923
R22 a_277_47.n11 a_277_47.t4 24.923
R23 a_277_47.n11 a_277_47.t3 24.923
R24 a_277_47.n2 a_277_47.n1 15.961
R25 a_277_47.n7 a_277_47.n4 13.187
R26 a_277_47.n10 a_277_47.n7 13.187
R27 a_277_47.n6 a_277_47.n5 8.763
R28 a_277_47.n9 a_277_47.n8 2.921
R29 X.n2 X.n1 215.715
R30 X.n5 X.n4 155.747
R31 X.n2 X.n0 152.468
R32 X.n5 X.n3 92.5
R33 X X.n2 45.552
R34 X X.n5 45.552
R35 X.n1 X.t3 26.595
R36 X.n1 X.t1 26.595
R37 X.n0 X.t0 26.595
R38 X.n0 X.t2 26.595
R39 X.n3 X.t7 24.923
R40 X.n3 X.t5 24.923
R41 X.n4 X.t6 24.923
R42 X.n4 X.t4 24.923
R43 X X.n6 21.082
R44 X.n6 X 6.4
R45 X.n6 X 4.517
R46 VPWR.n5 VPWR.t3 482.761
R47 VPWR.n2 VPWR.t2 404.781
R48 VPWR.n1 VPWR.n0 312.281
R49 VPWR.n14 VPWR.n13 312.281
R50 VPWR.n20 VPWR.n19 312.281
R51 VPWR.n25 VPWR.n24 312.281
R52 VPWR.n13 VPWR.t0 38.415
R53 VPWR.n0 VPWR.t4 26.595
R54 VPWR.n0 VPWR.t5 26.595
R55 VPWR.n13 VPWR.t8 26.595
R56 VPWR.n19 VPWR.t6 26.595
R57 VPWR.n19 VPWR.t7 26.595
R58 VPWR.n24 VPWR.t9 26.595
R59 VPWR.n24 VPWR.t1 26.595
R60 VPWR.n2 VPWR.n1 5.684
R61 VPWR.n4 VPWR.n3 4.65
R62 VPWR.n6 VPWR.n5 4.65
R63 VPWR.n8 VPWR.n7 4.65
R64 VPWR.n10 VPWR.n9 4.65
R65 VPWR.n12 VPWR.n11 4.65
R66 VPWR.n16 VPWR.n15 4.65
R67 VPWR.n18 VPWR.n17 4.65
R68 VPWR.n21 VPWR.n20 4.65
R69 VPWR.n23 VPWR.n22 4.65
R70 VPWR.n26 VPWR.n25 3.932
R71 VPWR.n4 VPWR.n2 0.465
R72 VPWR.n15 VPWR.n14 0.376
R73 VPWR.n26 VPWR.n23 0.137
R74 VPWR VPWR.n26 0.121
R75 VPWR.n6 VPWR.n4 0.119
R76 VPWR.n8 VPWR.n6 0.119
R77 VPWR.n10 VPWR.n8 0.119
R78 VPWR.n12 VPWR.n10 0.119
R79 VPWR.n16 VPWR.n12 0.119
R80 VPWR.n18 VPWR.n16 0.119
R81 VPWR.n21 VPWR.n18 0.119
R82 VPWR.n23 VPWR.n21 0.119
R83 VPB.t1 VPB.t5 556.386
R84 VPB.t2 VPB.t0 284.112
R85 VPB.t10 VPB.t2 284.112
R86 VPB.t6 VPB.t4 248.598
R87 VPB.t7 VPB.t6 248.598
R88 VPB.t5 VPB.t7 248.598
R89 VPB.t0 VPB.t1 248.598
R90 VPB.t8 VPB.t10 248.598
R91 VPB.t9 VPB.t8 248.598
R92 VPB.t11 VPB.t9 248.598
R93 VPB.t3 VPB.t11 248.598
R94 VPB VPB.t3 189.408
R95 A2.n1 A2.t1 241.534
R96 A2.n0 A2.t0 241.534
R97 A2.n2 A2.n1 174.543
R98 A2.n1 A2.t2 169.234
R99 A2.n0 A2.t3 169.234
R100 A2.n3 A2.n0 80.8
R101 A2.n3 A2.n2 17.643
R102 A2 A2.n3 5.44
R103 A2.n2 A2 3.805
R104 a_27_297.n1 a_27_297.t1 254.402
R105 a_27_297.n4 a_27_297.t3 242.31
R106 a_27_297.n5 a_27_297.n4 152.469
R107 a_27_297.n3 a_27_297.n2 152.468
R108 a_27_297.n1 a_27_297.n0 140.119
R109 a_27_297.n3 a_27_297.n1 84.546
R110 a_27_297.n4 a_27_297.n3 63.247
R111 a_27_297.n0 a_27_297.t2 38.415
R112 a_27_297.n2 a_27_297.t7 26.595
R113 a_27_297.n2 a_27_297.t4 26.595
R114 a_27_297.n0 a_27_297.t0 26.595
R115 a_27_297.n5 a_27_297.t5 26.595
R116 a_27_297.t6 a_27_297.n5 26.595
R117 A3 A3.n0 243.84
R118 A3.n0 A3.t0 241.534
R119 A3.n1 A3.t2 236.932
R120 A3.n0 A3.t1 169.234
R121 A3.n1 A3.t3 164.632
R122 A3.n2 A3.n1 76
R123 A3.n2 A3 9.728
R124 A3 A3.n2 1.877
R125 B1.n1 B1.t2 212.079
R126 B1.n0 B1.t0 212.079
R127 B1.n1 B1.t1 139.779
R128 B1.n0 B1.t3 139.779
R129 B1 B1.n1 120.09
R130 B1.n1 B1.n0 61.345
R131 A1.n0 A1.t0 221.719
R132 A1.n1 A1.t1 221.719
R133 A1.n0 A1.t2 149.419
R134 A1.n1 A1.t3 149.419
R135 A1 A1.n2 78.011
R136 A1.n2 A1.n0 37.488
R137 A1.n2 A1.n1 37.488
R138 VGND.n2 VGND.t5 185.711
R139 VGND.n29 VGND.t1 114.773
R140 VGND.n16 VGND.n15 108.892
R141 VGND.n1 VGND.n0 108.015
R142 VGND.n8 VGND.n7 92.5
R143 VGND.n10 VGND.n9 92.5
R144 VGND.n7 VGND.t2 39.692
R145 VGND.n9 VGND.t7 39.692
R146 VGND.n15 VGND.t0 32.307
R147 VGND.n15 VGND.t6 28.615
R148 VGND.n0 VGND.t3 24.923
R149 VGND.n0 VGND.t4 24.923
R150 VGND.n30 VGND.n29 6.908
R151 VGND.n2 VGND.n1 5.684
R152 VGND.n11 VGND.n8 5.316
R153 VGND.n4 VGND.n3 4.65
R154 VGND.n6 VGND.n5 4.65
R155 VGND.n12 VGND.n11 4.65
R156 VGND.n14 VGND.n13 4.65
R157 VGND.n18 VGND.n17 4.65
R158 VGND.n20 VGND.n19 4.65
R159 VGND.n22 VGND.n21 4.65
R160 VGND.n24 VGND.n23 4.65
R161 VGND.n26 VGND.n25 4.65
R162 VGND.n28 VGND.n27 4.65
R163 VGND.n11 VGND.n10 1.772
R164 VGND.n4 VGND.n2 0.465
R165 VGND.n17 VGND.n16 0.376
R166 VGND.n6 VGND.n4 0.119
R167 VGND.n12 VGND.n6 0.119
R168 VGND.n14 VGND.n12 0.119
R169 VGND.n18 VGND.n14 0.119
R170 VGND.n20 VGND.n18 0.119
R171 VGND.n22 VGND.n20 0.119
R172 VGND.n24 VGND.n22 0.119
R173 VGND.n26 VGND.n24 0.119
R174 VGND.n28 VGND.n26 0.119
R175 VGND.n30 VGND.n28 0.119
R176 VGND VGND.n30 0.02
R177 VNB VNB.t0 6053.91
R178 VNB.t7 VNB.t2 4545.05
R179 VNB.t1 VNB.t6 2320.88
R180 VNB.t8 VNB.t1 2320.88
R181 VNB.t3 VNB.t5 2030.77
R182 VNB.t4 VNB.t3 2030.77
R183 VNB.t2 VNB.t4 2030.77
R184 VNB.t6 VNB.t7 2030.77
R185 VNB.t11 VNB.t8 2030.77
R186 VNB.t10 VNB.t11 2030.77
R187 VNB.t9 VNB.t10 2030.77
R188 VNB.t0 VNB.t9 2030.77
R189 a_109_47.t0 a_109_47.t1 49.846
R190 a_193_47.t0 a_193_47.t1 49.846
R191 a_361_47.t0 a_361_47.t1 49.846
R192 a_445_47.t0 a_445_47.t1 60.923
C0 A3 A2 0.33fF
C1 VPWR VGND 0.15fF
C2 A2 A1 0.23fF
C3 VPB VPWR 0.13fF
C4 VPWR X 0.43fF
C5 X VGND 0.20fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__a31oi_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__a31oi_1 VGND VPWR Y B1 A2 A1 A3 VNB VPB
X0 Y.t1 A1.t0 a_181_47.t1 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 a_181_47.t0 A2.t0 a_109_47.t0 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 VGND.t0 B1.t0 Y.t0 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 VPWR.t0 A2.t1 a_109_297.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 Y.t2 B1.t1 a_109_297.t2 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 a_109_297.t1 A1.t1 VPWR.t1 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 a_109_297.t3 A3.t0 VPWR.t2 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 a_109_47.t1 A3.t1 VGND.t1 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
R0 A1.n0 A1.t1 241.534
R1 A1.n0 A1.t0 169.234
R2 A1 A1.n0 112.59
R3 a_181_47.t0 a_181_47.t1 67.384
R4 Y.n1 Y.n0 147.091
R5 Y.n3 Y.n2 130.604
R6 Y.n2 Y.t0 35.076
R7 Y.n0 Y.t2 28.565
R8 Y.n2 Y.t1 24.923
R9 Y Y.n1 10.551
R10 Y Y.n3 4.776
R11 Y.n1 Y 2.402
R12 VNB VNB.t3 6053.91
R13 VNB.t1 VNB.t2 2490.11
R14 VNB.t2 VNB.t0 2296.7
R15 VNB.t3 VNB.t1 1740.66
R16 A2.n0 A2.t1 241.534
R17 A2.n0 A2.t0 169.234
R18 A2 A2.n0 77.582
R19 a_109_47.t0 a_109_47.t1 38.769
R20 B1.n0 B1.t1 229.752
R21 B1.n0 B1.t0 157.452
R22 B1 B1.n0 78.909
R23 VGND.n0 VGND.t0 187.753
R24 VGND.n0 VGND.t1 107.117
R25 VGND VGND.n0 0.043
R26 a_109_297.n1 a_109_297.n0 680.992
R27 a_109_297.n0 a_109_297.t2 37.43
R28 a_109_297.n0 a_109_297.t1 26.595
R29 a_109_297.t0 a_109_297.n1 26.595
R30 a_109_297.n1 a_109_297.t3 26.595
R31 VPWR.n1 VPWR.n0 310.721
R32 VPWR.n1 VPWR.t2 149.637
R33 VPWR.n0 VPWR.t1 33.49
R34 VPWR.n0 VPWR.t0 26.595
R35 VPWR VPWR.n1 0.153
R36 VPB.t1 VPB.t2 281.152
R37 VPB.t0 VPB.t1 269.314
R38 VPB.t3 VPB.t0 248.598
R39 VPB VPB.t3 189.408
R40 A3.n0 A3.t0 230.154
R41 A3.n0 A3.t1 157.854
R42 A3 A3.n0 79.684
C0 B1 Y 0.11fF
C1 VGND Y 0.11fF
C2 VGND A2 0.11fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__a31oi_2.ext - technology: sky130A

.subckt sky130_fd_sc_hd__a31oi_2 A3 B1 Y A1 A2 VPWR VGND VNB VPB
X0 VGND.t3 B1.t0 Y.t4 VNB.t6 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 VPWR.t5 A1.t0 a_27_297.t7 VPB.t7 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 a_27_297.t4 A2.t0 VPWR.t2 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 a_27_297.t3 B1.t1 Y.t2 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 a_277_47.t1 A1.t1 Y.t0 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 VPWR.t0 A2.t1 a_27_297.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 a_27_297.t5 A3.t0 VPWR.t3 VPB.t5 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 a_27_47.t1 A3.t1 VGND.t0 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 a_27_47.t3 A2.t2 a_277_47.t3 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 a_27_297.t6 A1.t2 VPWR.t4 VPB.t6 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 Y.t1 B1.t2 a_27_297.t2 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 a_277_47.t2 A2.t3 a_27_47.t2 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 Y.t3 B1.t3 VGND.t2 VNB.t5 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 Y.t5 A1.t3 a_277_47.t0 VNB.t7 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14 VPWR.t1 A3.t2 a_27_297.t1 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 VGND.t1 A3.t3 a_27_47.t0 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
R0 B1.n4 B1.t1 212.079
R1 B1.n0 B1.t2 212.079
R2 B1.n4 B1.t3 139.779
R3 B1.n0 B1.t0 139.779
R4 B1.n5 B1.n4 104.481
R5 B1.n2 B1.n1 76
R6 B1.n1 B1.n0 51.851
R7 B1.n3 B1.n2 17.92
R8 B1.n3 B1 15.36
R9 B1.n2 B1 10.56
R10 B1 B1.n5 3.128
R11 B1.n5 B1.n3 0.853
R12 Y.n2 Y.t0 235.434
R13 Y Y.n0 171.29
R14 Y.n2 Y.t3 136.697
R15 Y.n3 Y.n1 50.795
R16 Y.n0 Y.t1 42.355
R17 Y.n1 Y.t4 39.692
R18 Y.n1 Y.t5 26.769
R19 Y.n0 Y.t2 26.595
R20 Y Y.n3 0.566
R21 Y.n3 Y.n2 0.446
R22 VGND.n2 VGND.n0 111.443
R23 VGND.n2 VGND.n1 110.657
R24 VGND.n0 VGND.t2 39.692
R25 VGND.n0 VGND.t3 24.923
R26 VGND.n1 VGND.t0 24.923
R27 VGND.n1 VGND.t1 24.923
R28 VGND VGND.n2 0.141
R29 VNB VNB.t4 6053.91
R30 VNB.t0 VNB.t2 4545.05
R31 VNB.t7 VNB.t6 2465.93
R32 VNB.t6 VNB.t5 2417.58
R33 VNB.t2 VNB.t7 2175.82
R34 VNB.t1 VNB.t0 2030.77
R35 VNB.t3 VNB.t1 2030.77
R36 VNB.t4 VNB.t3 2030.77
R37 A1.n3 A1.t0 212.079
R38 A1.n0 A1.t2 212.079
R39 A1.n0 A1.t3 139.779
R40 A1.n1 A1.t1 139.779
R41 A1 A1.n2 78.27
R42 A1.n4 A1.n3 76
R43 A1.n1 A1.n0 65.726
R44 A1.n2 A1.n1 13.145
R45 A1 A1.n4 6.606
R46 A1.n4 A1 3.303
R47 a_27_297.t3 a_27_297.n5 260.426
R48 a_27_297.n3 a_27_297.t1 242.31
R49 a_27_297.n4 a_27_297.n1 152.468
R50 a_27_297.n3 a_27_297.n2 152.468
R51 a_27_297.n5 a_27_297.n0 140.119
R52 a_27_297.n5 a_27_297.n4 123.699
R53 a_27_297.n4 a_27_297.n3 63.247
R54 a_27_297.n0 a_27_297.t6 44.325
R55 a_27_297.n2 a_27_297.t0 26.595
R56 a_27_297.n2 a_27_297.t5 26.595
R57 a_27_297.n1 a_27_297.t7 26.595
R58 a_27_297.n1 a_27_297.t4 26.595
R59 a_27_297.n0 a_27_297.t2 26.595
R60 VPWR.n7 VPWR.n6 312.281
R61 VPWR.n12 VPWR.n11 312.281
R62 VPWR.n3 VPWR.n2 294.905
R63 VPWR.n1 VPWR.n0 292.5
R64 VPWR.n0 VPWR.t5 49.25
R65 VPWR.n2 VPWR.t4 45.31
R66 VPWR.n6 VPWR.t2 26.595
R67 VPWR.n6 VPWR.t0 26.595
R68 VPWR.n11 VPWR.t3 26.595
R69 VPWR.n11 VPWR.t1 26.595
R70 VPWR.n5 VPWR.n4 4.65
R71 VPWR.n8 VPWR.n7 4.65
R72 VPWR.n10 VPWR.n9 4.65
R73 VPWR.n13 VPWR.n12 3.932
R74 VPWR.n3 VPWR.n1 2.41
R75 VPWR.n5 VPWR.n3 2.203
R76 VPWR.n13 VPWR.n10 0.137
R77 VPWR VPWR.n13 0.121
R78 VPWR.n8 VPWR.n5 0.119
R79 VPWR.n10 VPWR.n8 0.119
R80 VPB.t7 VPB.t6 574.143
R81 VPB.t6 VPB.t2 301.869
R82 VPB.t2 VPB.t3 295.95
R83 VPB.t4 VPB.t7 248.598
R84 VPB.t0 VPB.t4 248.598
R85 VPB.t5 VPB.t0 248.598
R86 VPB.t1 VPB.t5 248.598
R87 VPB VPB.t1 189.408
R88 A2.n2 A2.t1 212.079
R89 A2.n0 A2.t0 212.079
R90 A2.n2 A2.t3 139.779
R91 A2.n0 A2.t2 139.779
R92 A2 A2.n1 78.89
R93 A2.n3 A2.n2 76
R94 A2.n1 A2.n0 8.763
R95 A2.n3 A2 4.954
R96 A2 A2.n3 4.541
R97 a_277_47.n1 a_277_47.n0 289.658
R98 a_277_47.t1 a_277_47.n1 30.461
R99 a_277_47.n0 a_277_47.t3 24.923
R100 a_277_47.n0 a_277_47.t2 24.923
R101 a_277_47.n1 a_277_47.t0 24.923
R102 A3.n0 A3.t0 212.079
R103 A3.n1 A3.t2 212.079
R104 A3.n0 A3.t1 139.779
R105 A3.n1 A3.t3 139.779
R106 A3.n4 A3.n2 76
R107 A3.n2 A3.n0 41.627
R108 A3.n2 A3.n1 19.718
R109 A3.n4 A3.n3 7.432
R110 A3.n3 A3 1.961
R111 A3 A3.n4 0.103
R112 a_27_47.n0 a_27_47.t3 238.823
R113 a_27_47.n0 a_27_47.t0 238.823
R114 a_27_47.n1 a_27_47.n0 92.5
R115 a_27_47.n1 a_27_47.t2 24.923
R116 a_27_47.t1 a_27_47.n1 24.923
C0 A2 A1 0.14fF
C1 Y VGND 0.22fF
C2 A2 A3 0.14fF
C3 A1 Y 0.16fF
C4 Y B1 0.19fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__a31oi_4.ext - technology: sky130A

.subckt sky130_fd_sc_hd__a31oi_4 Y B1 A1 A3 A2 VPWR VGND VNB VPB
X0 a_27_47.t3 A2.t0 a_445_47.t4 VNB.t7 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 a_27_47.t2 A2.t1 a_445_47.t7 VNB.t6 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 VPWR.t11 A1.t0 a_27_297.t15 VPB.t15 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 a_27_297.t14 A1.t1 VPWR.t10 VPB.t14 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 a_27_297.t10 B1.t0 Y.t7 VPB.t10 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 VPWR.t6 A2.t2 a_27_297.t6 VPB.t6 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 a_27_297.t13 A1.t2 VPWR.t9 VPB.t13 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 a_27_297.t0 A3.t0 VPWR.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 VPWR.t8 A1.t3 a_27_297.t12 VPB.t12 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 Y.t6 B1.t1 a_27_297.t11 VPB.t11 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 a_27_297.t8 B1.t2 Y.t5 VPB.t8 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 a_445_47.t0 A1.t4 Y.t3 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 VPWR.t1 A3.t1 a_27_297.t1 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13 Y.t4 B1.t3 a_27_297.t9 VPB.t9 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14 a_445_47.t1 A1.t5 Y.t2 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X15 VGND.t7 B1.t4 Y.t11 VNB.t13 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X16 a_27_297.t2 A3.t2 VPWR.t2 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17 a_27_47.t4 A3.t3 VGND.t3 VNB.t10 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X18 a_27_47.t5 A3.t4 VGND.t2 VNB.t11 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X19 Y.t1 A1.t6 a_445_47.t2 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X20 a_27_297.t5 A2.t3 VPWR.t5 VPB.t5 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X21 Y.t0 A1.t7 a_445_47.t3 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X22 Y.t10 B1.t5 VGND.t6 VNB.t14 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X23 Y.t9 B1.t6 VGND.t5 VNB.t8 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X24 VGND.t1 A3.t5 a_27_47.t6 VNB.t12 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X25 a_445_47.t6 A2.t4 a_27_47.t1 VNB.t5 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X26 VPWR.t4 A2.t5 a_27_297.t4 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X27 a_445_47.t5 A2.t6 a_27_47.t0 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X28 a_27_297.t3 A2.t7 VPWR.t3 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X29 VGND.t4 B1.t7 Y.t8 VNB.t9 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X30 VPWR.t7 A3.t6 a_27_297.t7 VPB.t7 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X31 VGND.t0 A3.t7 a_27_47.t7 VNB.t15 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
R0 A2.n0 A2.t3 212.079
R1 A2.n2 A2.t5 212.079
R2 A2.n3 A2.t7 212.079
R3 A2.n4 A2.t2 212.079
R4 A2.n0 A2.t1 139.779
R5 A2.n2 A2.t6 139.779
R6 A2.n3 A2.t0 139.779
R7 A2.n4 A2.t4 139.779
R8 A2.n11 A2.n1 76
R9 A2.n10 A2.n9 76
R10 A2.n8 A2.n7 76
R11 A2.n6 A2.n5 76
R12 A2.n9 A2.n8 54.042
R13 A2.n5 A2.n3 52.581
R14 A2.n11 A2.n10 14.351
R15 A2.n1 A2.n0 13.145
R16 A2.n7 A2 12.8
R17 A2 A2.n6 9.309
R18 A2.n5 A2.n4 8.763
R19 A2.n6 A2 8.533
R20 A2.n9 A2.n2 5.842
R21 A2.n7 A2 5.042
R22 A2 A2.n11 1.939
R23 A2.n10 A2 1.551
R24 A2.n8 A2.n3 1.46
R25 a_445_47.n5 a_445_47.n4 155.747
R26 a_445_47.n3 a_445_47.n2 155.747
R27 a_445_47.n4 a_445_47.n3 102.4
R28 a_445_47.n4 a_445_47.n0 92.5
R29 a_445_47.n3 a_445_47.n1 92.5
R30 a_445_47.n2 a_445_47.t4 24.923
R31 a_445_47.n2 a_445_47.t6 24.923
R32 a_445_47.n1 a_445_47.t7 24.923
R33 a_445_47.n1 a_445_47.t5 24.923
R34 a_445_47.n0 a_445_47.t3 24.923
R35 a_445_47.n0 a_445_47.t1 24.923
R36 a_445_47.n5 a_445_47.t2 24.923
R37 a_445_47.t0 a_445_47.n5 24.923
R38 a_27_47.n2 a_27_47.t7 236.55
R39 a_27_47.n4 a_27_47.t2 229.593
R40 a_27_47.n2 a_27_47.n1 108.688
R41 a_27_47.n3 a_27_47.n0 108.688
R42 a_27_47.n5 a_27_47.n4 92.5
R43 a_27_47.n4 a_27_47.n3 63.247
R44 a_27_47.n3 a_27_47.n2 63.247
R45 a_27_47.n1 a_27_47.t6 24.923
R46 a_27_47.n1 a_27_47.t4 24.923
R47 a_27_47.n0 a_27_47.t1 24.923
R48 a_27_47.n0 a_27_47.t5 24.923
R49 a_27_47.n5 a_27_47.t0 24.923
R50 a_27_47.t3 a_27_47.n5 24.923
R51 VNB VNB.t15 6053.91
R52 VNB.t6 VNB.t1 4545.05
R53 VNB.t9 VNB.t8 2030.77
R54 VNB.t14 VNB.t9 2030.77
R55 VNB.t13 VNB.t14 2030.77
R56 VNB.t2 VNB.t13 2030.77
R57 VNB.t0 VNB.t2 2030.77
R58 VNB.t3 VNB.t0 2030.77
R59 VNB.t1 VNB.t3 2030.77
R60 VNB.t4 VNB.t6 2030.77
R61 VNB.t7 VNB.t4 2030.77
R62 VNB.t5 VNB.t7 2030.77
R63 VNB.t11 VNB.t5 2030.77
R64 VNB.t12 VNB.t11 2030.77
R65 VNB.t10 VNB.t12 2030.77
R66 VNB.t15 VNB.t10 2030.77
R67 A1.n8 A1.t3 213.914
R68 A1.n1 A1.t1 205.652
R69 A1.n5 A1.t0 205.652
R70 A1.n11 A1.t2 205.652
R71 A1.n0 A1.t6 204.047
R72 A1.n0 A1.t4 150.752
R73 A1.n10 A1.t5 139.779
R74 A1.n4 A1.t7 139.779
R75 A1.n3 A1.n2 76
R76 A1.n7 A1.n6 76
R77 A1.n13 A1.n12 76
R78 A1.n9 A1.n8 76
R79 A1.n4 A1.n3 34.428
R80 A1.n13 A1.n9 14.351
R81 A1 A1.n7 13.187
R82 A1.n3 A1.n1 12.394
R83 A1.n5 A1.n4 11.017
R84 A1.n2 A1 9.696
R85 A1.n12 A1.n10 9.64
R86 A1.n2 A1 8.145
R87 A1.n1 A1.n0 6.55
R88 A1.n6 A1.n5 5.508
R89 A1.n7 A1 4.654
R90 A1.n9 A1 2.327
R91 A1.n12 A1.n11 1.377
R92 A1 A1.n13 1.163
R93 a_27_297.n4 a_27_297.n3 292.5
R94 a_27_297.n11 a_27_297.t7 264.436
R95 a_27_297.n4 a_27_297.t10 190.107
R96 a_27_297.n7 a_27_297.n2 174.594
R97 a_27_297.n8 a_27_297.n1 174.594
R98 a_27_297.n9 a_27_297.n0 174.594
R99 a_27_297.n11 a_27_297.n10 174.594
R100 a_27_297.n13 a_27_297.n12 174.593
R101 a_27_297.n6 a_27_297.n5 138.16
R102 a_27_297.n5 a_27_297.t9 125.095
R103 a_27_297.n6 a_27_297.n4 117.076
R104 a_27_297.n7 a_27_297.n6 89.593
R105 a_27_297.n8 a_27_297.n7 64.752
R106 a_27_297.n9 a_27_297.n8 63.247
R107 a_27_297.n12 a_27_297.n9 63.247
R108 a_27_297.n12 a_27_297.n11 63.247
R109 a_27_297.n1 a_27_297.t12 30.535
R110 a_27_297.n5 a_27_297.t14 26.595
R111 a_27_297.n3 a_27_297.t11 26.595
R112 a_27_297.n3 a_27_297.t8 26.595
R113 a_27_297.n2 a_27_297.t15 26.595
R114 a_27_297.n2 a_27_297.t13 26.595
R115 a_27_297.n1 a_27_297.t5 26.595
R116 a_27_297.n0 a_27_297.t4 26.595
R117 a_27_297.n0 a_27_297.t3 26.595
R118 a_27_297.n10 a_27_297.t1 26.595
R119 a_27_297.n10 a_27_297.t2 26.595
R120 a_27_297.n13 a_27_297.t6 26.595
R121 a_27_297.t0 a_27_297.n13 26.595
R122 VPWR.n3 VPWR.n2 310.697
R123 VPWR.n1 VPWR.n0 164.214
R124 VPWR.n7 VPWR.n6 164.214
R125 VPWR.n11 VPWR.n10 164.214
R126 VPWR.n17 VPWR.n16 164.214
R127 VPWR.n22 VPWR.n21 164.214
R128 VPWR.n2 VPWR.t10 26.595
R129 VPWR.n2 VPWR.t11 26.595
R130 VPWR.n0 VPWR.t9 26.595
R131 VPWR.n0 VPWR.t8 26.595
R132 VPWR.n6 VPWR.t5 26.595
R133 VPWR.n6 VPWR.t4 26.595
R134 VPWR.n10 VPWR.t3 26.595
R135 VPWR.n10 VPWR.t6 26.595
R136 VPWR.n16 VPWR.t0 26.595
R137 VPWR.n16 VPWR.t1 26.595
R138 VPWR.n21 VPWR.t2 26.595
R139 VPWR.n21 VPWR.t7 26.595
R140 VPWR.n5 VPWR.n4 4.65
R141 VPWR.n9 VPWR.n8 4.65
R142 VPWR.n13 VPWR.n12 4.65
R143 VPWR.n15 VPWR.n14 4.65
R144 VPWR.n18 VPWR.n17 4.65
R145 VPWR.n20 VPWR.n19 4.65
R146 VPWR.n23 VPWR.n22 3.932
R147 VPWR.n3 VPWR.n1 3.407
R148 VPWR.n8 VPWR.n7 3.388
R149 VPWR.n12 VPWR.n11 0.376
R150 VPWR.n5 VPWR.n3 0.267
R151 VPWR.n23 VPWR.n20 0.137
R152 VPWR VPWR.n23 0.121
R153 VPWR.n9 VPWR.n5 0.119
R154 VPWR.n13 VPWR.n9 0.119
R155 VPWR.n15 VPWR.n13 0.119
R156 VPWR.n18 VPWR.n15 0.119
R157 VPWR.n20 VPWR.n18 0.119
R158 VPB.t14 VPB.t9 544.548
R159 VPB.t5 VPB.t12 260.436
R160 VPB.t11 VPB.t10 248.598
R161 VPB.t8 VPB.t11 248.598
R162 VPB.t9 VPB.t8 248.598
R163 VPB.t15 VPB.t14 248.598
R164 VPB.t13 VPB.t15 248.598
R165 VPB.t12 VPB.t13 248.598
R166 VPB.t4 VPB.t5 248.598
R167 VPB.t3 VPB.t4 248.598
R168 VPB.t6 VPB.t3 248.598
R169 VPB.t0 VPB.t6 248.598
R170 VPB.t1 VPB.t0 248.598
R171 VPB.t2 VPB.t1 248.598
R172 VPB.t7 VPB.t2 248.598
R173 VPB VPB.t7 189.408
R174 B1.n6 B1.t3 212.079
R175 B1.n1 B1.t0 212.079
R176 B1.n2 B1.t1 212.079
R177 B1.n0 B1.t2 212.079
R178 B1.n6 B1.t4 139.779
R179 B1.n1 B1.t6 139.779
R180 B1.n2 B1.t7 139.779
R181 B1.n0 B1.t5 139.779
R182 B1 B1.n3 79.225
R183 B1.n5 B1.n4 76
R184 B1.n7 B1.n6 76
R185 B1.n2 B1.n1 61.345
R186 B1.n6 B1.n5 54.042
R187 B1.n3 B1.n0 46.739
R188 B1.n3 B1.n2 14.606
R189 B1.n5 B1.n0 7.303
R190 B1 B1.n7 6.853
R191 B1.n4 B1 5.039
R192 B1.n4 B1 4.233
R193 B1.n7 B1 2.418
R194 Y.n2 Y.n0 353.111
R195 Y.n2 Y.n1 292.5
R196 Y.n6 Y.t2 229.593
R197 Y.n9 Y.t9 180.388
R198 Y.n8 Y.n3 108.688
R199 Y.n6 Y.n5 92.5
R200 Y.n7 Y.n4 92.5
R201 Y.n8 Y.n7 63.247
R202 Y.n7 Y.n6 63.247
R203 Y.n9 Y.n8 28.988
R204 Y.n0 Y.t5 26.595
R205 Y.n0 Y.t4 26.595
R206 Y.n1 Y.t7 26.595
R207 Y.n1 Y.t6 26.595
R208 Y.n4 Y.t11 24.923
R209 Y.n4 Y.t1 24.923
R210 Y.n5 Y.t3 24.923
R211 Y.n5 Y.t0 24.923
R212 Y.n3 Y.t8 24.923
R213 Y.n3 Y.t10 24.923
R214 Y Y.n2 13.76
R215 Y Y.n9 2.88
R216 A3.n1 A3.t0 212.079
R217 A3.n3 A3.t1 212.079
R218 A3.n0 A3.t2 212.079
R219 A3.n9 A3.t6 212.079
R220 A3.n1 A3.t4 139.779
R221 A3.n3 A3.t5 139.779
R222 A3.n0 A3.t3 139.779
R223 A3.n9 A3.t7 139.779
R224 A3.n10 A3.n9 103.021
R225 A3.n5 A3.n4 76
R226 A3.n8 A3.n7 76
R227 A3.n4 A3.n1 48.93
R228 A3.n3 A3.n2 41.627
R229 A3.n8 A3.n0 34.324
R230 A3.n9 A3.n8 27.021
R231 A3.n2 A3.n0 19.718
R232 A3.n7 A3.n6 14.351
R233 A3 A3.n5 12.606
R234 A3.n10 A3 12.606
R235 A3.n4 A3.n3 12.415
R236 A3.n5 A3 5.236
R237 A3 A3.n10 5.236
R238 A3.n6 A3 1.745
R239 A3.n7 A3 1.745
R240 VGND.n3 VGND.n0 110.725
R241 VGND.n2 VGND.n1 107.239
R242 VGND.n23 VGND.n22 107.239
R243 VGND.n28 VGND.n27 107.239
R244 VGND.n0 VGND.t5 24.923
R245 VGND.n0 VGND.t4 24.923
R246 VGND.n1 VGND.t6 24.923
R247 VGND.n1 VGND.t7 24.923
R248 VGND.n22 VGND.t2 24.923
R249 VGND.n22 VGND.t1 24.923
R250 VGND.n27 VGND.t3 24.923
R251 VGND.n27 VGND.t0 24.923
R252 VGND.n5 VGND.n4 4.65
R253 VGND.n7 VGND.n6 4.65
R254 VGND.n9 VGND.n8 4.65
R255 VGND.n11 VGND.n10 4.65
R256 VGND.n13 VGND.n12 4.65
R257 VGND.n15 VGND.n14 4.65
R258 VGND.n17 VGND.n16 4.65
R259 VGND.n19 VGND.n18 4.65
R260 VGND.n21 VGND.n20 4.65
R261 VGND.n24 VGND.n23 4.65
R262 VGND.n26 VGND.n25 4.65
R263 VGND.n29 VGND.n28 3.932
R264 VGND.n3 VGND.n2 3.759
R265 VGND.n5 VGND.n3 0.254
R266 VGND.n29 VGND.n26 0.137
R267 VGND VGND.n29 0.121
R268 VGND.n7 VGND.n5 0.119
R269 VGND.n9 VGND.n7 0.119
R270 VGND.n11 VGND.n9 0.119
R271 VGND.n13 VGND.n11 0.119
R272 VGND.n15 VGND.n13 0.119
R273 VGND.n17 VGND.n15 0.119
R274 VGND.n19 VGND.n17 0.119
R275 VGND.n21 VGND.n19 0.119
R276 VGND.n24 VGND.n21 0.119
R277 VGND.n26 VGND.n24 0.119
C0 Y B1 0.34fF
C1 Y A1 0.24fF
C2 VPB VPWR 0.15fF
C3 A3 A2 0.10fF
C4 VGND Y 0.34fF
C5 VGND VPWR 0.17fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__a32o_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__a32o_1 X A3 B2 B1 A1 A2 VGND VPWR VNB VPB
X0 a_93_21.t0 A1.t0 a_346_47.t0 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 a_93_21.t1 B1.t0 a_250_297.t2 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 a_584_47.t0 B1.t1 a_93_21.t2 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 VPWR.t1 a_93_21.t4 X.t1 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 VGND.t2 B2.t0 a_584_47.t1 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 a_256_47.t0 A3.t0 VGND.t1 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 a_250_297.t3 B2.t1 a_93_21.t3 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 VGND.t0 a_93_21.t5 X.t0 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 a_250_297.t4 A3.t1 VPWR.t3 VPB.t5 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 VPWR.t0 A2.t0 a_250_297.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 a_250_297.t1 A1.t1 VPWR.t2 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 a_346_47.t1 A2.t1 a_256_47.t1 VNB.t5 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
R0 A1.n0 A1.t1 241.534
R1 A1.n0 A1.t0 169.234
R2 A1 A1.n0 78.427
R3 a_346_47.t0 a_346_47.t1 83.076
R4 a_93_21.n3 a_93_21.n2 500.082
R5 a_93_21.n2 a_93_21.n1 257.164
R6 a_93_21.n0 a_93_21.t4 236.549
R7 a_93_21.n0 a_93_21.t5 164.249
R8 a_93_21.n2 a_93_21.n0 76
R9 a_93_21.n1 a_93_21.t2 41.538
R10 a_93_21.n1 a_93_21.t0 39.692
R11 a_93_21.n3 a_93_21.t3 27.58
R12 a_93_21.t1 a_93_21.n3 27.58
R13 VNB VNB.t0 6392.37
R14 VNB.t0 VNB.t4 3215.38
R15 VNB.t5 VNB.t1 2901.1
R16 VNB.t1 VNB.t3 2852.75
R17 VNB.t4 VNB.t5 2175.82
R18 VNB.t3 VNB.t2 1740.66
R19 B1.n0 B1.t0 241.534
R20 B1.n0 B1.t1 169.234
R21 B1 B1.n0 77.676
R22 a_250_297.n1 a_250_297.t3 243.969
R23 a_250_297.n2 a_250_297.n1 218.959
R24 a_250_297.n1 a_250_297.n0 143.026
R25 a_250_297.n0 a_250_297.t2 37.43
R26 a_250_297.n0 a_250_297.t1 35.46
R27 a_250_297.t0 a_250_297.n2 32.505
R28 a_250_297.n2 a_250_297.t4 32.505
R29 VPB.t1 VPB.t5 375.856
R30 VPB.t0 VPB.t2 355.14
R31 VPB.t2 VPB.t3 307.788
R32 VPB.t5 VPB.t0 284.112
R33 VPB.t3 VPB.t4 254.517
R34 VPB VPB.t1 230.841
R35 a_584_47.t0 a_584_47.t1 38.769
R36 X.n4 X.n3 292.5
R37 X.n5 X.n4 147.091
R38 X X.n0 94.028
R39 X.n2 X.n0 92.5
R40 X.n4 X.t1 40.385
R41 X.n0 X.t0 37.846
R42 X.n3 X 10.792
R43 X.n2 X.n1 8.282
R44 X.n1 X 6.776
R45 X.n6 X 6.525
R46 X.n3 X 6.274
R47 X.n6 X.n5 5.584
R48 X.n1 X 5.158
R49 X X.n6 4.967
R50 X.n5 X 2.402
R51 X X.n2 2.007
R52 VPWR.n2 VPWR.n1 310.847
R53 VPWR.n2 VPWR.n0 167.413
R54 VPWR.n0 VPWR.t3 51.22
R55 VPWR.n1 VPWR.t2 44.325
R56 VPWR.n1 VPWR.t0 44.325
R57 VPWR.n0 VPWR.t1 44.325
R58 VPWR VPWR.n2 0.178
R59 B2.n0 B2.t1 241.534
R60 B2.n0 B2.t0 169.234
R61 B2.n1 B2.n0 76
R62 B2 B2.n1 13.526
R63 B2.n1 B2 2.011
R64 VGND.n1 VGND.n0 111.392
R65 VGND.n1 VGND.t2 107.332
R66 VGND.n0 VGND.t1 68.307
R67 VGND.n0 VGND.t0 26.769
R68 VGND VGND.n1 0.149
R69 A3.n0 A3.t1 241.534
R70 A3.n0 A3.t0 169.234
R71 A3 A3.n0 82.4
R72 a_256_47.t0 a_256_47.t1 55.384
R73 A2.n0 A2.t0 241.534
R74 A2.n0 A2.t1 169.234
R75 A2 A2.n0 78.607
C0 VPWR X 0.12fF
C1 A1 B1 0.15fF
C2 A1 A2 0.14fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__a32o_2.ext - technology: sky130A

.subckt sky130_fd_sc_hd__a32o_2 B2 X A2 A3 A1 B1 VGND VPWR VNB VPB
X0 VPWR.t2 A3.t0 a_299_297.t0 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_299_297.t2 A2.t0 VPWR.t3 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 a_352_47.t1 B2.t0 VGND.t3 VNB.t5 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 a_549_47.t1 A1.t0 a_21_199.t1 VNB.t6 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 X.t1 a_21_199.t4 VPWR.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 VGND.t0 a_21_199.t5 X.t3 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 a_665_47.t1 A2.t1 a_549_47.t0 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 VPWR.t4 A1.t1 a_299_297.t4 VPB.t6 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 a_299_297.t3 B1.t0 a_21_199.t2 VPB.t5 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 a_21_199.t3 B2.t1 a_299_297.t1 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 VGND.t2 A3.t1 a_665_47.t0 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 VPWR.t1 a_21_199.t6 X.t0 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 X.t2 a_21_199.t7 VGND.t1 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 a_21_199.t0 B1.t1 a_352_47.t0 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
R0 A3.n0 A3.t0 230.154
R1 A3.n0 A3.t1 157.854
R2 A3.n1 A3.n0 76
R3 A3.n1 A3 15.2
R4 A3 A3.n1 2.933
R5 a_299_297.n1 a_299_297.t1 254.228
R6 a_299_297.n2 a_299_297.n1 239.509
R7 a_299_297.n1 a_299_297.n0 140.292
R8 a_299_297.n0 a_299_297.t4 26.595
R9 a_299_297.n0 a_299_297.t3 26.595
R10 a_299_297.t0 a_299_297.n2 26.595
R11 a_299_297.n2 a_299_297.t2 26.595
R12 VPWR.n12 VPWR.n11 312.281
R13 VPWR.n1 VPWR.n0 311.7
R14 VPWR.n2 VPWR.t2 194.535
R15 VPWR.n0 VPWR.t3 58.115
R16 VPWR.n0 VPWR.t4 26.595
R17 VPWR.n11 VPWR.t0 26.595
R18 VPWR.n11 VPWR.t1 26.595
R19 VPWR.n4 VPWR.n3 4.65
R20 VPWR.n6 VPWR.n5 4.65
R21 VPWR.n8 VPWR.n7 4.65
R22 VPWR.n10 VPWR.n9 4.65
R23 VPWR.n2 VPWR.n1 3.995
R24 VPWR.n13 VPWR.n12 3.932
R25 VPWR.n4 VPWR.n2 0.223
R26 VPWR.n13 VPWR.n10 0.137
R27 VPWR VPWR.n13 0.121
R28 VPWR.n6 VPWR.n4 0.119
R29 VPWR.n8 VPWR.n6 0.119
R30 VPWR.n10 VPWR.n8 0.119
R31 VPB.t0 VPB.t3 556.386
R32 VPB.t6 VPB.t4 343.302
R33 VPB.t4 VPB.t2 248.598
R34 VPB.t5 VPB.t6 248.598
R35 VPB.t3 VPB.t5 248.598
R36 VPB.t1 VPB.t0 248.598
R37 VPB VPB.t1 189.408
R38 A2.n0 A2.t0 241.534
R39 A2.n0 A2.t1 169.234
R40 A2.n1 A2.n0 76
R41 A2.n1 A2 11.957
R42 A2 A2.n1 1.852
R43 B2.n0 B2.t1 233.257
R44 B2.n0 B2.t0 139.779
R45 B2 B2.n0 124.435
R46 VGND.n9 VGND.t1 190.095
R47 VGND.n2 VGND.t2 107.68
R48 VGND.n1 VGND.n0 92.5
R49 VGND.n4 VGND.n3 92.5
R50 VGND.n0 VGND.t3 24.923
R51 VGND.n3 VGND.t0 24.923
R52 VGND.n2 VGND.n1 7.381
R53 VGND.n10 VGND.n9 4.65
R54 VGND.n6 VGND.n5 4.65
R55 VGND.n8 VGND.n7 4.65
R56 VGND.n5 VGND.n4 1.207
R57 VGND.n6 VGND.n2 0.134
R58 VGND.n8 VGND.n6 0.119
R59 VGND.n10 VGND.n8 0.119
R60 VGND VGND.n10 0.02
R61 a_352_47.t0 a_352_47.t1 65.538
R62 VNB VNB.t1 6053.91
R63 VNB.t0 VNB.t5 3843.96
R64 VNB.t6 VNB.t3 2804.4
R65 VNB.t5 VNB.t4 2441.76
R66 VNB.t4 VNB.t6 2320.88
R67 VNB.t3 VNB.t2 2030.77
R68 VNB.t1 VNB.t0 2030.77
R69 A1.n0 A1.t1 237.733
R70 A1.n0 A1.t0 165.433
R71 A1.n1 A1.n0 109.511
R72 A1 A1.n1 9.066
R73 A1.n1 A1 4.73
R74 a_21_199.n1 a_21_199.t4 212.079
R75 a_21_199.n2 a_21_199.t6 212.079
R76 a_21_199.n4 a_21_199.n3 185.927
R77 a_21_199.n5 a_21_199.n4 167.402
R78 a_21_199.n1 a_21_199.t5 139.779
R79 a_21_199.n2 a_21_199.t7 139.779
R80 a_21_199.n4 a_21_199.n0 126.999
R81 a_21_199.n3 a_21_199.n1 39.436
R82 a_21_199.n0 a_21_199.t1 32.307
R83 a_21_199.n0 a_21_199.t0 28.615
R84 a_21_199.t2 a_21_199.n5 26.595
R85 a_21_199.n5 a_21_199.t3 26.595
R86 a_21_199.n3 a_21_199.n2 21.909
R87 a_549_47.t0 a_549_47.t1 79.384
R88 X.n1 X.t1 235.91
R89 X.n0 X.t0 172.846
R90 X X.n2 119.246
R91 X.n2 X.t3 24.923
R92 X.n2 X.t2 24.923
R93 X.n1 X.n0 10.022
R94 X.n0 X 5.334
R95 X X.n1 5.18
R96 a_665_47.t0 a_665_47.t1 49.846
R97 B1.n0 B1.t0 241.534
R98 B1.n0 B1.t1 169.234
R99 B1 B1.n0 110.257
C0 X VPWR 0.24fF
C1 A2 A1 0.16fF
C2 A2 A3 0.11fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__a32o_4.ext - technology: sky130A

.subckt sky130_fd_sc_hd__a32o_4 A3 X A2 B1 B2 A1 VGND VPWR VNB VPB
X0 VGND.t7 A3.t0 a_445_47.t2 VNB.t13 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 a_445_297.t7 A2.t0 VPWR.t7 VPB.t11 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 VPWR.t6 A2.t1 a_445_297.t6 VPB.t10 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 a_635_47.t3 A2.t2 a_445_47.t0 VNB.t7 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 a_445_297.t9 A3.t1 VPWR.t9 VPB.t13 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 VPWR.t4 a_79_21.t8 X.t7 VPB.t6 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 a_445_297.t0 B2.t0 a_79_21.t2 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 a_79_21.t4 B1.t0 a_1142_47.t1 VNB.t9 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 a_79_21.t3 B2.t1 a_445_297.t1 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 X.t6 a_79_21.t9 VPWR.t5 VPB.t7 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 a_445_47.t1 A2.t3 a_635_47.t2 VNB.t8 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 a_79_21.t0 A1.t0 a_635_47.t0 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 VPWR.t0 a_79_21.t10 X.t5 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13 a_445_297.t4 B1.t1 a_79_21.t5 VPB.t8 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14 VGND.t0 a_79_21.t11 X.t3 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X15 VGND.t1 a_79_21.t12 X.t2 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X16 a_1142_47.t0 B1.t2 a_79_21.t6 VNB.t10 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X17 VGND.t4 B2.t2 a_1142_47.t3 VNB.t6 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X18 a_635_47.t1 A1.t1 a_79_21.t1 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X19 X.t1 a_79_21.t13 VGND.t2 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X20 a_445_47.t3 A3.t2 VGND.t6 VNB.t12 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X21 a_79_21.t7 B1.t3 a_445_297.t5 VPB.t9 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X22 a_1142_47.t2 B2.t3 VGND.t5 VNB.t11 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X23 VPWR.t8 A3.t3 a_445_297.t8 VPB.t12 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X24 a_445_297.t2 A1.t2 VPWR.t2 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X25 X.t4 a_79_21.t14 VPWR.t1 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X26 VPWR.t3 A1.t3 a_445_297.t3 VPB.t5 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X27 X.t0 a_79_21.t15 VGND.t3 VNB.t5 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
R0 A3.n0 A3.t3 212.079
R1 A3.n1 A3.t1 212.079
R2 A3.n0 A3.t0 139.779
R3 A3.n1 A3.t2 139.779
R4 A3.n3 A3.n0 97.279
R5 A3 A3.n2 80.363
R6 A3.n2 A3.n1 32.863
R7 A3.n2 A3.n0 28.481
R8 A3.n3 A3 15.418
R9 A3 A3.n3 11.345
R10 a_445_47.n1 a_445_47.n0 305.094
R11 a_445_47.n0 a_445_47.t2 24.923
R12 a_445_47.n0 a_445_47.t3 24.923
R13 a_445_47.t0 a_445_47.n1 24.923
R14 a_445_47.n1 a_445_47.t1 24.923
R15 VGND.n1 VGND.t7 190.315
R16 VGND.n15 VGND.t3 190.315
R17 VGND.n2 VGND.n0 111.717
R18 VGND.n6 VGND.n5 107.239
R19 VGND.n11 VGND.n10 107.239
R20 VGND.n0 VGND.t5 24.923
R21 VGND.n0 VGND.t4 24.923
R22 VGND.n5 VGND.t6 24.923
R23 VGND.n5 VGND.t1 24.923
R24 VGND.n10 VGND.t2 24.923
R25 VGND.n10 VGND.t0 24.923
R26 VGND.n2 VGND.n1 7.528
R27 VGND.n16 VGND.n15 4.65
R28 VGND.n4 VGND.n3 4.65
R29 VGND.n7 VGND.n6 4.65
R30 VGND.n9 VGND.n8 4.65
R31 VGND.n12 VGND.n11 4.65
R32 VGND.n14 VGND.n13 4.65
R33 VGND.n4 VGND.n2 0.134
R34 VGND.n7 VGND.n4 0.119
R35 VGND.n9 VGND.n7 0.119
R36 VGND.n12 VGND.n9 0.119
R37 VGND.n14 VGND.n12 0.119
R38 VGND.n16 VGND.n14 0.119
R39 VGND VGND.n16 0.02
R40 VNB.t1 VNB.t9 6164.83
R41 VNB VNB.t5 6053.91
R42 VNB.t13 VNB.t8 4545.05
R43 VNB.t10 VNB.t6 2248.35
R44 VNB.t6 VNB.t11 2030.77
R45 VNB.t9 VNB.t10 2030.77
R46 VNB.t0 VNB.t1 2030.77
R47 VNB.t7 VNB.t0 2030.77
R48 VNB.t8 VNB.t7 2030.77
R49 VNB.t12 VNB.t13 2030.77
R50 VNB.t3 VNB.t12 2030.77
R51 VNB.t4 VNB.t3 2030.77
R52 VNB.t2 VNB.t4 2030.77
R53 VNB.t5 VNB.t2 2030.77
R54 A2.n0 A2.t0 205.652
R55 A2.n2 A2.t1 205.652
R56 A2.n0 A2.t2 139.779
R57 A2.n2 A2.t3 139.779
R58 A2.n3 A2.n2 77.377
R59 A2.n4 A2.n1 76
R60 A2.n4 A2.n3 17.408
R61 A2.n1 A2.n0 12.394
R62 A2.n3 A2 5.632
R63 A2 A2.n4 0.512
R64 VPWR.n6 VPWR.t8 576.219
R65 VPWR.n3 VPWR.n0 311.04
R66 VPWR.n2 VPWR.n1 307.239
R67 VPWR.n21 VPWR.t1 190.809
R68 VPWR.n17 VPWR.n16 164.214
R69 VPWR.n12 VPWR.n11 164.214
R70 VPWR.n16 VPWR.t5 26.595
R71 VPWR.n16 VPWR.t0 26.595
R72 VPWR.n11 VPWR.t9 26.595
R73 VPWR.n11 VPWR.t4 26.595
R74 VPWR.n1 VPWR.t7 26.595
R75 VPWR.n1 VPWR.t6 26.595
R76 VPWR.n0 VPWR.t2 26.595
R77 VPWR.n0 VPWR.t3 26.595
R78 VPWR.n3 VPWR.n2 5.687
R79 VPWR.n5 VPWR.n4 4.65
R80 VPWR.n8 VPWR.n7 4.65
R81 VPWR.n10 VPWR.n9 4.65
R82 VPWR.n13 VPWR.n12 4.65
R83 VPWR.n15 VPWR.n14 4.65
R84 VPWR.n18 VPWR.n17 4.65
R85 VPWR.n20 VPWR.n19 4.65
R86 VPWR.n22 VPWR.n21 4.65
R87 VPWR.n7 VPWR.n6 3.388
R88 VPWR.n5 VPWR.n3 0.461
R89 VPWR.n8 VPWR.n5 0.119
R90 VPWR.n10 VPWR.n8 0.119
R91 VPWR.n13 VPWR.n10 0.119
R92 VPWR.n15 VPWR.n13 0.119
R93 VPWR.n18 VPWR.n15 0.119
R94 VPWR.n20 VPWR.n18 0.119
R95 VPWR.n22 VPWR.n20 0.119
R96 VPWR VPWR.n22 0.02
R97 a_445_297.n5 a_445_297.t6 547.361
R98 a_445_297.n5 a_445_297.n4 379.464
R99 a_445_297.n7 a_445_297.n6 308.688
R100 a_445_297.n1 a_445_297.n0 292.5
R101 a_445_297.n3 a_445_297.n2 292.5
R102 a_445_297.n1 a_445_297.t0 234.878
R103 a_445_297.n2 a_445_297.t2 203.895
R104 a_445_297.n6 a_445_297.n3 143.811
R105 a_445_297.n3 a_445_297.n1 63.247
R106 a_445_297.n6 a_445_297.n5 63.247
R107 a_445_297.n2 a_445_297.t5 26.595
R108 a_445_297.n0 a_445_297.t1 26.595
R109 a_445_297.n0 a_445_297.t4 26.595
R110 a_445_297.n4 a_445_297.t8 26.595
R111 a_445_297.n4 a_445_297.t9 26.595
R112 a_445_297.n7 a_445_297.t3 26.595
R113 a_445_297.t7 a_445_297.n7 26.595
R114 VPB.t4 VPB.t9 781.308
R115 VPB.t12 VPB.t10 556.386
R116 VPB.t3 VPB.t2 248.598
R117 VPB.t8 VPB.t3 248.598
R118 VPB.t9 VPB.t8 248.598
R119 VPB.t5 VPB.t4 248.598
R120 VPB.t11 VPB.t5 248.598
R121 VPB.t10 VPB.t11 248.598
R122 VPB.t13 VPB.t12 248.598
R123 VPB.t6 VPB.t13 248.598
R124 VPB.t7 VPB.t6 248.598
R125 VPB.t0 VPB.t7 248.598
R126 VPB.t1 VPB.t0 248.598
R127 VPB VPB.t1 189.408
R128 a_635_47.n1 a_635_47.t1 238.823
R129 a_635_47.t2 a_635_47.n1 238.823
R130 a_635_47.n1 a_635_47.n0 92.5
R131 a_635_47.n0 a_635_47.t0 24.923
R132 a_635_47.n0 a_635_47.t3 24.923
R133 a_79_21.n15 a_79_21.n14 355.747
R134 a_79_21.n13 a_79_21.n12 293.829
R135 a_79_21.n14 a_79_21.n0 292.5
R136 a_79_21.n9 a_79_21.t8 212.079
R137 a_79_21.n10 a_79_21.t9 212.079
R138 a_79_21.n6 a_79_21.t10 212.079
R139 a_79_21.n4 a_79_21.t14 212.079
R140 a_79_21.n3 a_79_21.n1 159.511
R141 a_79_21.n3 a_79_21.n2 153.111
R142 a_79_21.n9 a_79_21.t12 139.779
R143 a_79_21.n10 a_79_21.t13 139.779
R144 a_79_21.n6 a_79_21.t11 139.779
R145 a_79_21.n4 a_79_21.t15 139.779
R146 a_79_21.n8 a_79_21.n5 90.351
R147 a_79_21.n14 a_79_21.n13 88.197
R148 a_79_21.n8 a_79_21.n7 76
R149 a_79_21.n12 a_79_21.n11 76
R150 a_79_21.n13 a_79_21.n3 51.952
R151 a_79_21.n11 a_79_21.n9 48.93
R152 a_79_21.n5 a_79_21.n4 27.021
R153 a_79_21.n0 a_79_21.t5 26.595
R154 a_79_21.n0 a_79_21.t7 26.595
R155 a_79_21.t2 a_79_21.n15 26.595
R156 a_79_21.n15 a_79_21.t3 26.595
R157 a_79_21.n1 a_79_21.t6 24.923
R158 a_79_21.n1 a_79_21.t4 24.923
R159 a_79_21.n2 a_79_21.t1 24.923
R160 a_79_21.n2 a_79_21.t0 24.923
R161 a_79_21.n7 a_79_21.n6 19.718
R162 a_79_21.n12 a_79_21.n8 14.351
R163 a_79_21.n11 a_79_21.n10 12.415
R164 X.n2 X.n1 237.841
R165 X.n2 X.n0 174.594
R166 X.n5 X.n4 171.935
R167 X.n5 X.n3 108.688
R168 X X.n2 33.454
R169 X X.n5 28.218
R170 X.n1 X.t7 26.595
R171 X.n1 X.t6 26.595
R172 X.n0 X.t5 26.595
R173 X.n0 X.t4 26.595
R174 X.n3 X.t3 24.923
R175 X.n3 X.t0 24.923
R176 X.n4 X.t2 24.923
R177 X.n4 X.t1 24.923
R178 B2.n1 B2.t0 260.279
R179 B2.n2 B2.t1 212.079
R180 B2.n0 B2.t3 192.799
R181 B2.n2 B2.t2 149.419
R182 B2.n0 B2 98.562
R183 B2.n4 B2.n3 76
R184 B2.n3 B2.n2 44.183
R185 B2.n4 B2 17.163
R186 B2.n3 B2.n1 11.246
R187 B2.n5 B2 9.846
R188 B2 B2.n5 4.945
R189 B2.n1 B2.n0 4.82
R190 B2.n5 B2.n4 4.654
R191 B1.n0 B1.t1 219.309
R192 B1.n3 B1.t3 212.079
R193 B1.n4 B1.t0 155.741
R194 B1.n0 B1.t2 149.419
R195 B1.n2 B1.n1 76
R196 B1.n5 B1.n4 76
R197 B1.n5 B1 9.774
R198 B1.n1 B1.n0 7.23
R199 B1 B1.n2 6.981
R200 B1.n2 B1 3.723
R201 B1.n4 B1.n3 1.606
R202 B1 B1.n5 0.93
R203 a_1142_47.n1 a_1142_47.t2 250.855
R204 a_1142_47.t1 a_1142_47.n1 242.211
R205 a_1142_47.n1 a_1142_47.n0 92.5
R206 a_1142_47.n0 a_1142_47.t0 33.23
R207 a_1142_47.n0 a_1142_47.t3 24.923
R208 A1.n0 A1.t2 257.066
R209 A1.n2 A1.t3 205.652
R210 A1.n1 A1.t1 192.799
R211 A1.n2 A1.t0 149.419
R212 A1 A1.n1 93.971
R213 A1.n4 A1.n3 76
R214 A1.n3 A1.n2 33.137
R215 A1.n4 A1 13.312
R216 A1 A1.n4 10.24
R217 A1.n1 A1.n0 8.033
C0 B1 B2 0.11fF
C1 VPB VPWR 0.15fF
C2 VPWR X 0.46fF
C3 VGND X 0.32fF
C4 VGND VPWR 0.16fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__a32oi_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__a32oi_1 A2 Y A1 B2 B1 A3 VGND VPWR VNB VPB
X0 VPWR.t2 A3.t0 a_27_297.t3 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 VGND.t1 A3.t1 a_383_47.t1 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 a_309_47.t1 A1.t0 Y.t2 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 Y.t0 B1.t0 a_109_47.t0 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 a_27_297.t0 B1.t1 Y.t1 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 a_383_47.t0 A2.t0 a_309_47.t0 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 a_27_297.t2 A2.t1 VPWR.t1 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 Y.t3 B2.t0 a_27_297.t4 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 VPWR.t0 A1.t1 a_27_297.t1 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 a_109_47.t1 B2.t1 VGND.t0 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
R0 A3.n0 A3.t0 212.152
R1 A3.n0 A3.t1 150.442
R2 A3 A3.n0 77.696
R3 a_27_297.n1 a_27_297.t4 237.294
R4 a_27_297.n1 a_27_297.n0 219.925
R5 a_27_297.n2 a_27_297.n1 140.946
R6 a_27_297.t0 a_27_297.n2 58.115
R7 a_27_297.n0 a_27_297.t3 28.565
R8 a_27_297.n0 a_27_297.t2 26.595
R9 a_27_297.n2 a_27_297.t1 26.595
R10 VPWR.n1 VPWR.n0 317.385
R11 VPWR.n1 VPWR.t2 148.772
R12 VPWR.n0 VPWR.t1 26.595
R13 VPWR.n0 VPWR.t0 26.595
R14 VPWR VPWR.n1 0.476
R15 VPB.t0 VPB.t1 343.302
R16 VPB.t2 VPB.t3 254.517
R17 VPB.t1 VPB.t2 248.598
R18 VPB.t4 VPB.t0 248.598
R19 VPB VPB.t4 192.367
R20 a_383_47.t0 a_383_47.t1 60.923
R21 VGND.n0 VGND.t0 194.195
R22 VGND.n0 VGND.t1 106.955
R23 VGND VGND.n0 0.044
R24 VNB VNB.t0 6078.09
R25 VNB.t1 VNB.t2 2997.8
R26 VNB.t3 VNB.t4 2320.88
R27 VNB.t0 VNB.t1 1837.36
R28 VNB.t2 VNB.t3 1789.01
R29 A1.n0 A1.t1 241.534
R30 A1.n0 A1.t0 169.234
R31 A1 A1.n0 117.116
R32 Y Y.n1 300.362
R33 Y Y.n0 199.733
R34 Y.n0 Y.t2 58.153
R35 Y.n0 Y.t0 28.615
R36 Y.n1 Y.t1 26.595
R37 Y.n1 Y.t3 26.595
R38 a_309_47.t0 a_309_47.t1 40.615
R39 B1.n0 B1.t1 236.932
R40 B1.n0 B1.t0 164.632
R41 B1 B1.n0 105.046
R42 a_109_47.t0 a_109_47.t1 42.461
R43 A2.n0 A2.t1 229.395
R44 A2.n0 A2.t0 164.236
R45 A2 A2.n0 79.684
R46 B2.n0 B2.t0 230.154
R47 B2.n0 B2.t1 157.854
R48 B2 B2.n0 79.684
C0 A2 A1 0.15fF
C1 B1 Y 0.15fF
C2 A2 A3 0.11fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__a32oi_2.ext - technology: sky130A

.subckt sky130_fd_sc_hd__a32oi_2 B2 A3 A2 A1 Y B1 VGND VPWR VNB VPB
X0 Y.t4 A1.t0 a_478_47.t3 VNB.t5 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 a_27_297.t6 A1.t1 VPWR.t3 VPB.t6 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 a_27_297.t3 A2.t0 VPWR.t0 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 a_27_297.t8 A3.t0 VPWR.t4 VPB.t8 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 VPWR.t5 A3.t1 a_27_297.t9 VPB.t9 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 VPWR.t2 A1.t2 a_27_297.t5 VPB.t5 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 a_27_297.t1 B1.t0 Y.t1 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 a_478_47.t2 A1.t3 Y.t3 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 a_478_47.t0 A2.t1 a_730_47.t1 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 VGND.t3 A3.t2 a_730_47.t3 VNB.t8 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 Y.t2 B1.t1 a_27_297.t2 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 a_27_297.t7 B2.t0 Y.t7 VPB.t7 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 a_27_47.t1 B2.t1 VGND.t0 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 a_27_47.t3 B1.t2 Y.t5 VNB.t6 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14 Y.t6 B1.t3 a_27_47.t2 VNB.t7 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X15 a_730_47.t2 A3.t3 VGND.t2 VNB.t9 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X16 Y.t0 B2.t2 a_27_297.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17 VPWR.t1 A2.t2 a_27_297.t4 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X18 VGND.t1 B2.t3 a_27_47.t0 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X19 a_730_47.t0 A2.t3 a_478_47.t1 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
R0 A1.n2 A1.t2 322.581
R1 A1.n0 A1.t1 221.719
R2 A1.n0 A1.t3 165.485
R3 A1.n1 A1.t0 149.419
R4 A1 A1.n0 79.374
R5 A1.n3 A1.n2 76
R6 A1.n3 A1 6.167
R7 A1 A1.n3 4.538
R8 A1.n2 A1.n1 1.785
R9 a_478_47.n1 a_478_47.t3 239.576
R10 a_478_47.t0 a_478_47.n1 238.823
R11 a_478_47.n1 a_478_47.n0 92.5
R12 a_478_47.n0 a_478_47.t2 26.769
R13 a_478_47.n0 a_478_47.t1 24.923
R14 Y.n2 Y.n0 317.723
R15 Y.n2 Y.n1 220.561
R16 Y.n5 Y.n4 149.347
R17 Y.n5 Y.n3 126.005
R18 Y Y.n2 39.16
R19 Y.n0 Y.t1 26.595
R20 Y.n0 Y.t2 26.595
R21 Y.n1 Y.t7 26.595
R22 Y.n1 Y.t0 26.595
R23 Y.n4 Y.t3 24.923
R24 Y.n4 Y.t4 24.923
R25 Y.n3 Y.t5 24.923
R26 Y.n3 Y.t6 24.923
R27 Y Y.n5 1.488
R28 VNB VNB.t1 6053.91
R29 VNB.t2 VNB.t9 4810.99
R30 VNB.t6 VNB.t5 4810.99
R31 VNB.t9 VNB.t8 2514.28
R32 VNB.t4 VNB.t3 2079.12
R33 VNB.t3 VNB.t2 2030.77
R34 VNB.t5 VNB.t4 2030.77
R35 VNB.t7 VNB.t6 2030.77
R36 VNB.t0 VNB.t7 2030.77
R37 VNB.t1 VNB.t0 2030.77
R38 VPWR.n19 VPWR.n18 292.5
R39 VPWR.n21 VPWR.n20 292.5
R40 VPWR.n3 VPWR.n2 292.5
R41 VPWR.n1 VPWR.n0 292.5
R42 VPWR.n11 VPWR.n10 292.5
R43 VPWR.n9 VPWR.n8 292.5
R44 VPWR.n20 VPWR.t2 41.37
R45 VPWR.n18 VPWR.t3 40.385
R46 VPWR.n0 VPWR.t4 32.505
R47 VPWR.n2 VPWR.t5 32.505
R48 VPWR.n8 VPWR.t0 26.595
R49 VPWR.n10 VPWR.t1 26.595
R50 VPWR.n22 VPWR.n19 5.701
R51 VPWR.n17 VPWR.n16 4.65
R52 VPWR.n5 VPWR.n4 4.65
R53 VPWR.n7 VPWR.n6 4.65
R54 VPWR.n13 VPWR.n12 4.65
R55 VPWR.n15 VPWR.n14 4.65
R56 VPWR.n23 VPWR.n22 4.65
R57 VPWR.n5 VPWR.n1 4.642
R58 VPWR.n12 VPWR.n11 4.538
R59 VPWR.n12 VPWR.n9 3.374
R60 VPWR.n4 VPWR.n3 2.327
R61 VPWR.n22 VPWR.n21 2.21
R62 VPWR VPWR.n24 0.484
R63 VPWR.n24 VPWR.n23 0.134
R64 VPWR.n7 VPWR.n5 0.119
R65 VPWR.n13 VPWR.n7 0.119
R66 VPWR.n15 VPWR.n13 0.119
R67 VPWR.n17 VPWR.n15 0.119
R68 VPWR.n23 VPWR.n17 0.119
R69 a_27_297.n1 a_27_297.t8 270.524
R70 a_27_297.n4 a_27_297.t0 242.137
R71 a_27_297.n4 a_27_297.n3 152.295
R72 a_27_297.n7 a_27_297.n6 150.189
R73 a_27_297.n1 a_27_297.n0 150.188
R74 a_27_297.n5 a_27_297.n2 142.402
R75 a_27_297.n6 a_27_297.n5 107.462
R76 a_27_297.n6 a_27_297.n1 91.105
R77 a_27_297.n5 a_27_297.n4 70.946
R78 a_27_297.n7 a_27_297.t4 32.505
R79 a_27_297.n0 a_27_297.t9 27.58
R80 a_27_297.n3 a_27_297.t2 26.595
R81 a_27_297.n3 a_27_297.t7 26.595
R82 a_27_297.n2 a_27_297.t5 26.595
R83 a_27_297.n2 a_27_297.t1 26.595
R84 a_27_297.n0 a_27_297.t3 26.595
R85 a_27_297.t6 a_27_297.n7 26.595
R86 VPB.t5 VPB.t6 535.669
R87 VPB.t9 VPB.t8 485.358
R88 VPB.t4 VPB.t3 449.844
R89 VPB.t6 VPB.t4 266.355
R90 VPB.t3 VPB.t9 251.557
R91 VPB.t1 VPB.t5 248.598
R92 VPB.t2 VPB.t1 248.598
R93 VPB.t7 VPB.t2 248.598
R94 VPB.t0 VPB.t7 248.598
R95 VPB VPB.t0 189.408
R96 A2.n2 A2.t2 239.74
R97 A2.n0 A2.t0 227.967
R98 A2.n2 A2.t3 149.419
R99 A2.n1 A2.t1 149.419
R100 A2.n5 A2.n0 76
R101 A2.n4 A2.n3 76
R102 A2.n3 A2.n2 56.233
R103 A2.n3 A2.n1 18.744
R104 A2.n5 A2.n4 7.912
R105 A2 A2.n5 1.396
R106 A2.n4 A2 1.396
R107 A3.n3 A3.t1 275.274
R108 A3.n0 A3.t0 234.95
R109 A3.n0 A3.t2 162.65
R110 A3.n3 A3.t3 149.419
R111 A3 A3.n0 76.581
R112 A3.n2 A3.n1 76
R113 A3.n5 A3.n4 76
R114 A3.n4 A3.n2 60.696
R115 A3.n2 A3.n0 14.281
R116 A3.n1 A3 7.33
R117 A3 A3.n5 6.167
R118 A3.n5 A3 4.538
R119 A3.n4 A3.n3 4.462
R120 A3.n1 A3 3.374
R121 B1.n0 B1.t0 221.719
R122 B1.n1 B1.t1 221.719
R123 B1.n0 B1.t2 133.353
R124 B1.n1 B1.t3 133.353
R125 B1.n3 B1.n2 76
R126 B1.n2 B1.n0 58.743
R127 B1.n3 B1 14.42
R128 B1.n4 B1.n3 10.057
R129 B1.n4 B1 6.556
R130 B1 B1.n4 6.4
R131 B1.n2 B1.n1 4.518
R132 a_730_47.n1 a_730_47.n0 237.997
R133 a_730_47.n0 a_730_47.t3 38.769
R134 a_730_47.n0 a_730_47.t2 29.538
R135 a_730_47.t1 a_730_47.n1 24.923
R136 a_730_47.n1 a_730_47.t0 24.923
R137 VGND.n0 VGND.t2 142.095
R138 VGND.n19 VGND.n18 114.711
R139 VGND.n1 VGND.t3 107.786
R140 VGND.n18 VGND.t0 24.923
R141 VGND.n18 VGND.t1 24.923
R142 VGND.n3 VGND.n2 4.65
R143 VGND.n5 VGND.n4 4.65
R144 VGND.n7 VGND.n6 4.65
R145 VGND.n9 VGND.n8 4.65
R146 VGND.n11 VGND.n10 4.65
R147 VGND.n13 VGND.n12 4.65
R148 VGND.n15 VGND.n14 4.65
R149 VGND.n17 VGND.n16 4.65
R150 VGND.n21 VGND.n20 4.65
R151 VGND.n1 VGND.n0 3.99
R152 VGND.n20 VGND.n19 0.752
R153 VGND.n3 VGND.n1 0.223
R154 VGND.n5 VGND.n3 0.119
R155 VGND.n7 VGND.n5 0.119
R156 VGND.n9 VGND.n7 0.119
R157 VGND.n11 VGND.n9 0.119
R158 VGND.n13 VGND.n11 0.119
R159 VGND.n15 VGND.n13 0.119
R160 VGND.n17 VGND.n15 0.119
R161 VGND.n21 VGND.n17 0.119
R162 VGND.n22 VGND.n21 0.119
R163 VGND VGND.n22 0.02
R164 B2.n0 B2.t0 212.079
R165 B2.n2 B2.t2 212.079
R166 B2.n0 B2.t1 139.779
R167 B2.n2 B2.t3 139.779
R168 B2.n3 B2.n2 97.909
R169 B2.n1 B2 79.047
R170 B2.n1 B2.n0 33.593
R171 B2.n2 B2.n1 27.751
R172 B2.n3 B2 17.676
R173 B2.n4 B2 11.377
R174 B2.n4 B2.n3 5.18
R175 B2 B2.n4 5.18
R176 a_27_47.n0 a_27_47.t3 247.366
R177 a_27_47.n0 a_27_47.t0 162.126
R178 a_27_47.n1 a_27_47.n0 41.979
R179 a_27_47.n1 a_27_47.t2 24.923
R180 a_27_47.t1 a_27_47.n1 24.923
C0 B1 Y 0.24fF
C1 VPWR VGND 0.13fF
C2 A3 A2 0.11fF
C3 Y A1 0.15fF
C4 VPB VPWR 0.11fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__a32oi_4.ext - technology: sky130A

.subckt sky130_fd_sc_hd__a32oi_4 A3 A2 A1 B1 Y B2 VGND VPWR VNB VPB
X0 a_27_47.t3 B1.t0 Y.t7 VNB.t6 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 a_27_297.t19 A2.t0 VPWR.t10 VPB.t19 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 a_27_47.t2 B1.t1 Y.t6 VNB.t5 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 a_27_297.t0 A3.t0 VPWR.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 VPWR.t4 A1.t0 a_27_297.t12 VPB.t12 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 a_1249_47.t3 A3.t1 VGND.t7 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 VPWR.t9 A2.t1 a_27_297.t18 VPB.t18 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 a_1249_47.t2 A3.t2 VGND.t6 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 Y.t3 B1.t2 a_27_297.t4 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 a_27_297.t13 A1.t1 VPWR.t5 VPB.t13 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 VPWR.t1 A3.t3 a_27_297.t5 VPB.t5 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 a_27_297.t14 A1.t2 VPWR.t6 VPB.t14 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 a_803_47.t7 A2.t2 a_1249_47.t4 VNB.t17 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 a_27_297.t8 B2.t0 Y.t8 VPB.t8 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14 a_27_297.t6 A3.t4 VPWR.t2 VPB.t6 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 VPWR.t7 A1.t3 a_27_297.t15 VPB.t15 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16 a_803_47.t6 A2.t3 a_1249_47.t7 VNB.t18 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X17 Y.t12 A1.t4 a_803_47.t3 VNB.t13 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X18 Y.t9 B2.t1 a_27_297.t9 VPB.t9 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X19 VPWR.t3 A3.t5 a_27_297.t7 VPB.t7 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X20 Y.t13 A1.t5 a_803_47.t2 VNB.t14 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X21 a_27_297.t10 B2.t2 Y.t10 VPB.t10 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X22 a_1249_47.t6 A2.t4 a_803_47.t5 VNB.t19 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X23 a_27_297.t17 A2.t5 VPWR.t8 VPB.t17 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X24 a_27_47.t4 B2.t3 VGND.t0 VNB.t8 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X25 a_27_47.t5 B2.t4 VGND.t1 VNB.t10 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X26 a_1249_47.t5 A2.t6 a_803_47.t4 VNB.t9 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X27 VPWR.t11 A2.t7 a_27_297.t16 VPB.t16 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X28 a_803_47.t1 A1.t6 Y.t14 VNB.t15 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X29 a_27_297.t3 B1.t3 Y.t2 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X30 a_803_47.t0 A1.t7 Y.t15 VNB.t16 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X31 VGND.t2 B2.t5 a_27_47.t6 VNB.t11 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X32 Y.t5 B1.t4 a_27_47.t1 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X33 Y.t1 B1.t5 a_27_297.t2 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X34 Y.t4 B1.t6 a_27_47.t0 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X35 a_27_297.t1 B1.t7 Y.t0 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X36 VGND.t5 A3.t6 a_1249_47.t1 VNB.t7 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X37 Y.t11 B2.t6 a_27_297.t11 VPB.t11 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X38 VGND.t4 A3.t7 a_1249_47.t0 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X39 VGND.t3 B2.t7 a_27_47.t7 VNB.t12 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
R0 B1.n0 B1.t3 212.079
R1 B1.n3 B1.t5 212.079
R2 B1.n7 B1.t7 212.079
R3 B1.n6 B1.t2 212.079
R4 B1.n0 B1.t1 139.779
R5 B1.n3 B1.t6 139.779
R6 B1.n7 B1.t0 139.779
R7 B1.n6 B1.t4 139.779
R8 B1 B1.n8 85.309
R9 B1.n2 B1.n1 76
R10 B1.n5 B1.n4 76
R11 B1.n7 B1.n6 61.345
R12 B1.n8 B1.n7 14.606
R13 B1.n5 B1.n2 13.187
R14 B1.n1 B1.n0 8.763
R15 B1 B1.n5 3.878
R16 B1.n4 B1.n3 2.921
R17 B1.n2 B1 0.775
R18 Y.n13 Y.n10 187.875
R19 Y.n9 Y.n7 187.875
R20 Y.n2 Y.n0 155.747
R21 Y.n9 Y.n8 149.475
R22 Y.n12 Y.n11 146.767
R23 Y.n4 Y.n2 102.4
R24 Y.n2 Y.n1 92.5
R25 Y.n4 Y.n3 92.5
R26 Y.n6 Y.n5 92.5
R27 Y.n6 Y.n4 63.247
R28 Y.n10 Y.t2 26.595
R29 Y.n10 Y.t1 26.595
R30 Y.n7 Y.t10 26.595
R31 Y.n7 Y.t11 26.595
R32 Y.n8 Y.t8 26.595
R33 Y.n8 Y.t9 26.595
R34 Y.n11 Y.t0 26.595
R35 Y.n11 Y.t3 26.595
R36 Y.n5 Y.t7 24.923
R37 Y.n5 Y.t5 24.923
R38 Y.n3 Y.t6 24.923
R39 Y.n3 Y.t4 24.923
R40 Y.n1 Y.t15 24.923
R41 Y.n1 Y.t13 24.923
R42 Y.n0 Y.t14 24.923
R43 Y.n0 Y.t12 24.923
R44 Y Y.n6 23.726
R45 Y.n13 Y.n9 21.835
R46 Y.n14 Y 4.266
R47 Y Y.n14 3.025
R48 Y.n14 Y.n13 1.978
R49 Y.n12 Y 1.46
R50 Y.n13 Y.n12 1.436
R51 a_27_47.n4 a_27_47.t2 238.823
R52 a_27_47.n1 a_27_47.t7 236.55
R53 a_27_47.n1 a_27_47.n0 108.688
R54 a_27_47.n3 a_27_47.n2 92.5
R55 a_27_47.n5 a_27_47.n4 92.5
R56 a_27_47.n3 a_27_47.n1 76.047
R57 a_27_47.n4 a_27_47.n3 63.247
R58 a_27_47.n0 a_27_47.t6 24.923
R59 a_27_47.n0 a_27_47.t4 24.923
R60 a_27_47.n2 a_27_47.t1 24.923
R61 a_27_47.n2 a_27_47.t5 24.923
R62 a_27_47.n5 a_27_47.t0 24.923
R63 a_27_47.t3 a_27_47.n5 24.923
R64 VNB.t18 VNB.t0 4545.05
R65 VNB.t5 VNB.t14 4545.05
R66 VNB VNB.t12 3853.91
R67 VNB.t15 VNB.t19 2707.69
R68 VNB.t1 VNB.t2 2030.77
R69 VNB.t7 VNB.t1 2030.77
R70 VNB.t0 VNB.t7 2030.77
R71 VNB.t9 VNB.t18 2030.77
R72 VNB.t17 VNB.t9 2030.77
R73 VNB.t19 VNB.t17 2030.77
R74 VNB.t13 VNB.t15 2030.77
R75 VNB.t16 VNB.t13 2030.77
R76 VNB.t14 VNB.t16 2030.77
R77 VNB.t3 VNB.t5 2030.77
R78 VNB.t6 VNB.t3 2030.77
R79 VNB.t4 VNB.t6 2030.77
R80 VNB.t10 VNB.t4 2030.77
R81 VNB.t11 VNB.t10 2030.77
R82 VNB.t8 VNB.t11 2030.77
R83 VNB.t12 VNB.t8 2030.77
R84 A2.n2 A2.t1 205.652
R85 A2.n8 A2.t5 205.652
R86 A2.n9 A2.t7 205.652
R87 A2.n1 A2.t0 205.652
R88 A2.n1 A2.t3 144.599
R89 A2.n2 A2.t6 139.779
R90 A2.n8 A2.t2 139.779
R91 A2.n9 A2.t4 139.779
R92 A2.n4 A2.n3 76
R93 A2.n7 A2.n6 76
R94 A2.n11 A2.n10 76
R95 A2.n7 A2.n0 46.822
R96 A2.n10 A2.n8 45.445
R97 A2.n3 A2.n2 38.384
R98 A2.n3 A2.n1 21.582
R99 A2.n6 A2.n5 19.342
R100 A2.n11 A2 17.635
R101 A2 A2.n4 14.222
R102 A2.n10 A2.n9 12.394
R103 A2.n4 A2 11.946
R104 A2.n2 A2.n0 9.64
R105 A2 A2.n11 8.533
R106 A2.n5 A2 5.12
R107 A2.n6 A2 1.706
R108 A2.n8 A2.n7 1.377
R109 VPWR.n15 VPWR.n14 307.239
R110 VPWR.n7 VPWR.n6 167.722
R111 VPWR.n9 VPWR.n8 164.214
R112 VPWR.n18 VPWR.n17 164.214
R113 VPWR.n1 VPWR.n0 164.214
R114 VPWR.n24 VPWR.t4 66.98
R115 VPWR.n24 VPWR.t6 65.995
R116 VPWR.n10 VPWR.n5 34.635
R117 VPWR.n19 VPWR.n3 34.635
R118 VPWR.n26 VPWR.n25 30.979
R119 VPWR.n16 VPWR.n15 28.988
R120 VPWR.n10 VPWR.n9 27.482
R121 VPWR.n6 VPWR.t0 26.595
R122 VPWR.n6 VPWR.t1 26.595
R123 VPWR.n8 VPWR.t2 26.595
R124 VPWR.n8 VPWR.t3 26.595
R125 VPWR.n14 VPWR.t10 26.595
R126 VPWR.n14 VPWR.t9 26.595
R127 VPWR.n17 VPWR.t8 26.595
R128 VPWR.n17 VPWR.t11 26.595
R129 VPWR.n0 VPWR.t5 26.595
R130 VPWR.n0 VPWR.t7 26.595
R131 VPWR.n23 VPWR.n3 25.498
R132 VPWR.n15 VPWR.n5 15.435
R133 VPWR.n26 VPWR.n1 10.917
R134 VPWR.n18 VPWR.n16 9.411
R135 VPWR.n11 VPWR.n10 4.65
R136 VPWR.n12 VPWR.n5 4.65
R137 VPWR.n15 VPWR.n13 4.65
R138 VPWR.n16 VPWR.n4 4.65
R139 VPWR.n20 VPWR.n19 4.65
R140 VPWR.n21 VPWR.n3 4.65
R141 VPWR.n23 VPWR.n22 4.65
R142 VPWR.n25 VPWR.n2 4.65
R143 VPWR.n27 VPWR.n26 4.65
R144 VPWR.n28 VPWR.n1 4.126
R145 VPWR.n25 VPWR.n24 3.955
R146 VPWR.n9 VPWR.n7 3.671
R147 VPWR.n24 VPWR.n23 2.66
R148 VPWR VPWR.n28 0.942
R149 VPWR.n19 VPWR.n18 0.376
R150 VPWR.n11 VPWR.n7 0.256
R151 VPWR.n28 VPWR.n27 0.134
R152 VPWR.n12 VPWR.n11 0.119
R153 VPWR.n13 VPWR.n12 0.119
R154 VPWR.n13 VPWR.n4 0.119
R155 VPWR.n20 VPWR.n4 0.119
R156 VPWR.n21 VPWR.n20 0.119
R157 VPWR.n22 VPWR.n21 0.119
R158 VPWR.n22 VPWR.n2 0.119
R159 VPWR.n27 VPWR.n2 0.119
R160 a_27_297.n15 a_27_297.t11 624.727
R161 a_27_297.n11 a_27_297.n10 292.5
R162 a_27_297.n13 a_27_297.n12 292.5
R163 a_27_297.n15 a_27_297.n14 292.5
R164 a_27_297.n17 a_27_297.n16 292.5
R165 a_27_297.n5 a_27_297.t0 258.413
R166 a_27_297.n5 a_27_297.n4 168.571
R167 a_27_297.n6 a_27_297.n3 168.571
R168 a_27_297.n7 a_27_297.n2 168.571
R169 a_27_297.n8 a_27_297.n1 168.571
R170 a_27_297.n9 a_27_297.n0 168.571
R171 a_27_297.n3 a_27_297.t7 129.035
R172 a_27_297.n11 a_27_297.n9 103.152
R173 a_27_297.n6 a_27_297.n5 102.4
R174 a_27_297.n9 a_27_297.n8 93.741
R175 a_27_297.n8 a_27_297.n7 80.941
R176 a_27_297.n1 a_27_297.t16 72.89
R177 a_27_297.n7 a_27_297.n6 63.247
R178 a_27_297.n13 a_27_297.n11 63.247
R179 a_27_297.n16 a_27_297.n13 63.247
R180 a_27_297.n16 a_27_297.n15 63.247
R181 a_27_297.n10 a_27_297.t15 30.535
R182 a_27_297.n14 a_27_297.t9 26.595
R183 a_27_297.n14 a_27_297.t10 26.595
R184 a_27_297.n12 a_27_297.t2 26.595
R185 a_27_297.n12 a_27_297.t1 26.595
R186 a_27_297.n4 a_27_297.t5 26.595
R187 a_27_297.n4 a_27_297.t6 26.595
R188 a_27_297.n3 a_27_297.t19 26.595
R189 a_27_297.n2 a_27_297.t18 26.595
R190 a_27_297.n2 a_27_297.t17 26.595
R191 a_27_297.n1 a_27_297.t14 26.595
R192 a_27_297.n0 a_27_297.t12 26.595
R193 a_27_297.n0 a_27_297.t13 26.595
R194 a_27_297.n10 a_27_297.t3 26.595
R195 a_27_297.t4 a_27_297.n17 26.595
R196 a_27_297.n17 a_27_297.t8 26.595
R197 VPB.t19 VPB.t7 556.386
R198 VPB.t12 VPB.t14 488.317
R199 VPB.t14 VPB.t16 387.694
R200 VPB.t3 VPB.t15 260.436
R201 VPB.t5 VPB.t0 248.598
R202 VPB.t6 VPB.t5 248.598
R203 VPB.t7 VPB.t6 248.598
R204 VPB.t18 VPB.t19 248.598
R205 VPB.t17 VPB.t18 248.598
R206 VPB.t16 VPB.t17 248.598
R207 VPB.t13 VPB.t12 248.598
R208 VPB.t15 VPB.t13 248.598
R209 VPB.t2 VPB.t3 248.598
R210 VPB.t1 VPB.t2 248.598
R211 VPB.t4 VPB.t1 248.598
R212 VPB.t8 VPB.t4 248.598
R213 VPB.t9 VPB.t8 248.598
R214 VPB.t10 VPB.t9 248.598
R215 VPB.t11 VPB.t10 248.598
R216 VPB VPB.t11 139.096
R217 A3.n1 A3.t0 212.079
R218 A3.n4 A3.t3 212.079
R219 A3.n7 A3.t4 212.079
R220 A3.n5 A3.t5 212.079
R221 A3.n1 A3.t7 139.779
R222 A3.n4 A3.t2 139.779
R223 A3.n7 A3.t6 139.779
R224 A3.n5 A3.t1 139.779
R225 A3.n1 A3.n0 106.067
R226 A3.n3 A3.n2 76
R227 A3.n12 A3.n11 76
R228 A3.n10 A3.n9 76
R229 A3.n11 A3.n10 49.66
R230 A3.n7 A3.n6 48.2
R231 A3.n0 A3 26.726
R232 A3.n2 A3.n1 21.909
R233 A3.n9 A3.n8 21.229
R234 A3.n3 A3 20.604
R235 A3.n12 A3 15.609
R236 A3.n6 A3.n5 13.145
R237 A3 A3.n12 13.112
R238 A3.n11 A3.n4 10.224
R239 A3 A3.n3 8.117
R240 A3.n9 A3 5.619
R241 A3.n8 A3 1.873
R242 A3.n10 A3.n7 1.46
R243 A3.n0 A3 0.624
R244 A1.n1 A1.t2 230.864
R245 A1.n5 A1.t3 218.046
R246 A1.n11 A1.t0 205.652
R247 A1.n6 A1.t1 205.652
R248 A1.n2 A1.t6 169.865
R249 A1.n3 A1.t5 139.779
R250 A1.n12 A1.t7 139.779
R251 A1.n0 A1.t4 139.779
R252 A1 A1.n2 80.573
R253 A1.n14 A1.n13 76
R254 A1.n10 A1.n9 76
R255 A1.n8 A1.n7 76
R256 A1.n6 A1.n5 45.445
R257 A1.n10 A1.n3 37.182
R258 A1.n13 A1.n12 26.165
R259 A1.n8 A1.n4 20.723
R260 A1.n9 A1 18.895
R261 A1 A1.n14 16.457
R262 A1.n14 A1 11.58
R263 A1.n12 A1.n11 11.017
R264 A1.n1 A1.n0 10.328
R265 A1.n11 A1.n10 9.64
R266 A1.n7 A1.n3 9.64
R267 A1.n9 A1 9.142
R268 A1.n4 A1 5.485
R269 A1.n2 A1.n1 1.915
R270 A1 A1.n8 1.828
R271 A1.n7 A1.n6 1.377
R272 VGND.n14 VGND.t7 190.315
R273 VGND.n10 VGND.t4 187.869
R274 VGND.n12 VGND.n11 107.239
R275 VGND.n36 VGND.n2 107.239
R276 VGND.n39 VGND.n38 107.239
R277 VGND.n18 VGND.n8 34.635
R278 VGND.n19 VGND.n18 34.635
R279 VGND.n20 VGND.n19 34.635
R280 VGND.n20 VGND.n6 34.635
R281 VGND.n24 VGND.n6 34.635
R282 VGND.n25 VGND.n24 34.635
R283 VGND.n26 VGND.n25 34.635
R284 VGND.n26 VGND.n4 34.635
R285 VGND.n30 VGND.n4 34.635
R286 VGND.n31 VGND.n30 34.635
R287 VGND.n32 VGND.n31 34.635
R288 VGND.n32 VGND.n1 34.635
R289 VGND.n14 VGND.n8 30.494
R290 VGND.n36 VGND.n1 28.988
R291 VGND.n11 VGND.t6 24.923
R292 VGND.n11 VGND.t5 24.923
R293 VGND.n2 VGND.t1 24.923
R294 VGND.n2 VGND.t2 24.923
R295 VGND.n38 VGND.t0 24.923
R296 VGND.n38 VGND.t3 24.923
R297 VGND.n13 VGND.n12 24.47
R298 VGND.n39 VGND.n37 22.964
R299 VGND.n37 VGND.n36 15.435
R300 VGND.n14 VGND.n13 13.929
R301 VGND.n13 VGND.n9 4.65
R302 VGND.n15 VGND.n14 4.65
R303 VGND.n16 VGND.n8 4.65
R304 VGND.n18 VGND.n17 4.65
R305 VGND.n19 VGND.n7 4.65
R306 VGND.n21 VGND.n20 4.65
R307 VGND.n22 VGND.n6 4.65
R308 VGND.n24 VGND.n23 4.65
R309 VGND.n25 VGND.n5 4.65
R310 VGND.n27 VGND.n26 4.65
R311 VGND.n28 VGND.n4 4.65
R312 VGND.n30 VGND.n29 4.65
R313 VGND.n31 VGND.n3 4.65
R314 VGND.n33 VGND.n32 4.65
R315 VGND.n34 VGND.n1 4.65
R316 VGND.n36 VGND.n35 4.65
R317 VGND.n37 VGND.n0 4.65
R318 VGND.n40 VGND.n39 3.932
R319 VGND.n12 VGND.n10 3.75
R320 VGND.n10 VGND.n9 0.265
R321 VGND.n40 VGND.n0 0.137
R322 VGND.n15 VGND.n9 0.119
R323 VGND.n16 VGND.n15 0.119
R324 VGND.n17 VGND.n16 0.119
R325 VGND.n17 VGND.n7 0.119
R326 VGND.n21 VGND.n7 0.119
R327 VGND.n22 VGND.n21 0.119
R328 VGND.n23 VGND.n22 0.119
R329 VGND.n23 VGND.n5 0.119
R330 VGND.n27 VGND.n5 0.119
R331 VGND.n28 VGND.n27 0.119
R332 VGND.n29 VGND.n28 0.119
R333 VGND.n29 VGND.n3 0.119
R334 VGND.n33 VGND.n3 0.119
R335 VGND.n34 VGND.n33 0.119
R336 VGND.n35 VGND.n34 0.119
R337 VGND.n35 VGND.n0 0.119
R338 VGND VGND.n40 0.101
R339 a_1249_47.n4 a_1249_47.n0 171.935
R340 a_1249_47.n3 a_1249_47.n2 155.747
R341 a_1249_47.n5 a_1249_47.n4 108.688
R342 a_1249_47.n4 a_1249_47.n3 102.4
R343 a_1249_47.n3 a_1249_47.n1 92.5
R344 a_1249_47.n2 a_1249_47.t4 24.923
R345 a_1249_47.n2 a_1249_47.t6 24.923
R346 a_1249_47.n1 a_1249_47.t7 24.923
R347 a_1249_47.n1 a_1249_47.t5 24.923
R348 a_1249_47.n0 a_1249_47.t0 24.923
R349 a_1249_47.n0 a_1249_47.t2 24.923
R350 a_1249_47.n5 a_1249_47.t1 24.923
R351 a_1249_47.t3 a_1249_47.n5 24.923
R352 a_803_47.n1 a_803_47.t6 238.823
R353 a_803_47.n4 a_803_47.t2 238.823
R354 a_803_47.n1 a_803_47.n0 92.5
R355 a_803_47.n3 a_803_47.n2 92.5
R356 a_803_47.n5 a_803_47.n4 92.5
R357 a_803_47.n3 a_803_47.n1 73.788
R358 a_803_47.n4 a_803_47.n3 63.247
R359 a_803_47.n2 a_803_47.t5 50.769
R360 a_803_47.n2 a_803_47.t1 24.923
R361 a_803_47.n0 a_803_47.t4 24.923
R362 a_803_47.n0 a_803_47.t7 24.923
R363 a_803_47.t3 a_803_47.n5 24.923
R364 a_803_47.n5 a_803_47.t0 24.923
R365 B2.n0 B2.t0 212.079
R366 B2.n1 B2.t1 212.079
R367 B2.n8 B2.t2 212.079
R368 B2.n6 B2.t6 212.079
R369 B2.n0 B2.t4 139.779
R370 B2.n1 B2.t5 139.779
R371 B2.n8 B2.t3 139.779
R372 B2.n6 B2.t7 139.779
R373 B2.n6 B2.n5 106.898
R374 B2.n11 B2.n2 76
R375 B2.n10 B2.n9 76
R376 B2.n1 B2.n0 61.345
R377 B2.n9 B2.n2 49.66
R378 B2.n8 B2.n7 40.166
R379 B2.n7 B2.n6 21.178
R380 B2.n10 B2.n3 18.921
R381 B2.n5 B2 18.643
R382 B2 B2.n11 13.078
R383 B2.n11 B2 12.521
R384 B2.n9 B2.n8 9.493
R385 B2.n4 B2 8.145
R386 B2 B2.n10 6.4
R387 B2.n4 B2 3.895
R388 B2.n5 B2.n4 3.06
R389 B2.n2 B2.n1 2.19
R390 B2 B2.n3 0.278
C0 VPWR VGND 0.21fF
C1 VPWR VPB 0.19fF
C2 Y B1 0.33fF
C3 Y B2 0.24fF
C4 Y A1 0.19fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__a41o_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__a41o_1 VGND VPWR A3 A4 A2 X B1 A1 VNB VPB
X0 a_465_47.t1 A2.t0 a_381_47.t1 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 VGND.t1 A4.t0 a_561_47.t1 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 VPWR.t3 A3.t0 a_297_297.t4 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 a_297_297.t3 A2.t1 VPWR.t2 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 a_297_297.t2 A4.t1 VPWR.t1 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 VPWR.t0 A1.t0 a_297_297.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 a_381_47.t0 A1.t1 a_79_21.t2 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 a_297_297.t1 B1.t0 a_79_21.t1 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 VPWR.t4 a_79_21.t3 X.t0 VPB.t5 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 a_79_21.t0 B1.t1 VGND.t0 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 VGND.t2 a_79_21.t4 X.t1 VNB.t5 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 a_561_47.t0 A3.t1 a_465_47.t0 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
R0 A2.n0 A2.t1 241.534
R1 A2.n0 A2.t0 169.234
R2 A2.n1 A2.n0 114.109
R3 A2.n1 A2 14.875
R4 A2 A2.n1 4.995
R5 a_381_47.t0 a_381_47.t1 49.846
R6 a_465_47.t0 a_465_47.t1 60.923
R7 VNB VNB.t5 6053.91
R8 VNB.t2 VNB.t0 3457.14
R9 VNB.t5 VNB.t2 3118.68
R10 VNB.t3 VNB.t1 2320.88
R11 VNB.t4 VNB.t3 2320.88
R12 VNB.t0 VNB.t4 2030.77
R13 A4.n0 A4.t1 230.154
R14 A4.n0 A4.t0 157.854
R15 A4.n1 A4.n0 76
R16 A4.n1 A4 14.305
R17 A4 A4.n1 2.76
R18 a_561_47.t0 a_561_47.t1 60.923
R19 VGND.n1 VGND.n0 114.495
R20 VGND.n1 VGND.t1 107.695
R21 VGND.n0 VGND.t0 51.692
R22 VGND.n0 VGND.t2 39.692
R23 VGND VGND.n1 0.149
R24 A3.n0 A3.t0 241.534
R25 A3.n0 A3.t1 169.234
R26 A3.n1 A3.n0 76
R27 A3 A3.n1 9.6
R28 A3.n1 A3 1.852
R29 a_297_297.n1 a_297_297.t2 251.172
R30 a_297_297.n2 a_297_297.n1 215.544
R31 a_297_297.n1 a_297_297.n0 152.295
R32 a_297_297.n0 a_297_297.t4 38.415
R33 a_297_297.n0 a_297_297.t3 26.595
R34 a_297_297.t0 a_297_297.n2 26.595
R35 a_297_297.n2 a_297_297.t1 26.595
R36 VPWR.n8 VPWR.t4 580.936
R37 VPWR.n3 VPWR.n2 315.608
R38 VPWR.n1 VPWR.n0 311.956
R39 VPWR.n2 VPWR.t1 32.505
R40 VPWR.n2 VPWR.t3 32.505
R41 VPWR.n0 VPWR.t2 26.595
R42 VPWR.n0 VPWR.t0 26.595
R43 VPWR.n5 VPWR.n4 4.65
R44 VPWR.n7 VPWR.n6 4.65
R45 VPWR.n9 VPWR.n8 4.05
R46 VPWR.n3 VPWR.n1 3.962
R47 VPWR.n5 VPWR.n3 0.211
R48 VPWR.n9 VPWR.n7 0.134
R49 VPWR VPWR.n9 0.124
R50 VPWR.n7 VPWR.n5 0.119
R51 VPB.t5 VPB.t1 556.386
R52 VPB.t4 VPB.t2 284.112
R53 VPB.t3 VPB.t4 284.112
R54 VPB.t0 VPB.t3 248.598
R55 VPB.t1 VPB.t0 248.598
R56 VPB VPB.t5 189.408
R57 A1.n0 A1.t0 241.534
R58 A1.n0 A1.t1 169.234
R59 A1 A1.n0 87.414
R60 a_79_21.t1 a_79_21.n2 262.383
R61 a_79_21.n0 a_79_21.t3 235.47
R62 a_79_21.n0 a_79_21.t4 163.17
R63 a_79_21.n2 a_79_21.n1 125.224
R64 a_79_21.n2 a_79_21.n0 76
R65 a_79_21.n1 a_79_21.t2 72
R66 a_79_21.n1 a_79_21.t0 32.307
R67 B1.n0 B1.t0 229.752
R68 B1.n0 B1.t1 157.452
R69 B1.n1 B1.n0 76
R70 B1.n1 B1 11.054
R71 B1 B1.n1 2.133
R72 X.n2 X.n1 299.088
R73 X.n5 X.n2 292.5
R74 X.t1 X 174.774
R75 X.n4 X.t1 168.653
R76 X.n2 X.t0 26.595
R77 X X.n0 10.584
R78 X.n5 X 10.584
R79 X.n4 X.n3 8.123
R80 X.n3 X 6.646
R81 X X.n0 6.153
R82 X X.n5 6.153
R83 X X.n3 5.082
R84 X.n1 X 1.969
R85 X X.n4 1.969
R86 X.n1 X 1.505
C0 A2 A1 0.11fF
C1 A2 A3 0.14fF
C2 A3 A4 0.13fF
C3 B1 A1 0.13fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__a41o_2.ext - technology: sky130A

.subckt sky130_fd_sc_hd__a41o_2 B1 A1 X A2 A4 A3 VGND VPWR VNB VPB
X0 a_381_297.t0 A1.t0 VPWR.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 VPWR.t4 A2.t0 a_381_297.t3 VPB.t5 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 a_465_47.t0 A4.t0 VGND.t1 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 a_549_47.t1 A3.t0 a_465_47.t1 VNB.t6 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 VPWR.t2 a_79_21.t3 X.t3 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 VGND.t2 a_79_21.t4 X.t1 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 a_665_47.t1 A2.t1 a_549_47.t0 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 a_381_297.t4 A3.t1 VPWR.t5 VPB.t6 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 VPWR.t1 A4.t1 a_381_297.t2 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 a_381_297.t1 B1.t0 a_79_21.t1 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 a_79_21.t0 A1.t1 a_665_47.t0 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 VGND.t0 B1.t1 a_79_21.t2 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 X.t2 a_79_21.t5 VPWR.t3 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13 X.t0 a_79_21.t6 VGND.t3 VNB.t5 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
R0 A1.n0 A1.t0 231.476
R1 A1.n0 A1.t1 159.176
R2 A1.n1 A1.n0 76
R3 A1.n1 A1 16.581
R4 A1 A1.n1 3.2
R5 VPWR.n3 VPWR.n0 315.627
R6 VPWR.n2 VPWR.n1 311.956
R7 VPWR.n8 VPWR.t2 196.528
R8 VPWR.n12 VPWR.t3 145.867
R9 VPWR.n1 VPWR.t5 26.595
R10 VPWR.n1 VPWR.t1 26.595
R11 VPWR.n0 VPWR.t0 26.595
R12 VPWR.n0 VPWR.t4 26.595
R13 VPWR.n5 VPWR.n4 4.65
R14 VPWR.n7 VPWR.n6 4.65
R15 VPWR.n9 VPWR.n8 4.65
R16 VPWR.n11 VPWR.n10 4.65
R17 VPWR.n13 VPWR.n12 4.65
R18 VPWR.n3 VPWR.n2 4.021
R19 VPWR.n5 VPWR.n3 0.199
R20 VPWR.n7 VPWR.n5 0.119
R21 VPWR.n9 VPWR.n7 0.119
R22 VPWR.n11 VPWR.n9 0.119
R23 VPWR.n13 VPWR.n11 0.119
R24 VPWR VPWR.n13 0.02
R25 a_381_297.t0 a_381_297.n2 254.186
R26 a_381_297.n2 a_381_297.n1 215.542
R27 a_381_297.n2 a_381_297.n0 152.295
R28 a_381_297.n0 a_381_297.t3 58.115
R29 a_381_297.n1 a_381_297.t2 26.595
R30 a_381_297.n1 a_381_297.t1 26.595
R31 a_381_297.n0 a_381_297.t4 26.595
R32 VPB.t3 VPB.t1 556.386
R33 VPB.t6 VPB.t5 343.302
R34 VPB.t5 VPB.t0 248.598
R35 VPB.t2 VPB.t6 248.598
R36 VPB.t1 VPB.t2 248.598
R37 VPB.t4 VPB.t3 248.598
R38 VPB VPB.t4 189.408
R39 A2.n0 A2.t0 241.534
R40 A2.n0 A2.t1 169.234
R41 A2.n1 A2.n0 82.4
R42 A2.n1 A2 16.967
R43 A2 A2.n1 3.274
R44 A4.n0 A4.t1 241.534
R45 A4.n0 A4.t0 169.234
R46 A4.n1 A4.n0 76
R47 A4.n1 A4 10.889
R48 A4 A4.n1 2.101
R49 VGND.n1 VGND.t2 190.315
R50 VGND.n2 VGND.n0 110.767
R51 VGND.n5 VGND.t3 103.506
R52 VGND.n0 VGND.t1 24.923
R53 VGND.n0 VGND.t0 24.923
R54 VGND.n6 VGND.n5 4.65
R55 VGND.n4 VGND.n3 4.65
R56 VGND.n2 VGND.n1 3.921
R57 VGND.n4 VGND.n2 0.225
R58 VGND.n6 VGND.n4 0.119
R59 VGND VGND.n6 0.02
R60 a_465_47.t0 a_465_47.t1 49.846
R61 VNB VNB.t5 6053.91
R62 VNB.t4 VNB.t2 4545.05
R63 VNB.t6 VNB.t1 2804.4
R64 VNB.t1 VNB.t0 2030.77
R65 VNB.t3 VNB.t6 2030.77
R66 VNB.t2 VNB.t3 2030.77
R67 VNB.t5 VNB.t4 2030.77
R68 A3.n0 A3.t1 237.733
R69 A3.n0 A3.t0 165.433
R70 A3 A3.n0 105.799
R71 a_549_47.t0 a_549_47.t1 79.384
R72 a_79_21.n2 a_79_21.t0 352.14
R73 a_79_21.t1 a_79_21.n3 246.948
R74 a_79_21.n1 a_79_21.t3 212.079
R75 a_79_21.n0 a_79_21.t5 212.079
R76 a_79_21.n2 a_79_21.t2 175.4
R77 a_79_21.n1 a_79_21.t4 139.779
R78 a_79_21.n0 a_79_21.t6 139.779
R79 a_79_21.n3 a_79_21.n1 101.56
R80 a_79_21.n1 a_79_21.n0 61.345
R81 a_79_21.n3 a_79_21.n2 59.105
R82 X.n1 X.n0 146.413
R83 X X.n2 115.384
R84 X.n0 X.t3 26.595
R85 X.n0 X.t2 26.595
R86 X.n2 X.t1 24.923
R87 X.n2 X.t0 24.923
R88 X X.n1 17.138
R89 X.n1 X 5.564
R90 a_665_47.t0 a_665_47.t1 49.846
R91 B1.n0 B1.t0 228.822
R92 B1.n0 B1.t1 156.522
R93 B1 B1.n0 78.133
C0 A2 A1 0.17fF
C1 A2 A3 0.11fF
C2 VGND X 0.12fF
C3 VGND VPWR 0.11fF
C4 VPWR X 0.20fF
C5 A4 A3 0.11fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__a41o_4.ext - technology: sky130A

.subckt sky130_fd_sc_hd__a41o_4 X A4 A3 A2 A1 B1 VGND VPWR VNB VPB
X0 a_639_47.t3 A1.t0 a_79_21.t5 VNB.t9 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 a_639_47.t0 A2.t0 a_889_47.t1 VNB.t5 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 VPWR.t11 a_79_21.t6 X.t7 VPB.t13 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 VPWR.t4 A3.t0 a_467_297.t3 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 a_889_47.t0 A2.t1 a_639_47.t1 VNB.t6 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 a_889_47.t2 A3.t1 a_1079_47.t1 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 X.t6 a_79_21.t7 VPWR.t10 VPB.t12 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 VGND.t3 B1.t0 a_79_21.t1 VNB.t7 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 VPWR.t9 a_79_21.t8 X.t5 VPB.t11 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 a_467_297.t4 A4.t0 VPWR.t2 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 VGND.t7 a_79_21.t9 X.t4 VNB.t13 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 VGND.t6 a_79_21.t10 X.t3 VNB.t12 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 a_467_297.t6 B1.t1 a_79_21.t2 VPB.t6 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13 a_467_297.t1 A2.t2 VPWR.t1 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14 VPWR.t3 A4.t1 a_467_297.t5 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 a_1079_47.t0 A3.t2 a_889_47.t3 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X16 a_79_21.t3 B1.t2 a_467_297.t7 VPB.t7 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17 a_79_21.t0 B1.t3 VGND.t2 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X18 a_1079_47.t2 A4.t2 VGND.t0 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X19 VPWR.t0 A2.t3 a_467_297.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X20 X.t2 a_79_21.t11 VGND.t5 VNB.t11 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X21 a_467_297.t9 A1.t1 VPWR.t7 VPB.t9 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X22 a_79_21.t4 A1.t2 a_639_47.t2 VNB.t8 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X23 VPWR.t6 A1.t3 a_467_297.t8 VPB.t8 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X24 a_467_297.t2 A3.t3 VPWR.t5 VPB.t5 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X25 VGND.t1 A4.t3 a_1079_47.t3 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X26 X.t0 a_79_21.t12 VPWR.t8 VPB.t10 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X27 X.t1 a_79_21.t13 VGND.t4 VNB.t10 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
R0 A1.n0 A1.t1 212.079
R1 A1.n2 A1.t3 212.079
R2 A1.n0 A1.t0 139.779
R3 A1.n2 A1.t2 139.779
R4 A1 A1.n1 77.745
R5 A1.n4 A1.n3 76
R6 A1 A1.n4 18.036
R7 A1.n4 A1 8.727
R8 A1.n1 A1.n0 7.303
R9 A1.n3 A1.n2 4.381
R10 a_79_21.n15 a_79_21.n14 249.926
R11 a_79_21.n11 a_79_21.t6 212.079
R12 a_79_21.n3 a_79_21.t7 212.079
R13 a_79_21.n7 a_79_21.t8 212.079
R14 a_79_21.n5 a_79_21.t12 212.079
R15 a_79_21.n2 a_79_21.n1 194.9
R16 a_79_21.n11 a_79_21.t10 139.779
R17 a_79_21.n3 a_79_21.t11 139.779
R18 a_79_21.n7 a_79_21.t9 139.779
R19 a_79_21.n5 a_79_21.t13 139.779
R20 a_79_21.n2 a_79_21.n0 109.441
R21 a_79_21.n9 a_79_21.n6 101.6
R22 a_79_21.n10 a_79_21.n4 76
R23 a_79_21.n9 a_79_21.n8 76
R24 a_79_21.n13 a_79_21.n12 76
R25 a_79_21.n14 a_79_21.n2 58.728
R26 a_79_21.n6 a_79_21.n5 27.021
R27 a_79_21.t2 a_79_21.n15 26.595
R28 a_79_21.n15 a_79_21.t3 26.595
R29 a_79_21.n13 a_79_21.n10 25.6
R30 a_79_21.n10 a_79_21.n9 25.6
R31 a_79_21.n1 a_79_21.t5 24.923
R32 a_79_21.n1 a_79_21.t4 24.923
R33 a_79_21.n0 a_79_21.t1 24.923
R34 a_79_21.n0 a_79_21.t0 24.923
R35 a_79_21.n8 a_79_21.n7 15.336
R36 a_79_21.n14 a_79_21.n13 13.929
R37 a_79_21.n12 a_79_21.n11 8.033
R38 a_79_21.n4 a_79_21.n3 3.651
R39 a_639_47.t2 a_639_47.n1 252.375
R40 a_639_47.n1 a_639_47.t0 234.208
R41 a_639_47.n1 a_639_47.n0 92.5
R42 a_639_47.n0 a_639_47.t1 24.923
R43 a_639_47.n0 a_639_47.t3 24.923
R44 VNB VNB.t10 6053.91
R45 VNB.t5 VNB.t3 4545.05
R46 VNB.t7 VNB.t8 4545.05
R47 VNB.t12 VNB.t0 2127.47
R48 VNB.t2 VNB.t1 2030.77
R49 VNB.t4 VNB.t2 2030.77
R50 VNB.t3 VNB.t4 2030.77
R51 VNB.t6 VNB.t5 2030.77
R52 VNB.t9 VNB.t6 2030.77
R53 VNB.t8 VNB.t9 2030.77
R54 VNB.t0 VNB.t7 2030.77
R55 VNB.t11 VNB.t12 2030.77
R56 VNB.t13 VNB.t11 2030.77
R57 VNB.t10 VNB.t13 2030.77
R58 A2.n0 A2.t2 221.719
R59 A2.n2 A2.t3 221.719
R60 A2.n0 A2.t0 149.419
R61 A2.n2 A2.t1 149.419
R62 A2.n5 A2.n1 76
R63 A2.n4 A2.n3 76
R64 A2.n5 A2.n4 20.723
R65 A2.n3 A2.n2 12.496
R66 A2.n4 A2 6.704
R67 A2.n1 A2.n0 1.785
R68 A2 A2.n5 0.609
R69 a_889_47.n1 a_889_47.n0 287.4
R70 a_889_47.n0 a_889_47.t3 24.923
R71 a_889_47.n0 a_889_47.t2 24.923
R72 a_889_47.t1 a_889_47.n1 24.923
R73 a_889_47.n1 a_889_47.t0 24.923
R74 X.n5 X.n4 231.818
R75 X.n2 X.n1 171.935
R76 X.n5 X.n3 168.571
R77 X.n2 X.n0 108.688
R78 X.n6 X.n5 33.505
R79 X.n7 X.n2 33.505
R80 X.n4 X.t7 26.595
R81 X.n4 X.t6 26.595
R82 X.n3 X.t5 26.595
R83 X.n3 X.t0 26.595
R84 X.n0 X.t4 24.923
R85 X.n0 X.t1 24.923
R86 X.n1 X.t3 24.923
R87 X.n1 X.t2 24.923
R88 X.n7 X 22.588
R89 X X.n6 9.788
R90 X.n6 X 6.4
R91 X.n7 X 6.4
R92 X X.n7 3.011
R93 VPWR.n31 VPWR.t8 190.809
R94 VPWR.n22 VPWR.t11 189.787
R95 VPWR.n3 VPWR.n0 167.647
R96 VPWR.n27 VPWR.n26 164.214
R97 VPWR.n13 VPWR.n12 164.214
R98 VPWR.n9 VPWR.n8 164.214
R99 VPWR.n1 VPWR.t5 68.927
R100 VPWR.n1 VPWR.t4 68.926
R101 VPWR.n2 VPWR.n1 67.448
R102 VPWR.n26 VPWR.t10 26.595
R103 VPWR.n26 VPWR.t9 26.595
R104 VPWR.n12 VPWR.t7 26.595
R105 VPWR.n12 VPWR.t6 26.595
R106 VPWR.n8 VPWR.t1 26.595
R107 VPWR.n8 VPWR.t0 26.595
R108 VPWR.n0 VPWR.t2 26.595
R109 VPWR.n0 VPWR.t3 26.595
R110 VPWR.n5 VPWR.n4 4.65
R111 VPWR.n7 VPWR.n6 4.65
R112 VPWR.n11 VPWR.n10 4.65
R113 VPWR.n15 VPWR.n14 4.65
R114 VPWR.n17 VPWR.n16 4.65
R115 VPWR.n19 VPWR.n18 4.65
R116 VPWR.n21 VPWR.n20 4.65
R117 VPWR.n23 VPWR.n22 4.65
R118 VPWR.n25 VPWR.n24 4.65
R119 VPWR.n28 VPWR.n27 4.65
R120 VPWR.n30 VPWR.n29 4.65
R121 VPWR.n32 VPWR.n31 4.65
R122 VPWR.n3 VPWR.n2 3.548
R123 VPWR.n10 VPWR.n9 3.388
R124 VPWR.n14 VPWR.n13 0.376
R125 VPWR.n5 VPWR.n3 0.241
R126 VPWR.n7 VPWR.n5 0.119
R127 VPWR.n11 VPWR.n7 0.119
R128 VPWR.n15 VPWR.n11 0.119
R129 VPWR.n17 VPWR.n15 0.119
R130 VPWR.n19 VPWR.n17 0.119
R131 VPWR.n21 VPWR.n19 0.119
R132 VPWR.n23 VPWR.n21 0.119
R133 VPWR.n25 VPWR.n23 0.119
R134 VPWR.n28 VPWR.n25 0.119
R135 VPWR.n30 VPWR.n28 0.119
R136 VPWR.n32 VPWR.n30 0.119
R137 VPWR VPWR.n32 0.02
R138 VPB.t13 VPB.t7 556.386
R139 VPB.t4 VPB.t5 544.548
R140 VPB.t1 VPB.t4 260.436
R141 VPB.t6 VPB.t8 260.436
R142 VPB.t3 VPB.t2 248.598
R143 VPB.t5 VPB.t3 248.598
R144 VPB.t0 VPB.t1 248.598
R145 VPB.t9 VPB.t0 248.598
R146 VPB.t8 VPB.t9 248.598
R147 VPB.t7 VPB.t6 248.598
R148 VPB.t12 VPB.t13 248.598
R149 VPB.t11 VPB.t12 248.598
R150 VPB.t10 VPB.t11 248.598
R151 VPB VPB.t10 189.408
R152 A3.n5 A3.t0 237.785
R153 A3.n0 A3.t3 221.719
R154 A3.n0 A3.t2 149.419
R155 A3.n2 A3.t1 149.419
R156 A3.n1 A3 92.872
R157 A3.n4 A3.n3 76
R158 A3.n6 A3.n5 76
R159 A3.n2 A3.n1 51.77
R160 A3.n1 A3.n0 23.207
R161 A3.n6 A3.n4 20.945
R162 A3.n3 A3.n2 8.925
R163 A3 A3.n6 4.072
R164 A3.n4 A3 2.909
R165 a_467_297.n1 a_467_297.t4 261.425
R166 a_467_297.n4 a_467_297.t7 255.733
R167 a_467_297.n1 a_467_297.n0 171.583
R168 a_467_297.n5 a_467_297.n2 171.583
R169 a_467_297.n7 a_467_297.n6 171.582
R170 a_467_297.n4 a_467_297.n3 140.205
R171 a_467_297.n6 a_467_297.n1 100.894
R172 a_467_297.n5 a_467_297.n4 94.538
R173 a_467_297.n6 a_467_297.n5 64.752
R174 a_467_297.n3 a_467_297.t6 30.535
R175 a_467_297.t1 a_467_297.n7 30.535
R176 a_467_297.n0 a_467_297.t5 26.595
R177 a_467_297.n0 a_467_297.t2 26.595
R178 a_467_297.n2 a_467_297.t0 26.595
R179 a_467_297.n2 a_467_297.t9 26.595
R180 a_467_297.n3 a_467_297.t8 26.595
R181 a_467_297.n7 a_467_297.t3 26.595
R182 a_1079_47.n1 a_1079_47.t2 237.303
R183 a_1079_47.t1 a_1079_47.n1 234.208
R184 a_1079_47.n1 a_1079_47.n0 92.5
R185 a_1079_47.n0 a_1079_47.t3 24.923
R186 a_1079_47.n0 a_1079_47.t0 24.923
R187 B1.n0 B1.t1 228.145
R188 B1.n1 B1.t2 212.079
R189 B1.n2 B1.t3 158.766
R190 B1.n3 B1.t0 139.779
R191 B1.n2 B1 86.614
R192 B1 B1.n0 79.121
R193 B1.n5 B1.n4 76
R194 B1.n3 B1.n2 42.357
R195 B1 B1.n5 18.107
R196 B1.n5 B1 10.614
R197 B1.n4 B1.n3 7.303
R198 B1.n4 B1.n1 4.381
R199 VGND.n1 VGND.t3 190.315
R200 VGND.n15 VGND.t4 190.315
R201 VGND.n2 VGND.n0 111.504
R202 VGND.n11 VGND.n10 107.239
R203 VGND.n6 VGND.n5 106.397
R204 VGND.n5 VGND.t2 28.615
R205 VGND.n0 VGND.t0 24.923
R206 VGND.n0 VGND.t1 24.923
R207 VGND.n5 VGND.t6 24.923
R208 VGND.n10 VGND.t5 24.923
R209 VGND.n10 VGND.t7 24.923
R210 VGND.n2 VGND.n1 6.022
R211 VGND.n16 VGND.n15 4.65
R212 VGND.n4 VGND.n3 4.65
R213 VGND.n7 VGND.n6 4.65
R214 VGND.n9 VGND.n8 4.65
R215 VGND.n12 VGND.n11 4.65
R216 VGND.n14 VGND.n13 4.65
R217 VGND.n4 VGND.n2 0.134
R218 VGND.n7 VGND.n4 0.119
R219 VGND.n9 VGND.n7 0.119
R220 VGND.n12 VGND.n9 0.119
R221 VGND.n14 VGND.n12 0.119
R222 VGND.n16 VGND.n14 0.119
R223 VGND VGND.n16 0.02
R224 A4.n0 A4.t0 221.719
R225 A4.n1 A4.t1 221.719
R226 A4.n0 A4.t2 149.419
R227 A4.n1 A4.t3 149.419
R228 A4.n3 A4.n2 76
R229 A4.n4 A4.n0 50.848
R230 A4.n4 A4.n3 21.874
R231 A4.n2 A4.n1 16.066
R232 A4 A4.n4 4.132
R233 A4.n3 A4 0.581
C0 VPWR X 0.50fF
C1 VPB VPWR 0.16fF
C2 VGND X 0.32fF
C3 VGND VPWR 0.18fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__a41oi_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__a41oi_1 VGND VPWR A4 Y B1 A1 A2 A3 VNB VPB
X0 a_236_47.t1 A4.t0 VGND.t0 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 a_428_47.t0 A2.t0 a_336_47.t1 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 a_109_297.t2 A1.t0 VPWR.t1 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 Y.t2 A1.t1 a_428_47.t1 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 a_336_47.t0 A3.t0 a_236_47.t0 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 VPWR.t0 A4.t1 a_109_297.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 a_109_297.t1 B1.t0 Y.t0 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 a_109_297.t4 A3.t1 VPWR.t3 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 VPWR.t2 A2.t1 a_109_297.t3 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 VGND.t1 B1.t1 Y.t1 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
R0 A4.n0 A4.t1 241.534
R1 A4.n0 A4.t0 169.234
R2 A4.n1 A4.n0 76
R3 A4.n1 A4 12.579
R4 A4 A4.n1 2.427
R5 VGND VGND.n0 97.647
R6 VGND.n0 VGND.t0 45.23
R7 VGND.n0 VGND.t1 44.307
R8 a_236_47.t0 a_236_47.t1 64.615
R9 VNB.n1 VNB.n0 40700
R10 VNB VNB.n1 9350
R11 VNB.n1 VNB 3882.35
R12 VNB.t3 VNB.t4 2780.22
R13 VNB.t1 VNB.t0 2417.58
R14 VNB.n0 VNB.t1 2417.58
R15 VNB.t0 VNB.t3 2224.18
R16 VNB.n0 VNB.t2 652.747
R17 A2.n0 A2.t1 241.534
R18 A2.n0 A2.t0 169.234
R19 A2.n1 A2.n0 76
R20 A2.n1 A2 11.4
R21 A2 A2.n1 2.2
R22 a_336_47.t0 a_336_47.t1 57.23
R23 a_428_47.t0 a_428_47.t1 78.461
R24 A1.n0 A1.t0 230.361
R25 A1.n0 A1.t1 158.061
R26 A1.n1 A1.n0 76
R27 A1.n1 A1 11.96
R28 A1 A1.n1 2.308
R29 VPWR.n2 VPWR.n1 313.088
R30 VPWR.n2 VPWR.n0 312.8
R31 VPWR.n0 VPWR.t3 48.265
R32 VPWR.n1 VPWR.t2 47.28
R33 VPWR.n1 VPWR.t1 36.445
R34 VPWR.n0 VPWR.t0 32.505
R35 VPWR VPWR.n2 0.296
R36 a_109_297.n1 a_109_297.t2 246.703
R37 a_109_297.n2 a_109_297.n1 226.132
R38 a_109_297.n1 a_109_297.n0 151.425
R39 a_109_297.n2 a_109_297.t1 42.355
R40 a_109_297.t0 a_109_297.n2 41.37
R41 a_109_297.n0 a_109_297.t4 32.505
R42 a_109_297.n0 a_109_297.t3 28.565
R43 VPB.t3 VPB.t2 340.342
R44 VPB.t1 VPB.t0 340.342
R45 VPB.t0 VPB.t4 331.464
R46 VPB.t4 VPB.t3 272.274
R47 VPB VPB.t1 189.408
R48 Y.n3 Y.n2 292.5
R49 Y.n1 Y.t2 263.43
R50 Y.n4 Y.n3 147.091
R51 Y.n0 Y.t1 117.423
R52 Y.n2 Y.n1 45.511
R53 Y.n3 Y.t0 26.595
R54 Y.n1 Y.n0 12.311
R55 Y.n5 Y.n4 8.259
R56 Y.n2 Y 5.925
R57 Y.n5 Y 2.844
R58 Y.n4 Y 2.402
R59 Y Y.n5 2.292
R60 Y.n0 Y 1.254
R61 A3.n0 A3.t1 241.534
R62 A3.n0 A3.t0 169.234
R63 A3.n1 A3.n0 76
R64 A3.n1 A3 15.2
R65 A3 A3.n1 2.933
R66 B1.n0 B1.t0 233.868
R67 B1.n0 B1.t1 161.568
R68 B1.n1 B1.n0 76
R69  B1.n1 15.2
R70 B1.n1 B1 2.933
C0 B1 A4 0.16fF
C1 VGND Y 0.45fF
C2 A3 A4 0.14fF
C3 A3 A2 0.19fF
C4 Y B1 0.17fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__a41oi_2.ext - technology: sky130A

.subckt sky130_fd_sc_hd__a41oi_2 A4 A3 A2 B1 A1 Y VPWR VGND VNB VPB
X0 a_149_297.t6 B1.t0 Y.t1 VPB.t6 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_757_47.t2 A4.t0 VGND.t3 VNB.t5 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 a_757_47.t0 A3.t0 a_567_47.t3 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 VPWR.t7 A3.t1 a_149_297.t7 VPB.t7 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 Y.t0 B1.t1 a_149_297.t5 VPB.t5 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 Y.t3 B1.t2 VGND.t1 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 a_567_47.t2 A3.t2 a_757_47.t3 VNB.t7 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 VGND.t2 A4.t1 a_757_47.t1 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 VPWR.t5 A4.t2 a_149_297.t9 VPB.t9 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 a_149_297.t2 A4.t3 VPWR.t4 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 a_317_47.t2 A1.t0 Y.t4 VNB.t8 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 a_317_47.t3 A2.t0 a_567_47.t1 VNB.t6 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 a_149_297.t8 A3.t3 VPWR.t6 VPB.t8 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13 a_149_297.t3 A2.t1 VPWR.t2 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14 Y.t5 A1.t1 a_317_47.t1 VNB.t9 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X15 VPWR.t3 A2.t2 a_149_297.t4 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16 a_567_47.t0 A2.t3 a_317_47.t0 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X17 a_149_297.t0 A1.t2 VPWR.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X18 VGND.t0 B1.t3 Y.t2 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X19 VPWR.t1 A1.t3 a_149_297.t1 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
R0 B1.n0 B1.t0 228.145
R1 B1.n3 B1.t1 212.079
R2 B1.n1 B1.t2 161.688
R3 B1.n4 B1.t3 139.779
R4 B1 B1.n0 96.292
R5 B1.n6 B1.n5 76
R6 B1.n2 B1.n1 76
R7 B1.n6 B1.n2 21.229
R8 B1.n5 B1.n4 10.224
R9 B1.n2 B1 6.556
R10 B1.n5 B1.n3 4.381
R11 B1 B1.n6 0.936
R12 Y.n4 Y.n3 223.069
R13 Y.n2 Y.n1 194.9
R14 Y.n2 Y.n0 109.441
R15 Y.n5 Y.n2 40.658
R16 Y.n3 Y.t1 26.595
R17 Y.n3 Y.t0 26.595
R18 Y.n1 Y.t4 24.923
R19 Y.n1 Y.t5 24.923
R20 Y.n0 Y.t2 24.923
R21 Y.n0 Y.t3 24.923
R22 Y.n5 Y 21.835
R23 Y.n4 Y 6.4
R24 Y.n5 Y 6.4
R25 Y Y.n5 3.764
R26 Y Y.n4 0.752
R27 a_149_297.n3 a_149_297.t2 261.425
R28 a_149_297.n6 a_149_297.t5 254.228
R29 a_149_297.n3 a_149_297.n2 171.583
R30 a_149_297.n4 a_149_297.n1 171.583
R31 a_149_297.n5 a_149_297.n0 171.583
R32 a_149_297.n7 a_149_297.n6 140.206
R33 a_149_297.n4 a_149_297.n3 100.894
R34 a_149_297.n6 a_149_297.n5 94.538
R35 a_149_297.n5 a_149_297.n4 64.752
R36 a_149_297.n1 a_149_297.t3 30.535
R37 a_149_297.n2 a_149_297.t9 26.595
R38 a_149_297.n2 a_149_297.t8 26.595
R39 a_149_297.n1 a_149_297.t7 26.595
R40 a_149_297.n0 a_149_297.t4 26.595
R41 a_149_297.n0 a_149_297.t0 26.595
R42 a_149_297.n7 a_149_297.t1 26.595
R43 a_149_297.t6 a_149_297.n7 26.595
R44 VPB VPB.t5 553.426
R45 VPB.t7 VPB.t8 544.548
R46 VPB.t3 VPB.t7 260.436
R47 VPB.t9 VPB.t2 248.598
R48 VPB.t8 VPB.t9 248.598
R49 VPB.t4 VPB.t3 248.598
R50 VPB.t0 VPB.t4 248.598
R51 VPB.t1 VPB.t0 248.598
R52 VPB.t6 VPB.t1 248.598
R53 VPB.t5 VPB.t6 248.598
R54 A4.n3 A4.t2 221.719
R55 A4.n0 A4.t3 218.506
R56 A4.n3 A4.t1 149.419
R57 A4.n0 A4.t0 146.206
R58 A4.n0 A4 133.466
R59 A4.n2 A4.n1 76
R60 A4.n5 A4.n4 76
R61 A4.n2 A4 17.163
R62 A4.n5 A4 15.418
R63 A4.n4 A4.n3 12.496
R64 A4 A4.n5 10.181
R65 A4 A4.n2 9.6
R66 A4.n1 A4.n0 1.662
R67 VGND.n5 VGND.t1 190.315
R68 VGND.n1 VGND.t0 189.473
R69 VGND.n2 VGND.n0 111.573
R70 VGND.n0 VGND.t3 24.923
R71 VGND.n0 VGND.t2 24.923
R72 VGND.n6 VGND.n5 4.65
R73 VGND.n4 VGND.n3 4.65
R74 VGND.n2 VGND.n1 3.815
R75 VGND.n4 VGND.n2 0.143
R76 VGND.n6 VGND.n4 0.119
R77 VGND VGND.n6 0.022
R78 a_757_47.t2 a_757_47.n1 237.303
R79 a_757_47.n1 a_757_47.t3 234.208
R80 a_757_47.n1 a_757_47.n0 92.5
R81 a_757_47.n0 a_757_47.t1 24.923
R82 a_757_47.n0 a_757_47.t0 24.923
R83 VNB VNB.t3 6513.25
R84 VNB.t6 VNB.t7 4545.05
R85 VNB.t2 VNB.t9 4545.05
R86 VNB.t4 VNB.t5 2030.77
R87 VNB.t0 VNB.t4 2030.77
R88 VNB.t7 VNB.t0 2030.77
R89 VNB.t1 VNB.t6 2030.77
R90 VNB.t8 VNB.t1 2030.77
R91 VNB.t9 VNB.t8 2030.77
R92 VNB.t3 VNB.t2 2030.77
R93 A3.n3 A3.t1 237.785
R94 A3.n0 A3.t3 221.719
R95 A3.n0 A3.t0 149.419
R96 A3.n2 A3.t2 149.419
R97 A3.n3 A3 83.854
R98 A3 A3.n1 82.109
R99 A3.n5 A3.n4 76
R100 A3.n4 A3.n3 64.266
R101 A3.n1 A3.n0 23.207
R102 A3 A3.n5 13.672
R103 A3.n5 A3 13.09
R104 A3.n4 A3.n2 8.925
R105 a_567_47.n1 a_567_47.n0 287.4
R106 a_567_47.n0 a_567_47.t1 24.923
R107 a_567_47.n0 a_567_47.t0 24.923
R108 a_567_47.n1 a_567_47.t3 24.923
R109 a_567_47.t2 a_567_47.n1 24.923
R110 VPWR.n1 VPWR.n0 167.615
R111 VPWR.n8 VPWR.n7 164.214
R112 VPWR.n13 VPWR.n12 164.214
R113 VPWR.n2 VPWR.t7 77.815
R114 VPWR.n2 VPWR.t6 73.875
R115 VPWR.n0 VPWR.t4 26.595
R116 VPWR.n0 VPWR.t5 26.595
R117 VPWR.n7 VPWR.t2 26.595
R118 VPWR.n7 VPWR.t3 26.595
R119 VPWR.n12 VPWR.t0 26.595
R120 VPWR.n12 VPWR.t1 26.595
R121 VPWR.n4 VPWR.n3 4.65
R122 VPWR.n6 VPWR.n5 4.65
R123 VPWR.n9 VPWR.n8 4.65
R124 VPWR.n11 VPWR.n10 4.65
R125 VPWR.n14 VPWR.n13 4.027
R126 VPWR.n3 VPWR.n2 2.588
R127 VPWR VPWR.n14 0.482
R128 VPWR.n4 VPWR.n1 0.238
R129 VPWR.n14 VPWR.n11 0.137
R130 VPWR.n6 VPWR.n4 0.119
R131 VPWR.n9 VPWR.n6 0.119
R132 VPWR.n11 VPWR.n9 0.119
R133 A1.n0 A1.t2 212.079
R134 A1.n1 A1.t3 212.079
R135 A1.n0 A1.t0 139.779
R136 A1.n1 A1.t1 139.779
R137 A1 A1.n2 33.036
R138 A1.n2 A1.n0 28.327
R139 A1.n2 A1.n1 21.882
R140 a_317_47.n0 a_317_47.t1 252.375
R141 a_317_47.n0 a_317_47.t3 234.208
R142 a_317_47.n1 a_317_47.n0 92.5
R143 a_317_47.n1 a_317_47.t0 24.923
R144 a_317_47.t2 a_317_47.n1 24.923
R145 A2.n0 A2.t1 221.719
R146 A2.n1 A2.t2 221.719
R147 A2.n0 A2.t0 149.419
R148 A2.n1 A2.t3 149.419
R149 A2.n2 A2.n1 33.447
R150 A2 A2.n2 31.809
R151 A2.n2 A2.n0 25.748
C0 B1 Y 0.31fF
C1 VPB VPWR 0.12fF
C2 VGND VPWR 0.13fF
C3 VGND Y 0.24fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__a41oi_4.ext - technology: sky130A

.subckt sky130_fd_sc_hd__a41oi_4 B1 A2 A1 A4 A3 Y VGND VPWR VNB VPB
X0 VPWR.t9 A1.t0 a_27_297.t9 VPB.t9 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_27_297.t14 A2.t0 VPWR.t12 VPB.t14 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 Y.t3 A1.t1 a_493_47.t7 VNB.t11 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 VPWR.t3 A4.t0 a_27_297.t3 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 Y.t2 A1.t2 a_493_47.t6 VNB.t10 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 a_27_297.t8 A1.t3 VPWR.t8 VPB.t8 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 VPWR.t13 A2.t1 a_27_297.t15 VPB.t15 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 a_27_297.t4 A3.t0 VPWR.t4 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 a_911_47.t3 A2.t2 a_493_47.t3 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 a_911_47.t7 A3.t1 a_1269_47.t7 VNB.t7 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 VGND.t3 A4.t1 a_1269_47.t3 VNB.t6 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 VPWR.t5 A3.t2 a_27_297.t5 VPB.t5 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 VGND.t2 A4.t2 a_1269_47.t2 VNB.t16 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 a_27_297.t16 B1.t0 Y.t10 VPB.t16 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14 a_493_47.t5 A1.t4 Y.t1 VNB.t9 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X15 a_493_47.t2 A2.t3 a_911_47.t2 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X16 a_493_47.t4 A1.t5 Y.t0 VNB.t8 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X17 a_493_47.t1 A2.t4 a_911_47.t1 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X18 Y.t11 B1.t1 a_27_297.t17 VPB.t17 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X19 a_27_297.t10 B1.t2 Y.t4 VPB.t10 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X20 VGND.t4 B1.t3 Y.t5 VNB.t12 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X21 VGND.t5 B1.t4 Y.t6 VNB.t13 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X22 a_911_47.t0 A2.t5 a_493_47.t0 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X23 a_1269_47.t1 A4.t3 VGND.t1 VNB.t17 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X24 a_27_297.t0 A3.t3 VPWR.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X25 a_27_297.t7 A1.t6 VPWR.t7 VPB.t7 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X26 VPWR.t1 A3.t4 a_27_297.t1 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X27 a_911_47.t6 A3.t5 a_1269_47.t6 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X28 Y.t7 B1.t5 VGND.t6 VNB.t14 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X29 a_27_297.t19 A2.t6 VPWR.t15 VPB.t19 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X30 VPWR.t2 A2.t7 a_27_297.t2 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X31 a_27_297.t12 A4.t4 VPWR.t10 VPB.t12 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X32 VPWR.t11 A4.t5 a_27_297.t13 VPB.t13 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X33 a_1269_47.t5 A3.t6 a_911_47.t5 VNB.t5 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X34 a_27_297.t18 A4.t6 VPWR.t14 VPB.t18 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X35 Y.t8 B1.t6 a_27_297.t11 VPB.t11 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X36 VPWR.t6 A1.t7 a_27_297.t6 VPB.t6 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X37 a_1269_47.t4 A3.t7 a_911_47.t4 VNB.t18 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X38 Y.t9 B1.t7 VGND.t7 VNB.t15 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X39 a_1269_47.t0 A4.t7 VGND.t0 VNB.t19 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
R0 A1.n11 A1.t0 238.369
R1 A1.n1 A1.t6 212.079
R2 A1.n4 A1.t7 212.079
R3 A1.n0 A1.t3 212.079
R4 A1.n1 A1.t5 139.779
R5 A1.n4 A1.t2 139.779
R6 A1.n0 A1.t4 139.779
R7 A1.n10 A1.t1 139.779
R8 A1.n2 A1 83.757
R9 A1.n6 A1.n5 76
R10 A1.n9 A1.n8 76
R11 A1.n12 A1.n11 76
R12 A1.n5 A1.n2 49.66
R13 A1.n4 A1.n3 46.739
R14 A1.n9 A1.n0 35.054
R15 A1.n10 A1.n9 26.29
R16 A1.n11 A1.n10 23.369
R17 A1.n3 A1.n0 14.606
R18 A1.n8 A1.n7 13.187
R19 A1 A1.n6 12.412
R20 A1.n12 A1 9.309
R21 A1.n2 A1.n1 8.763
R22 A1 A1.n12 8.533
R23 A1.n6 A1 5.43
R24 A1.n8 A1 3.878
R25 A1.n5 A1.n4 2.921
R26 A1.n7 A1 0.775
R27 a_27_297.n9 a_27_297.t11 624.727
R28 a_27_297.n13 a_27_297.n6 331.276
R29 a_27_297.n12 a_27_297.n7 309.441
R30 a_27_297.n11 a_27_297.n10 292.5
R31 a_27_297.n9 a_27_297.n8 292.5
R32 a_27_297.n2 a_27_297.t12 266.581
R33 a_27_297.n2 a_27_297.n1 168.571
R34 a_27_297.n3 a_27_297.n0 168.571
R35 a_27_297.n15 a_27_297.n4 168.571
R36 a_27_297.n14 a_27_297.n5 168.571
R37 a_27_297.n17 a_27_297.n16 168.57
R38 a_27_297.n12 a_27_297.n11 102.399
R39 a_27_297.n15 a_27_297.n14 95.247
R40 a_27_297.n10 a_27_297.t16 87.665
R41 a_27_297.n11 a_27_297.n9 86.588
R42 a_27_297.n13 a_27_297.n12 75.294
R43 a_27_297.n14 a_27_297.n13 70.4
R44 a_27_297.n3 a_27_297.n2 63.247
R45 a_27_297.n16 a_27_297.n3 63.247
R46 a_27_297.n16 a_27_297.n15 63.247
R47 a_27_297.n6 a_27_297.t15 45.31
R48 a_27_297.n4 a_27_297.t14 30.535
R49 a_27_297.n1 a_27_297.t13 26.595
R50 a_27_297.n1 a_27_297.t18 26.595
R51 a_27_297.n0 a_27_297.t3 26.595
R52 a_27_297.n0 a_27_297.t4 26.595
R53 a_27_297.n4 a_27_297.t1 26.595
R54 a_27_297.n5 a_27_297.t2 26.595
R55 a_27_297.n5 a_27_297.t19 26.595
R56 a_27_297.n6 a_27_297.t7 26.595
R57 a_27_297.n7 a_27_297.t6 26.595
R58 a_27_297.n7 a_27_297.t8 26.595
R59 a_27_297.n8 a_27_297.t17 26.595
R60 a_27_297.n8 a_27_297.t10 26.595
R61 a_27_297.n10 a_27_297.t9 26.595
R62 a_27_297.n17 a_27_297.t5 26.595
R63 a_27_297.t0 a_27_297.n17 26.595
R64 VPWR.n7 VPWR.n6 307.239
R65 VPWR.n35 VPWR.n34 292.5
R66 VPWR.n33 VPWR.n0 292.5
R67 VPWR.n9 VPWR.n8 167.719
R68 VPWR.n11 VPWR.n10 164.214
R69 VPWR.n18 VPWR.n17 164.214
R70 VPWR.n26 VPWR.n25 164.214
R71 VPWR.n31 VPWR.n30 164.214
R72 VPWR.n34 VPWR.n33 66.98
R73 VPWR.n4 VPWR.t2 66.98
R74 VPWR.n4 VPWR.t12 65.995
R75 VPWR.n20 VPWR.n19 34.635
R76 VPWR.n16 VPWR.n7 32.752
R77 VPWR.n12 VPWR.n11 26.729
R78 VPWR.n31 VPWR.n2 26.729
R79 VPWR.n34 VPWR.t8 26.595
R80 VPWR.n33 VPWR.t9 26.595
R81 VPWR.n8 VPWR.t10 26.595
R82 VPWR.n8 VPWR.t11 26.595
R83 VPWR.n10 VPWR.t14 26.595
R84 VPWR.n10 VPWR.t3 26.595
R85 VPWR.n6 VPWR.t4 26.595
R86 VPWR.n6 VPWR.t5 26.595
R87 VPWR.n17 VPWR.t0 26.595
R88 VPWR.n17 VPWR.t1 26.595
R89 VPWR.n25 VPWR.t15 26.595
R90 VPWR.n25 VPWR.t13 26.595
R91 VPWR.n30 VPWR.t7 26.595
R92 VPWR.n30 VPWR.t6 26.595
R93 VPWR.n26 VPWR.n24 25.6
R94 VPWR.n35 VPWR.n32 24.545
R95 VPWR.n24 VPWR.n23 19.102
R96 VPWR.n26 VPWR.n2 18.823
R97 VPWR.n32 VPWR.n31 17.694
R98 VPWR.n12 VPWR.n7 11.67
R99 VPWR.n20 VPWR.n4 8.205
R100 VPWR.n36 VPWR.n0 7.447
R101 VPWR.n38 VPWR.n0 7.382
R102 VPWR.n18 VPWR.n16 5.647
R103 VPWR.n37 VPWR.n36 4.65
R104 VPWR.n13 VPWR.n12 4.65
R105 VPWR.n14 VPWR.n7 4.65
R106 VPWR.n16 VPWR.n15 4.65
R107 VPWR.n19 VPWR.n5 4.65
R108 VPWR.n21 VPWR.n20 4.65
R109 VPWR.n23 VPWR.n22 4.65
R110 VPWR.n24 VPWR.n3 4.65
R111 VPWR.n27 VPWR.n26 4.65
R112 VPWR.n28 VPWR.n2 4.65
R113 VPWR.n31 VPWR.n29 4.65
R114 VPWR.n32 VPWR.n1 4.65
R115 VPWR.n19 VPWR.n18 4.141
R116 VPWR.n11 VPWR.n9 3.695
R117 VPWR.n23 VPWR.n4 1.15
R118 VPWR VPWR.n38 0.583
R119 VPWR.n36 VPWR.n35 0.465
R120 VPWR.n13 VPWR.n9 0.255
R121 VPWR.n38 VPWR.n37 0.134
R122 VPWR.n14 VPWR.n13 0.119
R123 VPWR.n15 VPWR.n14 0.119
R124 VPWR.n15 VPWR.n5 0.119
R125 VPWR.n21 VPWR.n5 0.119
R126 VPWR.n22 VPWR.n21 0.119
R127 VPWR.n22 VPWR.n3 0.119
R128 VPWR.n27 VPWR.n3 0.119
R129 VPWR.n28 VPWR.n27 0.119
R130 VPWR.n29 VPWR.n28 0.119
R131 VPWR.n29 VPWR.n1 0.119
R132 VPWR.n37 VPWR.n1 0.119
R133 VPB.t2 VPB.t14 488.317
R134 VPB.t9 VPB.t8 449.844
R135 VPB.t16 VPB.t9 432.087
R136 VPB.t7 VPB.t15 304.828
R137 VPB.t14 VPB.t1 260.436
R138 VPB.t13 VPB.t12 248.598
R139 VPB.t18 VPB.t13 248.598
R140 VPB.t3 VPB.t18 248.598
R141 VPB.t4 VPB.t3 248.598
R142 VPB.t5 VPB.t4 248.598
R143 VPB.t0 VPB.t5 248.598
R144 VPB.t1 VPB.t0 248.598
R145 VPB.t19 VPB.t2 248.598
R146 VPB.t15 VPB.t19 248.598
R147 VPB.t6 VPB.t7 248.598
R148 VPB.t8 VPB.t6 248.598
R149 VPB.t17 VPB.t16 248.598
R150 VPB.t10 VPB.t17 248.598
R151 VPB.t11 VPB.t10 248.598
R152 VPB VPB.t11 142.056
R153 A2.n0 A2.t0 218.601
R154 A2.n7 A2.t6 205.652
R155 A2.n4 A2.t1 205.652
R156 A2.n1 A2.t7 203.433
R157 A2.n4 A2.t2 152.861
R158 A2.n12 A2.t3 144.599
R159 A2.n6 A2.t4 139.779
R160 A2.n3 A2.t5 139.779
R161 A2 A2.n0 79.047
R162 A2.n14 A2.n13 76
R163 A2.n11 A2.n10 76
R164 A2.n9 A2.n8 76
R165 A2.n12 A2.n11 38.847
R166 A2.n5 A2.n4 29.608
R167 A2.n8 A2.n3 26.165
R168 A2.n9 A2.n2 20.723
R169 A2.n8 A2.n7 18.591
R170 A2 A2.n14 17.676
R171 A2.n10 A2 17.676
R172 A2.n6 A2.n5 15.148
R173 A2.n7 A2.n6 13.082
R174 A2.n3 A2.n1 12.251
R175 A2.n14 A2 10.361
R176 A2.n10 A2 10.361
R177 A2.n13 A2.n12 10.071
R178 A2.n11 A2.n1 7.821
R179 A2.n2 A2 4.266
R180 A2 A2.n9 3.047
R181 a_493_47.n4 a_493_47.t2 238.823
R182 a_493_47.n2 a_493_47.t7 238.823
R183 a_493_47.n3 a_493_47.n0 92.5
R184 a_493_47.n2 a_493_47.n1 92.5
R185 a_493_47.n5 a_493_47.n4 92.5
R186 a_493_47.n4 a_493_47.n3 63.247
R187 a_493_47.n3 a_493_47.n2 63.247
R188 a_493_47.n1 a_493_47.t6 24.923
R189 a_493_47.n1 a_493_47.t5 24.923
R190 a_493_47.n0 a_493_47.t3 24.923
R191 a_493_47.n0 a_493_47.t4 24.923
R192 a_493_47.t0 a_493_47.n5 24.923
R193 a_493_47.n5 a_493_47.t1 24.923
R194 Y.n2 Y.n0 187.498
R195 Y.n5 Y.n4 171.935
R196 Y.n8 Y.n6 155.747
R197 Y.n2 Y.n1 149.428
R198 Y.n5 Y.n3 105.676
R199 Y.n8 Y.n7 92.5
R200 Y.n9 Y.n8 64.376
R201 Y.n9 Y.n5 31.247
R202 Y Y.n2 27.952
R203 Y.n0 Y.t4 26.595
R204 Y.n0 Y.t8 26.595
R205 Y.n1 Y.t10 26.595
R206 Y.n1 Y.t11 26.595
R207 Y.n7 Y.t1 24.923
R208 Y.n7 Y.t3 24.923
R209 Y.n6 Y.t0 24.923
R210 Y.n6 Y.t2 24.923
R211 Y.n4 Y.t5 24.923
R212 Y.n4 Y.t9 24.923
R213 Y.n3 Y.t6 24.923
R214 Y.n3 Y.t7 24.923
R215 Y Y.n9 2.618
R216 VNB.t13 VNB.t11 5173.63
R217 VNB.t2 VNB.t4 4545.05
R218 VNB VNB.t15 3878.09
R219 VNB.t16 VNB.t17 2030.77
R220 VNB.t19 VNB.t16 2030.77
R221 VNB.t6 VNB.t19 2030.77
R222 VNB.t18 VNB.t6 2030.77
R223 VNB.t7 VNB.t18 2030.77
R224 VNB.t5 VNB.t7 2030.77
R225 VNB.t4 VNB.t5 2030.77
R226 VNB.t0 VNB.t2 2030.77
R227 VNB.t1 VNB.t0 2030.77
R228 VNB.t3 VNB.t1 2030.77
R229 VNB.t8 VNB.t3 2030.77
R230 VNB.t10 VNB.t8 2030.77
R231 VNB.t9 VNB.t10 2030.77
R232 VNB.t11 VNB.t9 2030.77
R233 VNB.t14 VNB.t13 2030.77
R234 VNB.t12 VNB.t14 2030.77
R235 VNB.t15 VNB.t12 2030.77
R236 A4.n0 A4.t4 212.079
R237 A4.n9 A4.t5 212.079
R238 A4.n3 A4.t6 212.079
R239 A4.n1 A4.t0 212.079
R240 A4.n0 A4.t3 139.779
R241 A4.n9 A4.t2 139.779
R242 A4.n3 A4.t7 139.779
R243 A4.n1 A4.t1 139.779
R244 A4 A4.n0 106.691
R245 A4.n11 A4.n10 76
R246 A4.n8 A4.n7 76
R247 A4.n6 A4.n4 76
R248 A4.n8 A4.n4 49.66
R249 A4.n3 A4.n2 48.2
R250 A4.n10 A4.n9 39.436
R251 A4.n6 A4.n5 21.229
R252 A4 A4.n11 20.604
R253 A4.n7 A4 15.609
R254 A4.n2 A4.n1 13.145
R255 A4.n7 A4 13.112
R256 A4.n9 A4.n8 10.224
R257 A4.n11 A4 8.117
R258 A4 A4.n6 5.619
R259 A4.n5 A4 1.873
R260 A4.n4 A4.n3 1.46
R261 A3.n8 A3.t2 205.652
R262 A3.n5 A3.t3 205.652
R263 A3.n2 A3.t4 205.652
R264 A3.n0 A3.t0 205.652
R265 A3.n0 A3.t7 144.599
R266 A3.n8 A3.t1 139.779
R267 A3.n5 A3.t6 139.779
R268 A3.n2 A3.t5 139.779
R269 A3 A3.n1 92.497
R270 A3.n10 A3.n9 76
R271 A3.n7 A3.n6 76
R272 A3.n4 A3.n3 76
R273 A3.n5 A3.n4 45.445
R274 A3.n1 A3.n0 21.582
R275 A3.n10 A3.n7 19.342
R276 A3.n3 A3 15.36
R277 A3.n4 A3.n2 12.394
R278 A3.n3 A3 10.808
R279 A3.n9 A3.n8 9.64
R280 A3.n7 A3 3.982
R281 A3 A3.n10 2.844
R282 A3.n6 A3.n5 1.377
R283 a_911_47.n5 a_911_47.n4 155.747
R284 a_911_47.n2 a_911_47.n0 155.747
R285 a_911_47.n4 a_911_47.n2 102.4
R286 a_911_47.n2 a_911_47.n1 92.5
R287 a_911_47.n4 a_911_47.n3 92.5
R288 a_911_47.n3 a_911_47.t2 24.923
R289 a_911_47.n3 a_911_47.t0 24.923
R290 a_911_47.n1 a_911_47.t5 24.923
R291 a_911_47.n1 a_911_47.t6 24.923
R292 a_911_47.n0 a_911_47.t4 24.923
R293 a_911_47.n0 a_911_47.t7 24.923
R294 a_911_47.n5 a_911_47.t1 24.923
R295 a_911_47.t3 a_911_47.n5 24.923
R296 a_1269_47.t6 a_1269_47.n5 238.823
R297 a_1269_47.n1 a_1269_47.t1 229.866
R298 a_1269_47.n1 a_1269_47.n0 108.688
R299 a_1269_47.n3 a_1269_47.n2 92.5
R300 a_1269_47.n5 a_1269_47.n4 92.5
R301 a_1269_47.n3 a_1269_47.n1 76.047
R302 a_1269_47.n5 a_1269_47.n3 63.247
R303 a_1269_47.n4 a_1269_47.t7 24.923
R304 a_1269_47.n4 a_1269_47.t5 24.923
R305 a_1269_47.n0 a_1269_47.t2 24.923
R306 a_1269_47.n0 a_1269_47.t0 24.923
R307 a_1269_47.n2 a_1269_47.t3 24.923
R308 a_1269_47.n2 a_1269_47.t4 24.923
R309 VGND.n33 VGND.t5 190.315
R310 VGND.n39 VGND.t7 190.095
R311 VGND.n11 VGND.n10 110.744
R312 VGND.n13 VGND.n12 107.239
R313 VGND.n37 VGND.n2 107.239
R314 VGND.n15 VGND.n14 34.635
R315 VGND.n15 VGND.n8 34.635
R316 VGND.n19 VGND.n8 34.635
R317 VGND.n20 VGND.n19 34.635
R318 VGND.n21 VGND.n20 34.635
R319 VGND.n21 VGND.n6 34.635
R320 VGND.n25 VGND.n6 34.635
R321 VGND.n26 VGND.n25 34.635
R322 VGND.n27 VGND.n26 34.635
R323 VGND.n27 VGND.n4 34.635
R324 VGND.n31 VGND.n4 34.635
R325 VGND.n32 VGND.n31 34.635
R326 VGND.n33 VGND.n32 32
R327 VGND.n14 VGND.n13 26.729
R328 VGND.n37 VGND.n1 25.976
R329 VGND.n10 VGND.t1 24.923
R330 VGND.n10 VGND.t2 24.923
R331 VGND.n12 VGND.t0 24.923
R332 VGND.n12 VGND.t3 24.923
R333 VGND.n2 VGND.t6 24.923
R334 VGND.n2 VGND.t4 24.923
R335 VGND.n39 VGND.n38 19.952
R336 VGND.n38 VGND.n37 18.447
R337 VGND.n33 VGND.n1 12.423
R338 VGND VGND.n39 4.65
R339 VGND.n14 VGND.n9 4.65
R340 VGND.n16 VGND.n15 4.65
R341 VGND.n17 VGND.n8 4.65
R342 VGND.n19 VGND.n18 4.65
R343 VGND.n20 VGND.n7 4.65
R344 VGND.n22 VGND.n21 4.65
R345 VGND.n23 VGND.n6 4.65
R346 VGND.n25 VGND.n24 4.65
R347 VGND.n26 VGND.n5 4.65
R348 VGND.n28 VGND.n27 4.65
R349 VGND.n29 VGND.n4 4.65
R350 VGND.n31 VGND.n30 4.65
R351 VGND.n32 VGND.n3 4.65
R352 VGND.n34 VGND.n33 4.65
R353 VGND.n35 VGND.n1 4.65
R354 VGND.n37 VGND.n36 4.65
R355 VGND.n38 VGND.n0 4.65
R356 VGND.n13 VGND.n11 3.695
R357 VGND.n11 VGND.n9 0.255
R358 VGND.n16 VGND.n9 0.119
R359 VGND.n17 VGND.n16 0.119
R360 VGND.n18 VGND.n17 0.119
R361 VGND.n18 VGND.n7 0.119
R362 VGND.n22 VGND.n7 0.119
R363 VGND.n23 VGND.n22 0.119
R364 VGND.n24 VGND.n23 0.119
R365 VGND.n24 VGND.n5 0.119
R366 VGND.n28 VGND.n5 0.119
R367 VGND.n29 VGND.n28 0.119
R368 VGND.n30 VGND.n29 0.119
R369 VGND.n30 VGND.n3 0.119
R370 VGND.n34 VGND.n3 0.119
R371 VGND.n35 VGND.n34 0.119
R372 VGND.n36 VGND.n35 0.119
R373 VGND.n36 VGND.n0 0.119
R374 VGND VGND.n0 0.119
R375 B1.n0 B1.t0 212.079
R376 B1.n1 B1.t1 212.079
R377 B1.n4 B1.t2 212.079
R378 B1.n7 B1.t6 212.079
R379 B1.n0 B1.t4 139.779
R380 B1.n1 B1.t5 139.779
R381 B1.n4 B1.t3 139.779
R382 B1.n7 B1.t7 139.779
R383 B1.n3 B1.n2 76
R384 B1.n6 B1.n5 76
R385 B1.n9 B1.n8 76
R386 B1.n1 B1.n0 61.345
R387 B1.n5 B1.n3 49.66
R388 B1.n8 B1.n7 20.448
R389 B1.n9 B1.n6 18.921
R390 B1 B1.n11 18.643
R391 B1.n2 B1 13.078
R392 B1.n2 B1 12.521
R393 B1.n5 B1.n4 8.763
R394 B1.n10 B1 8.145
R395 B1.n6 B1 6.4
R396 B1.n10 B1 3.895
R397 B1.n11 B1.n10 3.06
R398 B1.n3 B1.n1 2.921
R399 B1 B1.n9 0.278
C0 VGND VPWR 0.22fF
C1 VGND Y 0.35fF
C2 Y A1 0.30fF
C3 B1 Y 0.41fF
C4 VPB VPWR 0.19fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__a211o_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__a211o_1 VGND VPWR X A2 B1 A1 C1 VNB VPB
X0 VPWR.t1 a_80_21.t4 X.t0 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_80_21.t2 C1.t0 a_472_297.t0 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 VPWR.t0 A2.t0 a_217_297.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 VGND.t3 B1.t0 a_80_21.t0 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 VGND.t2 a_80_21.t5 X.t1 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 a_300_47.t1 A2.t1 VGND.t1 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 a_217_297.t1 A1.t0 VPWR.t2 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 a_80_21.t1 A1.t1 a_300_47.t0 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 a_472_297.t1 B1.t1 a_217_297.t2 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 a_80_21.t3 C1.t1 VGND.t0 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
R0 a_80_21.t2 a_80_21.n3 354.605
R1 a_80_21.n0 a_80_21.t4 231.014
R2 a_80_21.n2 a_80_21.t3 177.965
R3 a_80_21.n0 a_80_21.t5 158.714
R4 a_80_21.n3 a_80_21.n2 102.069
R5 a_80_21.n2 a_80_21.n1 92.5
R6 a_80_21.n3 a_80_21.n0 76
R7 a_80_21.n1 a_80_21.t0 25.846
R8 a_80_21.n1 a_80_21.t1 25.846
R9 X.n1 X.t0 541.537
R10 X X.t0 527.204
R11 X.n0 X.t1 82.027
R12 X.n1 X 7.832
R13 X X.n0 6.906
R14 X X.n1 6.167
R15 X.n0 X 5.674
R16 VPWR.n1 VPWR.n0 310.027
R17 VPWR.n1 VPWR.t1 195.138
R18 VPWR.n0 VPWR.t2 27.58
R19 VPWR.n0 VPWR.t0 27.58
R20 VPWR VPWR.n1 0.217
R21 VPB.t2 VPB.t0 562.305
R22 VPB.t4 VPB.t1 272.274
R23 VPB.t3 VPB.t4 254.517
R24 VPB.t0 VPB.t3 254.517
R25 VPB VPB.t2 201.246
R26 C1.n0 C1.t0 231.014
R27 C1.n0 C1.t1 158.714
R28 C1 C1.n0 78.607
R29 a_472_297.t0 a_472_297.t1 61.07
R30 A2.n0 A2.t0 231.014
R31 A2.n0 A2.t1 158.714
R32 A2 A2.n0 81.43
R33 a_217_297.t0 a_217_297.n0 365.578
R34 a_217_297.n0 a_217_297.t2 27.58
R35 a_217_297.n0 a_217_297.t1 27.58
R36 B1.n0 B1.t1 241.534
R37 B1.n0 B1.t0 169.234
R38 B1 B1.n0 81.042
R39 VGND.n3 VGND.n0 110.205
R40 VGND.n2 VGND.n1 92.5
R41 VGND.n5 VGND.n4 92.5
R42 VGND.n1 VGND.t1 40.615
R43 VGND.n4 VGND.t2 40.615
R44 VGND.n0 VGND.t0 28.615
R45 VGND.n0 VGND.t3 28.615
R46 VGND.n6 VGND.n5 5.987
R47 VGND.n3 VGND.n2 4.446
R48 VGND.n6 VGND.n3 0.162
R49 VGND VGND.n6 0.129
R50 VNB VNB.t3 6150.61
R51 VNB.t3 VNB.t2 4593.41
R52 VNB.t4 VNB.t1 2224.18
R53 VNB.t0 VNB.t4 2079.12
R54 VNB.t2 VNB.t0 2079.12
R55 a_300_47.t0 a_300_47.t1 51.692
R56 A1.n0 A1.t0 241.534
R57 A1.n0 A1.t1 169.234
R58 A1 A1.n0 88.024
C0 X VPWR 0.13fF
C1 A2 A1 0.11fF
C2 B1 C1 0.11fF
C3 A1 B1 0.11fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__a211o_2.ext - technology: sky130A

.subckt sky130_fd_sc_hd__a211o_2 X A2 A1 B1 C1 VGND VPWR VNB VPB
X0 a_79_21.t0 A1.t0 a_348_47.t0 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 a_79_21.t2 C1.t0 VGND.t2 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 VGND.t4 a_79_21.t4 X.t3 VNB.t5 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 VPWR.t3 a_79_21.t5 X.t1 VPB.t5 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 a_79_21.t3 C1.t1 a_585_297.t0 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 VPWR.t1 A2.t0 a_299_297.t0 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 a_299_297.t1 A1.t1 VPWR.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 a_585_297.t1 B1.t0 a_299_297.t2 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 a_348_47.t1 A2.t1 VGND.t0 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 X.t0 a_79_21.t6 VPWR.t2 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 X.t2 a_79_21.t7 VGND.t3 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 VGND.t1 B1.t1 a_79_21.t1 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
R0 A1.n0 A1.t1 239.038
R1 A1.n0 A1.t0 166.738
R2 A1 A1.n0 92.973
R3 a_348_47.t0 a_348_47.t1 75.692
R4 a_79_21.n2 a_79_21.t4 1296.58
R5 a_79_21.t3 a_79_21.n5 346.634
R6 a_79_21.n1 a_79_21.t5 212.079
R7 a_79_21.n0 a_79_21.t6 212.079
R8 a_79_21.n0 a_79_21.t7 141.386
R9 a_79_21.n4 a_79_21.t2 136.734
R10 a_79_21.n5 a_79_21.n2 85.64
R11 a_79_21.n5 a_79_21.n4 84.105
R12 a_79_21.n1 a_79_21.n0 62.289
R13 a_79_21.n4 a_79_21.n3 52.624
R14 a_79_21.n3 a_79_21.t1 39.692
R15 a_79_21.n3 a_79_21.t0 25.846
R16 a_79_21.n2 a_79_21.n1 19.28
R17 VNB VNB.t4 6053.91
R18 VNB.t5 VNB.t1 3698.9
R19 VNB.t1 VNB.t0 2707.69
R20 VNB.t0 VNB.t2 2441.76
R21 VNB.t2 VNB.t3 2320.88
R22 VNB.t4 VNB.t5 2079.12
R23 C1.n0 C1.t1 230.154
R24 C1.n0 C1.t0 157.854
R25 C1 C1.n0 79.895
R26 VGND.n3 VGND.n0 113.053
R27 VGND.n10 VGND.t3 108.016
R28 VGND.n2 VGND.n1 92.5
R29 VGND.n5 VGND.n4 92.5
R30 VGND.n0 VGND.t2 30.461
R31 VGND.n0 VGND.t1 30.461
R32 VGND.n1 VGND.t0 24.923
R33 VGND.n4 VGND.t4 24.923
R34 VGND.n3 VGND.n2 7.732
R35 VGND.n11 VGND.n10 4.65
R36 VGND.n7 VGND.n6 4.65
R37 VGND.n9 VGND.n8 4.65
R38 VGND.n6 VGND.n5 0.966
R39 VGND.n7 VGND.n3 0.147
R40 VGND.n9 VGND.n7 0.119
R41 VGND.n11 VGND.n9 0.119
R42 VGND VGND.n11 0.02
R43 X.n2 X.n1 140.375
R44 X.n2 X.n0 110.316
R45 X.n1 X.t1 26.595
R46 X.n1 X.t0 26.595
R47 X.n0 X.t3 26.262
R48 X.n0 X.t2 25.427
R49 X X.n2 15.091
R50 VPWR.n2 VPWR.n0 313.113
R51 VPWR.n1 VPWR.t3 196.066
R52 VPWR.n5 VPWR.t2 148.63
R53 VPWR.n0 VPWR.t1 39.4
R54 VPWR.n0 VPWR.t0 37.43
R55 VPWR.n4 VPWR.n3 4.65
R56 VPWR.n6 VPWR.n5 4.65
R57 VPWR.n2 VPWR.n1 3.955
R58 VPWR.n4 VPWR.n2 0.207
R59 VPWR.n6 VPWR.n4 0.119
R60 VPWR VPWR.n6 0.02
R61 VPB.t5 VPB.t1 556.386
R62 VPB.t1 VPB.t0 319.626
R63 VPB.t0 VPB.t3 284.112
R64 VPB.t4 VPB.t5 248.598
R65 VPB.t3 VPB.t2 213.084
R66 VPB VPB.t4 189.408
R67 a_585_297.t0 a_585_297.t1 41.37
R68 A2.n0 A2.t1 929.507
R69 A2.n0 A2.t0 232.213
R70 A2 A2.n0 82.956
R71 a_299_297.t0 a_299_297.n0 379.331
R72 a_299_297.n0 a_299_297.t1 36.445
R73 a_299_297.n0 a_299_297.t2 28.565
R74 B1.n0 B1.t0 241.534
R75 B1.n0 B1.t1 169.234
R76 B1 B1.n0 82.121
C0 VPWR X 0.17fF
C1 X VGND 0.16fF
C2 VPWR VGND 0.10fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__a211o_4.ext - technology: sky130A

.subckt sky130_fd_sc_hd__a211o_4 VGND VPWR C1 B1 X A2 A1 VNB VPB
X0 X.t3 a_79_204.t8 VPWR.t5 VPB.t7 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 VPWR.t0 A1.t0 a_473_297.t3 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 a_473_297.t2 A1.t1 VPWR.t1 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 X.t7 a_79_204.t9 VGND.t7 VNB sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 VGND.t9 C1.t0 a_79_204.t7 VNB sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 a_79_204.t2 B1.t0 VGND.t2 VNB sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 VPWR.t4 a_79_204.t10 X.t2 VPB.t6 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 a_473_297.t4 A2.t0 VPWR.t6 VPB.t10 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 a_473_297.t0 B1.t1 a_727_297.t1 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 X.t6 a_79_204.t11 VGND.t6 VNB sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 VGND.t3 B1.t2 a_79_204.t3 VNB sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 a_79_204.t4 C1.t1 VGND.t8 VNB sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 VGND.t5 a_79_204.t12 X.t5 VNB sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 a_1123_47.t1 A1.t2 a_79_204.t0 VNB sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14 a_555_297.t1 B1.t3 a_473_297.t1 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 VPWR.t7 A2.t1 a_473_297.t5 VPB.t11 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16 VGND.t0 A2.t2 a_1123_47.t0 VNB sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X17 a_951_47.t0 A2.t3 VGND.t1 VNB sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X18 VPWR.t3 a_79_204.t13 X.t1 VPB.t5 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X19 VGND.t4 a_79_204.t14 X.t4 VNB sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X20 a_79_204.t1 A1.t3 a_951_47.t1 VNB sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X21 a_79_204.t5 C1.t2 a_555_297.t0 VPB.t8 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X22 a_727_297.t0 C1.t3 a_79_204.t6 VPB.t9 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X23 X.t0 a_79_204.t15 VPWR.t2 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
R0 a_79_204.n18 a_79_204.n17 400.504
R1 a_79_204.n5 a_79_204.t15 243.482
R2 a_79_204.n15 a_79_204.t12 207.697
R3 a_79_204.n15 a_79_204.t10 204.046
R4 a_79_204.n11 a_79_204.t8 204.046
R5 a_79_204.n7 a_79_204.t13 204.046
R6 a_79_204.n6 a_79_204.t9 147.813
R7 a_79_204.n10 a_79_204.t14 147.813
R8 a_79_204.n14 a_79_204.t11 147.813
R9 a_79_204.n2 a_79_204.n0 130.82
R10 a_79_204.n4 a_79_204.n3 92.5
R11 a_79_204.n9 a_79_204.n5 91.542
R12 a_79_204.n13 a_79_204.n12 76
R13 a_79_204.n9 a_79_204.n8 76
R14 a_79_204.n16 a_79_204.n15 76
R15 a_79_204.n4 a_79_204.n2 53.164
R16 a_79_204.n17 a_79_204.n4 49.97
R17 a_79_204.n2 a_79_204.n1 46.25
R18 a_79_204.n1 a_79_204.t4 36.923
R19 a_79_204.n1 a_79_204.t3 35.076
R20 a_79_204.n3 a_79_204.t7 33.23
R21 a_79_204.n18 a_79_204.t6 27.58
R22 a_79_204.t5 a_79_204.n18 27.58
R23 a_79_204.n8 a_79_204.n7 26.29
R24 a_79_204.n3 a_79_204.t2 25.846
R25 a_79_204.n0 a_79_204.t0 25.846
R26 a_79_204.n0 a_79_204.t1 25.846
R27 a_79_204.n17 a_79_204.n16 23.542
R28 a_79_204.n16 a_79_204.n13 15.542
R29 a_79_204.n13 a_79_204.n9 15.542
R30 a_79_204.n12 a_79_204.n11 13.145
R31 a_79_204.n15 a_79_204.n14 5.112
R32 a_79_204.n11 a_79_204.n10 5.112
R33 a_79_204.n7 a_79_204.n6 5.112
R34 VPWR.n3 VPWR.n0 310.018
R35 VPWR.n2 VPWR.n1 306.463
R36 VPWR.n14 VPWR.t4 196.528
R37 VPWR.n24 VPWR.t2 190.907
R38 VPWR.n20 VPWR.n19 164.584
R39 VPWR.n1 VPWR.t1 49.25
R40 VPWR.n19 VPWR.t5 27.58
R41 VPWR.n19 VPWR.t3 27.58
R42 VPWR.n1 VPWR.t7 27.58
R43 VPWR.n0 VPWR.t6 27.58
R44 VPWR.n0 VPWR.t0 27.58
R45 VPWR.n5 VPWR.n4 4.65
R46 VPWR.n7 VPWR.n6 4.65
R47 VPWR.n9 VPWR.n8 4.65
R48 VPWR.n11 VPWR.n10 4.65
R49 VPWR.n13 VPWR.n12 4.65
R50 VPWR.n16 VPWR.n15 4.65
R51 VPWR.n18 VPWR.n17 4.65
R52 VPWR.n21 VPWR.n20 4.65
R53 VPWR.n23 VPWR.n22 4.65
R54 VPWR.n25 VPWR.n24 4.65
R55 VPWR.n3 VPWR.n2 3.922
R56 VPWR.n15 VPWR.n14 0.752
R57 VPWR.n5 VPWR.n3 0.218
R58 VPWR.n7 VPWR.n5 0.119
R59 VPWR.n9 VPWR.n7 0.119
R60 VPWR.n11 VPWR.n9 0.119
R61 VPWR.n13 VPWR.n11 0.119
R62 VPWR.n16 VPWR.n13 0.119
R63 VPWR.n18 VPWR.n16 0.119
R64 VPWR.n21 VPWR.n18 0.119
R65 VPWR.n23 VPWR.n21 0.119
R66 VPWR.n25 VPWR.n23 0.119
R67 VPWR VPWR.n25 0.022
R68 X.n2 X.n1 215.904
R69 X.n2 X.n0 163.941
R70 X.n5 X.n4 148.458
R71 X.n5 X.n3 105.636
R72 X X.n2 62.941
R73 X X.n5 39.577
R74 X.n4 X.t5 28.615
R75 X.n1 X.t2 27.58
R76 X.n1 X.t3 27.58
R77 X.n0 X.t1 27.58
R78 X.n0 X.t0 27.58
R79 X.n3 X.t4 25.846
R80 X.n3 X.t7 25.846
R81 X.n4 X.t6 25.846
R82 VPB.t6 VPB.t3 556.386
R83 VPB.t11 VPB.t1 319.626
R84 VPB.t2 VPB.t11 319.626
R85 VPB.t9 VPB.t2 278.193
R86 VPB.t0 VPB.t10 254.517
R87 VPB.t1 VPB.t0 254.517
R88 VPB.t8 VPB.t9 254.517
R89 VPB.t3 VPB.t8 254.517
R90 VPB.t7 VPB.t6 254.517
R91 VPB.t5 VPB.t7 254.517
R92 VPB.t4 VPB.t5 254.517
R93 VPB VPB.t4 192.367
R94 A1.n0 A1.t0 204.046
R95 A1.n1 A1.t1 204.046
R96 A1.n0 A1.t2 147.813
R97 A1.n1 A1.t3 147.813
R98 A1 A1.n2 78.04
R99 A1.n2 A1.n0 49.66
R100 A1.n2 A1.n1 13.145
R101 a_473_297.n1 a_473_297.t1 649.657
R102 a_473_297.n2 a_473_297.t4 313.864
R103 a_473_297.n3 a_473_297.n2 307.761
R104 a_473_297.n1 a_473_297.n0 143.121
R105 a_473_297.n2 a_473_297.n1 47.132
R106 a_473_297.n0 a_473_297.t5 41.37
R107 a_473_297.n0 a_473_297.t0 35.46
R108 a_473_297.t3 a_473_297.n3 27.58
R109 a_473_297.n3 a_473_297.t2 27.58
R110 VGND.n20 VGND.t7 188.748
R111 VGND.n2 VGND.t0 107.823
R112 VGND.n6 VGND.n5 106.463
R113 VGND.n16 VGND.n15 106.463
R114 VGND.n11 VGND.n10 106.255
R115 VGND.n1 VGND.n0 92.5
R116 VGND.n0 VGND.t1 46.153
R117 VGND.n0 VGND.t3 33.23
R118 VGND.n5 VGND.t8 33.23
R119 VGND.n5 VGND.t9 28.615
R120 VGND.n10 VGND.t5 26.769
R121 VGND.n10 VGND.t2 25.846
R122 VGND.n15 VGND.t6 25.846
R123 VGND.n15 VGND.t4 25.846
R124 VGND.n4 VGND.n3 4.65
R125 VGND.n7 VGND.n6 4.65
R126 VGND.n9 VGND.n8 4.65
R127 VGND.n12 VGND.n11 4.65
R128 VGND.n14 VGND.n13 4.65
R129 VGND.n17 VGND.n16 4.65
R130 VGND.n19 VGND.n18 4.65
R131 VGND.n2 VGND.n1 4.354
R132 VGND.n21 VGND.n20 3.876
R133 VGND.n4 VGND.n2 0.139
R134 VGND.n21 VGND.n19 0.139
R135 VGND VGND.n21 0.122
R136 VGND.n7 VGND.n4 0.119
R137 VGND.n9 VGND.n7 0.119
R138 VGND.n12 VGND.n9 0.119
R139 VGND.n14 VGND.n12 0.119
R140 VGND.n17 VGND.n14 0.119
R141 VGND.n19 VGND.n17 0.119
R142 C1.n0 C1.t3 202.439
R143 C1.n1 C1.t2 202.439
R144 C1.n1 C1.t0 145.436
R145 C1.n0 C1.t1 138.173
R146 C1 C1.n2 32.873
R147 C1.n2 C1.n0 27.696
R148 C1.n2 C1.n1 19.574
R149 B1.n1 B1.t1 231.797
R150 B1.n0 B1.t3 231.797
R151 B1.n0 B1.t0 168.261
R152 B1.n1 B1.t2 162.126
R153 B1 B1.n0 148.47
R154 B1 B1.n1 87.054
R155 A2.n1 A2.t0 231.797
R156 A2.n0 A2.t1 223.033
R157 A2.n0 A2.t3 168.261
R158 A2.n1 A2.t2 166.508
R159 A2 A2.n0 157.58
R160 A2 A2.n1 97.272
R161 a_727_297.t0 a_727_297.t1 63.04
R162 a_1123_47.t0 a_1123_47.t1 51.692
R163 a_555_297.t0 a_555_297.t1 55.16
R164 a_951_47.t0 a_951_47.t1 51.692
C0 VPB VPWR 0.13fF
C1 VGND VPWR 0.14fF
C2 X VPWR 0.53fF
C3 B1 C1 0.37fF
C4 X VGND 0.35fF
C5 A1 A2 0.27fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__a211oi_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__a211oi_1 A1 C1 B1 Y A2 VPWR VGND VNB VPB
X0 a_56_297.t0 A1.t0 VPWR.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 VPWR.t1 A2.t0 a_56_297.t1 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 Y.t1 C1.t0 VGND.t0 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 a_139_47.t1 A2.t1 VGND.t1 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 a_311_297.t1 B1.t0 a_56_297.t2 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 Y.t0 C1.t1 a_311_297.t0 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 VGND.t2 B1.t1 Y.t3 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 Y.t2 A1.t1 a_139_47.t0 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
R0 A1.n0 A1.t0 241.534
R1 A1.n0 A1.t1 169.234
R2 A1.n1 A1.n0 76
R3 A1.n2 A1.n1 12.024
R4 A1.n2 A1 11.776
R5 A1 A1.n2 4.848
R6 A1.n1 A1 0.969
R7 VPWR VPWR.n0 166.831
R8 VPWR.n0 VPWR.t0 27.58
R9 VPWR.n0 VPWR.t1 27.58
R10 a_56_297.n0 a_56_297.t1 398.771
R11 a_56_297.n0 a_56_297.t2 27.58
R12 a_56_297.t0 a_56_297.n0 27.58
R13 VPB VPB.t1 281.152
R14 VPB.t3 VPB.t2 272.274
R15 VPB.t0 VPB.t3 254.517
R16 VPB.t1 VPB.t0 254.517
R17 A2.n0 A2.t0 228.647
R18 A2.n0 A2.t1 156.347
R19 A2 A2.n0 78.07
R20 C1.n0 C1.t1 231.014
R21 C1.n0 C1.t0 158.714
R22 C1.n1 C1.n0 76
R23 C1.n1 C1 12.16
R24 C1 C1.n1 2.346
R25 VGND.n1 VGND.t1 168.187
R26 VGND.n1 VGND.n0 110.131
R27 VGND.n0 VGND.t0 28.615
R28 VGND.n0 VGND.t2 28.615
R29 VGND VGND.n1 0.052
R30 Y.n2 Y.t0 173.83
R31 Y.n1 Y.n0 154.283
R32 Y.n1 Y.t1 118.346
R33 Y.n0 Y.t3 25.846
R34 Y.n0 Y.t2 25.846
R35 Y Y.n1 16.703
R36 Y.n2 Y 5.54
R37 Y Y.n2 3.247
R38 VNB VNB.t2 6803.36
R39 VNB.t3 VNB.t0 2224.18
R40 VNB.t1 VNB.t3 2079.12
R41 VNB.t2 VNB.t1 2079.12
R42 a_139_47.t0 a_139_47.t1 51.692
R43 B1.n0 B1.t0 241.534
R44 B1.n0 B1.t1 169.234
R45 B1.n1 B1.n0 76
R46 B1 B1.n1 13.078
R47 B1.n1 B1 2.133
R48 a_311_297.t0 a_311_297.t1 61.07
C0 A1 B1 0.11fF
C1 B1 C1 0.13fF
C2 Y C1 0.18fF
C3 Y B1 0.19fF
C4 VPWR Y 0.13fF
C5 VGND Y 0.24fF
C6 A2 A1 0.16fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__a211oi_2.ext - technology: sky130A

.subckt sky130_fd_sc_hd__a211oi_2 A2 C1 B1 Y A1 VPWR VGND VNB VPB
X0 VGND.t3 A2.t0 a_485_47.t1 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 VPWR.t1 A1.t0 a_292_297.t1 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 a_37_297.t1 B1.t0 a_292_297.t5 VPB.t7 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 Y.t5 B1.t1 VGND.t4 VNB.t6 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 a_485_47.t0 A2.t1 VGND.t2 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 a_292_297.t2 A2.t2 VPWR.t3 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 VGND.t5 B1.t2 Y.t4 VNB.t7 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 VPWR.t2 A2.t3 a_292_297.t3 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 a_485_47.t2 A1.t1 Y.t1 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 VGND.t0 C1.t0 Y.t2 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 Y.t3 C1.t1 VGND.t1 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 a_37_297.t2 C1.t2 Y.t6 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 Y.t0 A1.t2 a_485_47.t3 VNB.t5 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 Y.t7 C1.t3 a_37_297.t3 VPB.t5 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14 a_292_297.t0 A1.t3 VPWR.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 a_292_297.t4 B1.t3 a_37_297.t0 VPB.t6 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
R0 A2.n0 A2.t3 212.079
R1 A2.n1 A2.t2 212.079
R2 A2.n0 A2.t1 139.779
R3 A2.n1 A2.t0 139.779
R4 A2.n4 A2.n0 106.672
R5 A2.n3 A2.n2 76
R6 A2.n2 A2.n1 43.818
R7 A2.n4 A2.n3 12.8
R8 A2.n4 A2 11.224
R9 A2.n3 A2 5.12
R10 A2 A2.n4 2.166
R11 a_485_47.n1 a_485_47.t3 230.945
R12 a_485_47.t0 a_485_47.n1 180.949
R13 a_485_47.n1 a_485_47.n0 92.5
R14 a_485_47.n0 a_485_47.t1 25.846
R15 a_485_47.n0 a_485_47.t2 25.846
R16 VGND.n1 VGND.t5 188.748
R17 VGND.n10 VGND.t1 148.554
R18 VGND.n2 VGND.n0 110.29
R19 VGND.n6 VGND.n5 107.239
R20 VGND.n0 VGND.t2 25.846
R21 VGND.n0 VGND.t3 25.846
R22 VGND.n5 VGND.t4 25.846
R23 VGND.n5 VGND.t0 25.846
R24 VGND.n11 VGND.n10 4.65
R25 VGND.n4 VGND.n3 4.65
R26 VGND.n7 VGND.n6 4.65
R27 VGND.n9 VGND.n8 4.65
R28 VGND.n2 VGND.n1 3.998
R29 VGND.n4 VGND.n2 0.139
R30 VGND.n7 VGND.n4 0.119
R31 VGND.n9 VGND.n7 0.119
R32 VGND.n11 VGND.n9 0.119
R33 VGND VGND.n11 0.027
R34 VNB VNB.t1 6440.72
R35 VNB.t7 VNB.t5 4593.41
R36 VNB.t3 VNB.t2 2079.12
R37 VNB.t4 VNB.t3 2079.12
R38 VNB.t5 VNB.t4 2079.12
R39 VNB.t6 VNB.t7 2079.12
R40 VNB.t0 VNB.t6 2079.12
R41 VNB.t1 VNB.t0 2079.12
R42 A1.n0 A1.t0 212.079
R43 A1.n1 A1.t3 212.079
R44 A1.n0 A1.t1 139.779
R45 A1.n1 A1.t2 139.779
R46 A1.n4 A1.n2 76
R47 A1.n2 A1.n0 43.818
R48 A1.n2 A1.n1 18.987
R49 A1.n4 A1.n3 17.408
R50 A1.n3 A1 5.632
R51 A1 A1.n4 0.512
R52 a_292_297.n2 a_292_297.n0 222.279
R53 a_292_297.n2 a_292_297.n1 146.859
R54 a_292_297.n3 a_292_297.n2 109.1
R55 a_292_297.n1 a_292_297.t3 27.58
R56 a_292_297.n1 a_292_297.t2 27.58
R57 a_292_297.n0 a_292_297.t5 27.58
R58 a_292_297.n0 a_292_297.t4 27.58
R59 a_292_297.n3 a_292_297.t1 27.58
R60 a_292_297.t0 a_292_297.n3 27.58
R61 VPWR.n2 VPWR.t2 203.499
R62 VPWR.n5 VPWR.t0 199.56
R63 VPWR.n1 VPWR.n0 171.98
R64 VPWR.n0 VPWR.t3 27.58
R65 VPWR.n0 VPWR.t1 27.58
R66 VPWR.n4 VPWR.n3 4.65
R67 VPWR.n6 VPWR.n5 4.039
R68 VPWR.n2 VPWR.n1 3.963
R69 VPWR VPWR.n6 0.607
R70 VPWR.n4 VPWR.n2 0.233
R71 VPWR.n6 VPWR.n4 0.137
R72 VPB.t7 VPB.t0 562.305
R73 VPB.t3 VPB.t2 254.517
R74 VPB.t1 VPB.t3 254.517
R75 VPB.t0 VPB.t1 254.517
R76 VPB.t6 VPB.t7 254.517
R77 VPB.t4 VPB.t6 254.517
R78 VPB.t5 VPB.t4 254.517
R79 VPB VPB.t5 236.76
R80 B1.n0 B1.t0 212.079
R81 B1.n1 B1.t3 212.079
R82 B1.n0 B1.t2 139.779
R83 B1.n1 B1.t1 139.779
R84 B1 B1.n2 80.864
R85 B1.n2 B1.n0 31.403
R86 B1.n2 B1.n1 31.403
R87 B1 B1.n3 18.432
R88 B1.n3 B1 9.309
R89 B1.n3 B1 5.12
R90 a_37_297.n1 a_37_297.t3 238.364
R91 a_37_297.t1 a_37_297.n1 227.26
R92 a_37_297.n1 a_37_297.n0 151.212
R93 a_37_297.n0 a_37_297.t0 27.58
R94 a_37_297.n0 a_37_297.t2 27.58
R95 Y.n6 Y.n5 180.82
R96 Y.n1 Y.n0 146.685
R97 Y Y.n2 92.746
R98 Y.n4 Y.n3 92.5
R99 Y.n8 Y.n2 92.5
R100 Y.n7 Y.n6 47.68
R101 Y.n0 Y.t6 27.58
R102 Y.n0 Y.t7 27.58
R103 Y.n5 Y.t1 25.846
R104 Y.n5 Y.t0 25.846
R105 Y.n3 Y.t4 25.846
R106 Y.n3 Y.t5 25.846
R107 Y.n2 Y.t2 25.846
R108 Y.n2 Y.t3 25.846
R109 Y.n7 Y 15.894
R110 Y Y.n1 12.384
R111 Y.n4 Y 9.768
R112 Y.n6 Y.n4 5.726
R113 Y.n1 Y 3.095
R114 Y Y.n8 0.228
R115 Y.n8 Y.n7 0.228
R116 C1.n0 C1.t2 212.079
R117 C1.n1 C1.t3 212.079
R118 C1.n0 C1.t0 139.779
R119 C1.n1 C1.t1 139.779
R120 C1.n2 C1.n1 106.672
R121 C1.n1 C1.n0 62.806
R122 C1.n2 C1 11.96
R123 C1 C1.n2 2.308
C0 A1 Y 0.17fF
C1 Y VGND 0.44fF
C2 Y B1 0.27fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__a211oi_4.ext - technology: sky130A

.subckt sky130_fd_sc_hd__a211oi_4 A2 A1 C1 Y B1 VPWR VGND VNB VPB
X0 Y.t6 A1.t0 a_109_47.t7 VNB.t10 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 VGND.t3 C1.t0 Y.t7 VNB.t11 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 VGND.t6 A2.t0 a_109_47.t1 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 VGND.t11 B1.t0 Y.t15 VNB.t15 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 VPWR.t7 A1.t1 a_27_297.t9 VPB.t15 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 a_27_297.t8 A1.t2 VPWR.t6 VPB.t14 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 VPWR.t3 A2.t1 a_27_297.t3 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 a_949_297.t0 B1.t1 a_27_297.t7 VPB.t7 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 a_27_297.t2 A2.t2 VPWR.t2 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 Y.t8 C1.t1 a_949_297.t1 VPB.t11 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 a_781_297.t3 C1.t2 Y.t9 VPB.t10 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 a_27_297.t5 B1.t2 a_781_297.t1 VPB.t6 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 VGND.t7 A2.t3 a_109_47.t2 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 Y.t5 A1.t3 a_109_47.t6 VNB.t9 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14 a_781_297.t0 B1.t3 a_27_297.t4 VPB.t5 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 a_1301_297.t1 C1.t3 Y.t10 VPB.t9 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16 a_27_297.t1 A2.t4 VPWR.t1 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17 Y.t11 C1.t4 a_781_297.t2 VPB.t8 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X18 a_109_47.t3 A2.t5 VGND.t8 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X19 a_109_47.t5 A1.t4 Y.t4 VNB.t8 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X20 Y.t12 C1.t5 VGND.t2 VNB.t12 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X21 VPWR.t5 A1.t5 a_27_297.t11 VPB.t13 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X22 a_109_47.t4 A1.t6 Y.t3 VNB.t7 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X23 Y.t13 C1.t6 VGND.t1 VNB.t13 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X24 Y.t1 B1.t4 VGND.t9 VNB.t5 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X25 a_27_297.t10 A1.t7 VPWR.t4 VPB.t12 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X26 Y.t2 B1.t5 VGND.t10 VNB.t6 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X27 VPWR.t0 A2.t6 a_27_297.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X28 a_27_297.t6 B1.t6 a_1301_297.t0 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X29 VGND.t0 C1.t7 Y.t14 VNB.t14 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X30 a_109_47.t0 A2.t7 VGND.t5 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X31 VGND.t4 B1.t7 Y.t0 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
R0 A1.n0 A1.t5 221.719
R1 A1.n2 A1.t7 221.719
R2 A1.n5 A1.t1 221.719
R3 A1.n8 A1.t2 221.719
R4 A1.n0 A1.t6 149.419
R5 A1.n2 A1.t0 149.419
R6 A1.n5 A1.t4 149.419
R7 A1.n8 A1.t3 149.419
R8 A1.n4 A1.n1 94.133
R9 A1 A1.n9 85.066
R10 A1.n4 A1.n3 76
R11 A1.n7 A1.n6 76
R12 A1.n1 A1.n0 26.777
R13 A1.n7 A1.n4 18.133
R14 A1.n9 A1.n8 16.066
R15 A1.n3 A1.n2 12.496
R16 A1 A1.n7 9.066
R17 A1.n6 A1.n5 1.785
R18 a_109_47.n5 a_109_47.n4 155.927
R19 a_109_47.n2 a_109_47.n0 135.508
R20 a_109_47.n4 a_109_47.n3 92.5
R21 a_109_47.n2 a_109_47.n1 92.5
R22 a_109_47.n4 a_109_47.n2 43.008
R23 a_109_47.n0 a_109_47.t1 24.923
R24 a_109_47.n0 a_109_47.t4 24.923
R25 a_109_47.n1 a_109_47.t7 24.923
R26 a_109_47.n1 a_109_47.t5 24.923
R27 a_109_47.n3 a_109_47.t6 24.923
R28 a_109_47.n3 a_109_47.t3 24.923
R29 a_109_47.n5 a_109_47.t2 24.923
R30 a_109_47.t0 a_109_47.n5 24.923
R31 Y.n2 Y.n1 343.7
R32 Y.n2 Y.n0 292.5
R33 Y.n8 Y.n7 149.089
R34 Y Y.n13 94.12
R35 Y.n8 Y.n6 92.5
R36 Y.n13 Y.n3 92.5
R37 Y.n10 Y.n8 79.26
R38 Y.n11 Y.n5 49.651
R39 Y.n12 Y.n4 49.651
R40 Y.n10 Y.n9 49.045
R41 Y Y.n2 48.649
R42 Y.n13 Y.n12 46.396
R43 Y.n12 Y.n11 44.437
R44 Y.n11 Y.n10 39.593
R45 Y.n9 Y.t15 33.23
R46 Y.n0 Y.t11 31.52
R47 Y.n9 Y.t1 28.615
R48 Y.n1 Y.t9 27.58
R49 Y.n1 Y.t8 27.58
R50 Y.n0 Y.t10 27.58
R51 Y.n3 Y.t13 26.769
R52 Y.n5 Y.t2 25.846
R53 Y.n3 Y.t0 24.923
R54 Y.n4 Y.t7 24.923
R55 Y.n4 Y.t12 24.923
R56 Y.n5 Y.t14 24.923
R57 Y.n6 Y.t3 24.923
R58 Y.n6 Y.t6 24.923
R59 Y.n7 Y.t4 24.923
R60 Y.n7 Y.t5 24.923
R61 VNB VNB.t1 6053.91
R62 VNB.t5 VNB.t15 2345.05
R63 VNB.t13 VNB.t0 2079.12
R64 VNB.t15 VNB.t6 2079.12
R65 VNB.t6 VNB.t14 2054.95
R66 VNB.t11 VNB.t13 2030.77
R67 VNB.t12 VNB.t11 2030.77
R68 VNB.t14 VNB.t12 2030.77
R69 VNB.t2 VNB.t5 2030.77
R70 VNB.t7 VNB.t2 2030.77
R71 VNB.t10 VNB.t7 2030.77
R72 VNB.t8 VNB.t10 2030.77
R73 VNB.t9 VNB.t8 2030.77
R74 VNB.t4 VNB.t9 2030.77
R75 VNB.t3 VNB.t4 2030.77
R76 VNB.t1 VNB.t3 2030.77
R77 C1.n11 C1.t1 218.651
R78 C1.n0 C1.t3 212.079
R79 C1.n3 C1.t4 212.079
R80 C1.n7 C1.t2 212.079
R81 C1.n0 C1.t6 139.779
R82 C1.n10 C1.t7 139.779
R83 C1.n6 C1.t5 139.779
R84 C1.n2 C1.t0 139.779
R85 C1.n5 C1.n1 94.133
R86 C1 C1.n11 78.4
R87 C1.n5 C1.n4 76
R88 C1.n9 C1.n8 76
R89 C1.n1 C1.n0 35.784
R90 C1.n4 C1.n3 19.718
R91 C1.n9 C1.n5 18.133
R92 C1 C1.n9 15.733
R93 C1.n8 C1.n7 6.572
R94 C1.n7 C1.n6 5.842
R95 C1.n3 C1.n2 4.381
R96 C1.n11 C1.n10 0.73
R97 VGND.n2 VGND.t4 192.143
R98 VGND.n32 VGND.t5 191.789
R99 VGND.n16 VGND.n15 113.205
R100 VGND.n28 VGND.n27 112.108
R101 VGND.n1 VGND.n0 106.463
R102 VGND.n6 VGND.n5 106.463
R103 VGND.n11 VGND.n10 106.463
R104 VGND.n10 VGND.t10 25.846
R105 VGND.n10 VGND.t11 25.846
R106 VGND.n0 VGND.t1 24.923
R107 VGND.n0 VGND.t3 24.923
R108 VGND.n5 VGND.t2 24.923
R109 VGND.n5 VGND.t0 24.923
R110 VGND.n15 VGND.t9 24.923
R111 VGND.n15 VGND.t6 24.923
R112 VGND.n27 VGND.t8 24.923
R113 VGND.n27 VGND.t7 24.923
R114 VGND.n17 VGND.n16 12.8
R115 VGND.n33 VGND.n32 4.65
R116 VGND.n4 VGND.n3 4.65
R117 VGND.n7 VGND.n6 4.65
R118 VGND.n9 VGND.n8 4.65
R119 VGND.n12 VGND.n11 4.65
R120 VGND.n14 VGND.n13 4.65
R121 VGND.n18 VGND.n17 4.65
R122 VGND.n20 VGND.n19 4.65
R123 VGND.n22 VGND.n21 4.65
R124 VGND.n24 VGND.n23 4.65
R125 VGND.n26 VGND.n25 4.65
R126 VGND.n29 VGND.n28 4.65
R127 VGND.n31 VGND.n30 4.65
R128 VGND.n2 VGND.n1 3.791
R129 VGND.n4 VGND.n2 0.261
R130 VGND.n7 VGND.n4 0.119
R131 VGND.n9 VGND.n7 0.119
R132 VGND.n12 VGND.n9 0.119
R133 VGND.n14 VGND.n12 0.119
R134 VGND.n18 VGND.n14 0.119
R135 VGND.n20 VGND.n18 0.119
R136 VGND.n22 VGND.n20 0.119
R137 VGND.n24 VGND.n22 0.119
R138 VGND.n26 VGND.n24 0.119
R139 VGND.n29 VGND.n26 0.119
R140 VGND.n31 VGND.n29 0.119
R141 VGND.n33 VGND.n31 0.119
R142 VGND VGND.n33 0.02
R143 A2.n0 A2.t4 241.534
R144 A2.n3 A2.n0 226.39
R145 A2.n1 A2.t1 221.719
R146 A2.n5 A2.t2 221.719
R147 A2.n4 A2.t6 221.719
R148 A2.n0 A2.t0 169.234
R149 A2.n1 A2.t5 149.419
R150 A2.n5 A2.t3 149.419
R151 A2.n4 A2.t7 149.419
R152 A2.n3 A2.n2 76
R153 A2.n6 A2.n4 35.492
R154 A2 A2.n6 32.916
R155 A2.n6 A2.n5 22.746
R156 A2.n2 A2.n1 16.066
R157 A2 A2.n3 3.254
R158 B1.n0 B1.t6 240.999
R159 B1.n4 B1.t2 212.079
R160 B1.n1 B1.t1 212.079
R161 B1.n6 B1.t3 212.079
R162 B1.n0 B1.t7 168.699
R163 B1.n1 B1.t5 150.733
R164 B1.n6 B1.t4 139.779
R165 B1.n3 B1.t0 139.779
R166 B1.n9 B1.n0 105.233
R167 B1.n5 B1.n2 87.567
R168 B1.n8 B1.n7 76.11
R169 B1.n5 B1.n4 76
R170 B1.n2 B1.n1 11.684
R171 B1.n7 B1.n6 11.684
R172 B1.n4 B1.n3 9.493
R173 B1.n8 B1.n5 7.393
R174 B1.n9 B1.n8 4.65
R175 B1 B1.n9 0.046
R176 a_27_297.n2 a_27_297.t6 722.394
R177 a_27_297.n2 a_27_297.n1 292.5
R178 a_27_297.t0 a_27_297.n9 212.804
R179 a_27_297.n9 a_27_297.n8 149.831
R180 a_27_297.n7 a_27_297.n6 149.831
R181 a_27_297.n5 a_27_297.n4 149.831
R182 a_27_297.n3 a_27_297.n0 143.481
R183 a_27_297.n3 a_27_297.n2 56.741
R184 a_27_297.n5 a_27_297.n3 40.224
R185 a_27_297.n7 a_27_297.n5 34.683
R186 a_27_297.n9 a_27_297.n7 34.683
R187 a_27_297.n1 a_27_297.t7 26.595
R188 a_27_297.n1 a_27_297.t5 26.595
R189 a_27_297.n0 a_27_297.t4 26.595
R190 a_27_297.n0 a_27_297.t1 26.595
R191 a_27_297.n4 a_27_297.t11 26.595
R192 a_27_297.n4 a_27_297.t10 26.595
R193 a_27_297.n6 a_27_297.t9 26.595
R194 a_27_297.n6 a_27_297.t8 26.595
R195 a_27_297.n8 a_27_297.t3 26.595
R196 a_27_297.n8 a_27_297.t2 26.595
R197 VPWR.n3 VPWR.n2 310.69
R198 VPWR.n12 VPWR.n11 307.239
R199 VPWR.n1 VPWR.n0 306.463
R200 VPWR.n7 VPWR.n6 306.463
R201 VPWR.n2 VPWR.t1 26.595
R202 VPWR.n2 VPWR.t5 26.595
R203 VPWR.n0 VPWR.t4 26.595
R204 VPWR.n0 VPWR.t7 26.595
R205 VPWR.n6 VPWR.t6 26.595
R206 VPWR.n6 VPWR.t3 26.595
R207 VPWR.n11 VPWR.t2 26.595
R208 VPWR.n11 VPWR.t0 26.595
R209 VPWR.n5 VPWR.n4 4.65
R210 VPWR.n8 VPWR.n7 4.65
R211 VPWR.n10 VPWR.n9 4.65
R212 VPWR.n3 VPWR.n1 4.222
R213 VPWR.n13 VPWR.n12 3.932
R214 VPWR.n5 VPWR.n3 0.42
R215 VPWR.n13 VPWR.n10 0.137
R216 VPWR VPWR.n13 0.121
R217 VPWR.n8 VPWR.n5 0.119
R218 VPWR.n10 VPWR.n8 0.119
R219 VPB.t9 VPB.t4 272.274
R220 VPB.t8 VPB.t9 266.355
R221 VPB.t7 VPB.t11 266.355
R222 VPB.t10 VPB.t8 254.517
R223 VPB.t11 VPB.t10 254.517
R224 VPB.t6 VPB.t7 248.598
R225 VPB.t5 VPB.t6 248.598
R226 VPB.t1 VPB.t5 248.598
R227 VPB.t13 VPB.t1 248.598
R228 VPB.t12 VPB.t13 248.598
R229 VPB.t15 VPB.t12 248.598
R230 VPB.t14 VPB.t15 248.598
R231 VPB.t3 VPB.t14 248.598
R232 VPB.t2 VPB.t3 248.598
R233 VPB.t0 VPB.t2 248.598
R234 VPB VPB.t0 189.408
R235 a_949_297.t0 a_949_297.t1 59.1
R236 a_781_297.n1 a_781_297.n0 669.75
R237 a_781_297.n0 a_781_297.t2 27.58
R238 a_781_297.n0 a_781_297.t3 27.58
R239 a_781_297.t1 a_781_297.n1 26.595
R240 a_781_297.n1 a_781_297.t0 26.595
R241 a_1301_297.t0 a_1301_297.t1 61.07
C0 VPB VPWR 0.13fF
C1 A2 B1 0.17fF
C2 Y VGND 0.68fF
C3 A1 Y 0.22fF
C4 B1 VPWR 0.17fF
C5 B1 C1 0.22fF
C6 A2 A1 0.51fF
C7 VPWR VGND 0.10fF
C8 B1 VGND 0.13fF
C9 C1 Y 0.44fF
C10 B1 Y 0.45fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__a221o_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__a221o_1 X B1 A1 B2 A2 VGND VPWR C1 VNB VPB
X0 a_465_47.t1 A1.t0 a_27_47.t2 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 X.t1 a_27_47.t4 VPWR.t2 VPB.t5 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 a_109_297.t1 B1.t0 a_193_297.t3 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 a_193_297.t0 B2.t0 a_109_297.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 X.t0 a_27_47.t5 VGND.t3 VNB.t5 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 a_205_47.t0 B2.t1 VGND.t0 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 VPWR.t0 A2.t0 a_193_297.t1 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 a_193_297.t2 A1.t1 VPWR.t1 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 a_27_47.t0 B1.t1 a_205_47.t1 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 a_109_297.t2 C1.t0 a_27_47.t3 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 VGND.t1 C1.t1 a_27_47.t1 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 VGND.t2 A2.t1 a_465_47.t0 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
R0 A1.n0 A1.t1 236.549
R1 A1.n0 A1.t0 164.249
R2 A1 A1.n0 78.47
R3 a_27_47.t3 a_27_47.n3 523.051
R4 a_27_47.n0 a_27_47.t4 241.534
R5 a_27_47.n1 a_27_47.t1 233.992
R6 a_27_47.n0 a_27_47.t5 169.234
R7 a_27_47.n1 a_27_47.t0 157.115
R8 a_27_47.n2 a_27_47.t2 157.115
R9 a_27_47.n3 a_27_47.n2 108.528
R10 a_27_47.n3 a_27_47.n0 76
R11 a_27_47.n2 a_27_47.n1 26.624
R12 a_465_47.t0 a_465_47.t1 60.923
R13 VNB VNB.t2 6053.91
R14 VNB.t1 VNB.t4 4545.05
R15 VNB.t4 VNB.t3 2320.88
R16 VNB.t2 VNB.t0 2320.88
R17 VNB.t3 VNB.t5 2248.35
R18 VNB.t0 VNB.t1 1740.66
R19 VPWR.n1 VPWR.t1 546.316
R20 VPWR.n2 VPWR.n0 169.305
R21 VPWR.n0 VPWR.t0 35.46
R22 VPWR.n9 VPWR 33.261
R23 VPWR.n0 VPWR.t2 26.595
R24 VPWR VPWR.n8 6.023
R25 VPWR.n6 VPWR.n5 4.65
R26 VPWR.n8 VPWR.n7 4.65
R27 VPWR.n4 VPWR.n3 4.65
R28 VPWR.n2 VPWR.n1 3.849
R29 VPWR.n4 VPWR.n2 0.23
R30 VPWR.n6 VPWR.n4 0.119
R31 VPWR.n7 VPWR.n6 0.119
R32 VPWR.n9 VPWR.n7 0.119
R33 VPWR VPWR.n9 0.02
R34 X.n0 X.t1 172.967
R35 X X.t0 157.365
R36 X.n1 X.n0 102.923
R37 X X.n1 11.07
R38 X.n1 X 8.031
R39 X.n0 X 4.145
R40 VPB.t2 VPB.t3 556.386
R41 VPB.t3 VPB.t1 284.112
R42 VPB.t1 VPB.t5 275.233
R43 VPB.t0 VPB.t2 248.598
R44 VPB.t4 VPB.t0 248.598
R45 VPB VPB.t4 189.408
R46 B1.n0 B1.t0 239.503
R47 B1.n0 B1.t1 167.203
R48 B1 B1.n0 81.12
R49 a_193_297.n1 a_193_297.n0 514.223
R50 a_193_297.n0 a_193_297.t1 33.49
R51 a_193_297.n0 a_193_297.t2 31.52
R52 a_193_297.n1 a_193_297.t3 26.595
R53 a_193_297.t0 a_193_297.n1 26.595
R54 a_109_297.n0 a_109_297.t1 762.514
R55 a_109_297.t0 a_109_297.n0 26.595
R56 a_109_297.n0 a_109_297.t2 26.595
R57 B2.n0 B2.t0 241.534
R58 B2.n0 B2.t1 169.234
R59 B2 B2.n0 93.92
R60 VGND.n3 VGND.n2 112.002
R61 VGND.n1 VGND.n0 109.566
R62 VGND.n0 VGND.t0 36
R63 VGND.n2 VGND.t3 33.23
R64 VGND.n0 VGND.t1 24.923
R65 VGND.n2 VGND.t2 24.923
R66 VGND.n3 VGND.n1 3.418
R67 VGND.n1 VGND 3.296
R68 VGND VGND.n3 0.142
R69 a_205_47.t0 a_205_47.t1 38.769
R70 A2.n0 A2.t0 241.534
R71 A2.n0 A2.t1 169.234
R72 A2 A2.n0 88.8
R73 C1.n0 C1.t0 231.716
R74 C1.n0 C1.t1 159.416
R75 C1 C1.n0 83.619
C0 VPWR X 0.14fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__a221o_2.ext - technology: sky130A

.subckt sky130_fd_sc_hd__a221o_2 X B1 A1 B2 A2 VGND VPWR C1 VNB VPB
X0 VPWR.t1 a_27_47.t4 X.t1 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_465_47.t0 A1.t0 a_27_47.t2 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 X.t0 a_27_47.t5 VPWR.t0 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 a_109_297.t2 B1.t0 a_193_297.t3 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 a_193_297.t2 B2.t0 a_109_297.t1 VPB.t6 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 X.t3 a_27_47.t6 VGND.t2 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 a_205_47.t0 B2.t1 VGND.t4 VNB.t6 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 VPWR.t3 A2.t0 a_193_297.t1 VPB.t5 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 a_193_297.t0 A1.t1 VPWR.t2 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 a_27_47.t3 B1.t1 a_205_47.t1 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 VGND.t1 a_27_47.t7 X.t2 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 a_109_297.t0 C1.t0 a_27_47.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 VGND.t0 C1.t1 a_27_47.t1 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 VGND.t3 A2.t1 a_465_47.t1 VNB.t5 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
R0 a_27_47.t0 a_27_47.n4 523.051
R1 a_27_47.n2 a_27_47.t1 233.992
R2 a_27_47.n0 a_27_47.t4 212.079
R3 a_27_47.n1 a_27_47.t5 212.079
R4 a_27_47.n2 a_27_47.t3 157.115
R5 a_27_47.n3 a_27_47.t2 157.115
R6 a_27_47.n0 a_27_47.t7 139.779
R7 a_27_47.n1 a_27_47.t6 139.779
R8 a_27_47.n4 a_27_47.n3 108.528
R9 a_27_47.n4 a_27_47.n1 82.572
R10 a_27_47.n1 a_27_47.n0 61.345
R11 a_27_47.n3 a_27_47.n2 26.624
R12 X.n1 X.n0 146.372
R13 X.n3 X.n1 102.923
R14 X X.n2 92.75
R15 X.n0 X.t1 26.595
R16 X.n0 X.t0 26.595
R17 X.n2 X.t2 24.923
R18 X.n2 X.t3 24.923
R19 X X.n3 11.07
R20 X.n3 X 8.031
R21 X.n1 X 4.145
R22 VPWR.n5 VPWR.t2 546.316
R23 VPWR.n2 VPWR.t1 171.49
R24 VPWR.n1 VPWR.n0 165.765
R25 VPWR.n0 VPWR.t3 35.46
R26 VPWR.n13 VPWR 33.261
R27 VPWR.n0 VPWR.t0 26.595
R28 VPWR VPWR.n12 6.023
R29 VPWR.n4 VPWR.n3 4.65
R30 VPWR.n6 VPWR.n5 4.65
R31 VPWR.n10 VPWR.n9 4.65
R32 VPWR.n12 VPWR.n11 4.65
R33 VPWR.n8 VPWR.n7 4.65
R34 VPWR.n2 VPWR.n1 3.779
R35 VPWR.n4 VPWR.n2 0.305
R36 VPWR.n6 VPWR.n4 0.119
R37 VPWR.n8 VPWR.n6 0.119
R38 VPWR.n10 VPWR.n8 0.119
R39 VPWR.n11 VPWR.n10 0.119
R40 VPWR.n13 VPWR.n11 0.119
R41 VPWR VPWR.n13 0.02
R42 VPB.t4 VPB.t3 556.386
R43 VPB.t3 VPB.t5 284.112
R44 VPB.t5 VPB.t1 275.233
R45 VPB.t1 VPB.t2 248.598
R46 VPB.t6 VPB.t4 248.598
R47 VPB.t0 VPB.t6 248.598
R48 VPB VPB.t0 189.408
R49 A1.n0 A1.t1 236.549
R50 A1.n0 A1.t0 164.249
R51 A1 A1.n0 78.47
R52 a_465_47.t0 a_465_47.t1 60.923
R53 VNB VNB.t1 6053.91
R54 VNB.t4 VNB.t0 4545.05
R55 VNB.t0 VNB.t5 2320.88
R56 VNB.t1 VNB.t6 2320.88
R57 VNB.t5 VNB.t3 2248.35
R58 VNB.t3 VNB.t2 2030.77
R59 VNB.t6 VNB.t4 1740.66
R60 B1.n0 B1.t0 239.503
R61 B1.n0 B1.t1 167.203
R62 B1 B1.n0 81.12
R63 a_193_297.n1 a_193_297.n0 514.222
R64 a_193_297.n1 a_193_297.t1 33.49
R65 a_193_297.t0 a_193_297.n1 31.52
R66 a_193_297.n0 a_193_297.t3 26.595
R67 a_193_297.n0 a_193_297.t2 26.595
R68 a_109_297.n0 a_109_297.t2 762.514
R69 a_109_297.n0 a_109_297.t1 26.595
R70 a_109_297.t0 a_109_297.n0 26.595
R71 B2.n0 B2.t0 241.534
R72 B2.n0 B2.t1 169.234
R73 B2 B2.n0 93.92
R74 VGND.n2 VGND.t1 110.999
R75 VGND.n12 VGND.n11 109.566
R76 VGND.n1 VGND.n0 108.015
R77 VGND.n11 VGND.t4 36
R78 VGND.n0 VGND.t2 33.23
R79 VGND.n11 VGND.t0 24.923
R80 VGND.n0 VGND.t3 24.923
R81 VGND.n4 VGND.n3 4.65
R82 VGND.n6 VGND.n5 4.65
R83 VGND.n8 VGND.n7 4.65
R84 VGND.n10 VGND.n9 4.65
R85 VGND.n13 VGND.n12 3.932
R86 VGND.n2 VGND.n1 3.863
R87 VGND.n12 VGND 3.296
R88 VGND.n4 VGND.n2 0.287
R89 VGND.n13 VGND.n10 0.138
R90 VGND VGND.n13 0.122
R91 VGND.n6 VGND.n4 0.119
R92 VGND.n8 VGND.n6 0.119
R93 VGND.n10 VGND.n8 0.119
R94 a_205_47.t0 a_205_47.t1 38.769
R95 A2.n0 A2.t0 241.534
R96 A2.n0 A2.t1 169.234
R97 A2 A2.n0 88.8
R98 C1.n0 C1.t0 231.716
R99 C1.n0 C1.t1 159.416
R100 C1 C1.n0 83.619
C0 VPWR X 0.31fF
C1 VGND X 0.20fF
C2 VGND VPWR 0.11fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__a221o_4.ext - technology: sky130A

.subckt sky130_fd_sc_hd__a221o_4 A1 B1 C1 B2 X A2 VPWR VGND VNB VPB
X0 VGND.t6 A2.t0 a_445_47.t1 VNB.t7 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 VGND.t8 B2.t0 a_1053_47.t2 VNB.t12 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 a_804_297.t5 B1.t0 a_445_297.t5 VPB.t8 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 a_79_21.t1 A1.t0 a_445_47.t2 VNB.t9 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 a_445_297.t3 A2.t1 VPWR.t7 VPB.t6 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 a_804_297.t2 C1.t0 a_79_21.t2 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 a_445_297.t4 B1.t1 a_804_297.t4 VPB.t7 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 VPWR.t5 a_79_21.t8 X.t3 VPB.t9 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 a_1053_47.t1 B2.t1 VGND.t9 VNB.t13 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 a_79_21.t3 C1.t1 a_804_297.t3 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 a_1053_47.t0 B1.t2 a_79_21.t7 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 X.t2 a_79_21.t9 VPWR.t4 VPB.t10 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 a_445_47.t3 A1.t1 a_79_21.t0 VNB.t11 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 VGND.t3 C1.t2 a_79_21.t4 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14 VPWR.t3 a_79_21.t10 X.t1 VPB.t11 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 VGND.t7 a_79_21.t11 X.t7 VNB.t10 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X16 VGND.t0 a_79_21.t12 X.t6 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X17 a_804_297.t1 B2.t2 a_445_297.t1 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X18 a_79_21.t6 B1.t3 a_1053_47.t3 VNB.t8 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X19 a_79_21.t5 C1.t3 VGND.t4 VNB.t5 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X20 a_445_297.t0 B2.t3 a_804_297.t0 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X21 X.t5 a_79_21.t13 VGND.t1 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X22 a_445_47.t0 A2.t2 VGND.t5 VNB.t6 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X23 a_445_297.t6 A1.t2 VPWR.t1 VPB.t12 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X24 VPWR.t6 A2.t3 a_445_297.t2 VPB.t5 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X25 VPWR.t0 A1.t3 a_445_297.t7 VPB.t13 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X26 X.t0 a_79_21.t14 VPWR.t2 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X27 X.t4 a_79_21.t15 VGND.t2 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
R0 A2.n0 A2.t3 212.079
R1 A2.n1 A2.t1 212.079
R2 A2.n0 A2.t0 139.779
R3 A2.n1 A2.t2 139.779
R4 A2 A2.n2 77.696
R5 A2.n2 A2.n1 40.896
R6 A2.n2 A2.n0 20.448
R7 a_445_47.n1 a_445_47.n0 175.689
R8 a_445_47.n0 a_445_47.t2 24.923
R9 a_445_47.n0 a_445_47.t3 24.923
R10 a_445_47.n1 a_445_47.t1 24.923
R11 a_445_47.t0 a_445_47.n1 24.923
R12 VGND.n10 VGND.t6 219.525
R13 VGND.n27 VGND.t2 193.925
R14 VGND.n1 VGND.n0 124.063
R15 VGND.n3 VGND.n2 115.464
R16 VGND.n16 VGND.n15 115.464
R17 VGND.n22 VGND.n21 115.464
R18 VGND.n0 VGND.t9 24.923
R19 VGND.n0 VGND.t8 24.923
R20 VGND.n2 VGND.t4 24.923
R21 VGND.n2 VGND.t3 24.923
R22 VGND.n15 VGND.t5 24.923
R23 VGND.n15 VGND.t0 24.923
R24 VGND.n21 VGND.t1 24.923
R25 VGND.n21 VGND.t7 24.923
R26 VGND.n11 VGND.n10 15.811
R27 VGND.n4 VGND.n3 14.305
R28 VGND.n17 VGND.n16 9.788
R29 VGND.n28 VGND.n27 6.908
R30 VGND.n5 VGND.n4 4.65
R31 VGND.n7 VGND.n6 4.65
R32 VGND.n9 VGND.n8 4.65
R33 VGND.n12 VGND.n11 4.65
R34 VGND.n14 VGND.n13 4.65
R35 VGND.n18 VGND.n17 4.65
R36 VGND.n20 VGND.n19 4.65
R37 VGND.n24 VGND.n23 4.65
R38 VGND.n26 VGND.n25 4.65
R39 VGND.n23 VGND.n22 3.764
R40 VGND.n5 VGND.n1 0.134
R41 VGND.n7 VGND.n5 0.119
R42 VGND.n9 VGND.n7 0.119
R43 VGND.n12 VGND.n9 0.119
R44 VGND.n14 VGND.n12 0.119
R45 VGND.n18 VGND.n14 0.119
R46 VGND.n20 VGND.n18 0.119
R47 VGND.n24 VGND.n20 0.119
R48 VGND.n26 VGND.n24 0.119
R49 VGND.n28 VGND.n26 0.119
R50 VGND VGND.n28 0.019
R51 VNB VNB.t3 6029.73
R52 VNB.t8 VNB.t12 4545.05
R53 VNB.t7 VNB.t11 4545.05
R54 VNB.t12 VNB.t13 2030.77
R55 VNB.t0 VNB.t8 2030.77
R56 VNB.t5 VNB.t0 2030.77
R57 VNB.t4 VNB.t5 2030.77
R58 VNB.t9 VNB.t4 2030.77
R59 VNB.t11 VNB.t9 2030.77
R60 VNB.t6 VNB.t7 2030.77
R61 VNB.t1 VNB.t6 2030.77
R62 VNB.t2 VNB.t1 2030.77
R63 VNB.t10 VNB.t2 2030.77
R64 VNB.t3 VNB.t10 2030.77
R65 B2.n3 B2.t3 218.651
R66 B2.n0 B2.t2 212.079
R67 B2.n0 B2.t1 152.924
R68 B2.n2 B2.t0 139.779
R69 B2 B2.n1 92.152
R70 B2 B2.n3 80.571
R71 B2.n3 B2.n2 6.572
R72 B2.n1 B2.n0 5.112
R73 a_1053_47.t2 a_1053_47.n1 175.576
R74 a_1053_47.n1 a_1053_47.n0 138.776
R75 a_1053_47.n1 a_1053_47.t1 136.341
R76 a_1053_47.n0 a_1053_47.t3 24.923
R77 a_1053_47.n0 a_1053_47.t0 24.923
R78 B1.n0 B1.t0 212.079
R79 B1.n2 B1.t1 212.079
R80 B1.n2 B1.t2 141.382
R81 B1.n1 B1.t3 139.779
R82 B1.n4 B1.n3 76
R83 B1.n3 B1.n2 48.2
R84 B1 B1.n4 17.371
R85 B1.n3 B1.n1 11.684
R86 B1.n1 B1.n0 1.46
R87 a_445_297.n5 a_445_297.n4 237.912
R88 a_445_297.n2 a_445_297.n0 198.996
R89 a_445_297.n2 a_445_297.n1 154.412
R90 a_445_297.n4 a_445_297.n2 146.54
R91 a_445_297.n4 a_445_297.n3 143.026
R92 a_445_297.n1 a_445_297.t6 27.58
R93 a_445_297.n0 a_445_297.t2 26.595
R94 a_445_297.n0 a_445_297.t3 26.595
R95 a_445_297.n1 a_445_297.t7 26.595
R96 a_445_297.n3 a_445_297.t5 26.595
R97 a_445_297.n3 a_445_297.t4 26.595
R98 a_445_297.n5 a_445_297.t1 26.595
R99 a_445_297.t0 a_445_297.n5 26.595
R100 a_804_297.n2 a_804_297.t3 569.933
R101 a_804_297.n2 a_804_297.n1 292.5
R102 a_804_297.t1 a_804_297.n5 228.169
R103 a_804_297.n3 a_804_297.n0 146.25
R104 a_804_297.n5 a_804_297.n4 146.25
R105 a_804_297.n3 a_804_297.n2 40.279
R106 a_804_297.n4 a_804_297.t0 26.595
R107 a_804_297.n0 a_804_297.t5 26.595
R108 a_804_297.n1 a_804_297.t4 26.595
R109 a_804_297.n1 a_804_297.t2 26.595
R110 a_804_297.n5 a_804_297.n3 8.023
R111 VPB.t13 VPB.t4 559.345
R112 VPB.t8 VPB.t1 497.196
R113 VPB.t12 VPB.t13 251.557
R114 VPB.t1 VPB.t2 248.598
R115 VPB.t7 VPB.t8 248.598
R116 VPB.t3 VPB.t7 248.598
R117 VPB.t4 VPB.t3 248.598
R118 VPB.t5 VPB.t12 248.598
R119 VPB.t6 VPB.t5 248.598
R120 VPB.t9 VPB.t6 248.598
R121 VPB.t10 VPB.t9 248.598
R122 VPB.t11 VPB.t10 248.598
R123 VPB.t0 VPB.t11 248.598
R124 VPB VPB.t0 186.448
R125 A1.n3 A1.t2 216.46
R126 A1.n0 A1.t3 212.079
R127 A1.n2 A1.t0 147.812
R128 A1.n1 A1.t1 139.779
R129 A1 A1.n2 78.133
R130 A1.n4 A1.n3 76
R131 A1 A1.n4 55.261
R132 A1.n2 A1.n1 53.312
R133 A1.n1 A1.n0 13.875
R134 A1.n4 A1 6.4
R135 a_79_21.n12 a_79_21.n0 292.5
R136 a_79_21.n16 a_79_21.t0 235.764
R137 a_79_21.n14 a_79_21.t6 228.739
R138 a_79_21.n12 a_79_21.n11 223.459
R139 a_79_21.n9 a_79_21.t8 212.079
R140 a_79_21.n6 a_79_21.t9 212.079
R141 a_79_21.n3 a_79_21.t10 212.079
R142 a_79_21.n1 a_79_21.t14 212.079
R143 a_79_21.n9 a_79_21.t12 139.779
R144 a_79_21.n6 a_79_21.t13 139.779
R145 a_79_21.n3 a_79_21.t11 139.779
R146 a_79_21.n1 a_79_21.t15 139.779
R147 a_79_21.n5 a_79_21.n2 96.723
R148 a_79_21.n8 a_79_21.n7 76
R149 a_79_21.n5 a_79_21.n4 76
R150 a_79_21.n11 a_79_21.n10 76
R151 a_79_21.n15 a_79_21.n12 72.914
R152 a_79_21.n16 a_79_21.n15 48.575
R153 a_79_21.n17 a_79_21.n16 42.273
R154 a_79_21.n14 a_79_21.n13 42.273
R155 a_79_21.n2 a_79_21.n1 27.751
R156 a_79_21.n0 a_79_21.t2 26.595
R157 a_79_21.n0 a_79_21.t3 26.595
R158 a_79_21.n13 a_79_21.t7 24.923
R159 a_79_21.n13 a_79_21.t5 24.923
R160 a_79_21.n17 a_79_21.t4 24.923
R161 a_79_21.t1 a_79_21.n17 24.923
R162 a_79_21.n11 a_79_21.n8 20.723
R163 a_79_21.n8 a_79_21.n5 20.723
R164 a_79_21.n4 a_79_21.n3 16.066
R165 a_79_21.n15 a_79_21.n14 12.308
R166 a_79_21.n10 a_79_21.n9 7.303
R167 a_79_21.n7 a_79_21.n6 4.381
R168 VPWR.n2 VPWR.t0 557.771
R169 VPWR.n1 VPWR.n0 314.004
R170 VPWR.n16 VPWR.t2 200.801
R171 VPWR.n12 VPWR.n11 171.981
R172 VPWR.n6 VPWR.n5 171.981
R173 VPWR.n11 VPWR.t4 26.595
R174 VPWR.n11 VPWR.t3 26.595
R175 VPWR.n5 VPWR.t7 26.595
R176 VPWR.n5 VPWR.t5 26.595
R177 VPWR.n0 VPWR.t1 26.595
R178 VPWR.n0 VPWR.t6 26.595
R179 VPWR.n2 VPWR.n1 10.207
R180 VPWR.n4 VPWR.n3 4.65
R181 VPWR.n8 VPWR.n7 4.65
R182 VPWR.n10 VPWR.n9 4.65
R183 VPWR.n13 VPWR.n12 4.65
R184 VPWR.n15 VPWR.n14 4.65
R185 VPWR.n17 VPWR.n16 4.65
R186 VPWR.n4 VPWR.n2 0.463
R187 VPWR.n7 VPWR.n6 0.376
R188 VPWR.n8 VPWR.n4 0.119
R189 VPWR.n10 VPWR.n8 0.119
R190 VPWR.n13 VPWR.n10 0.119
R191 VPWR.n15 VPWR.n13 0.119
R192 VPWR.n17 VPWR.n15 0.119
R193 VPWR VPWR.n17 0.019
R194 C1.n0 C1.t0 213.734
R195 C1.n1 C1.t1 212.079
R196 C1.n1 C1.t2 141.372
R197 C1.n0 C1.t3 139.779
R198 C1 C1.n2 88.495
R199 C1.n2 C1.n0 35.054
R200 C1.n2 C1.n1 24.83
R201 X.n5 X.n3 155.183
R202 X.n5 X.n4 110.761
R203 X.n2 X.n0 88.89
R204 X.n2 X.n1 52.624
R205 X.n3 X.t3 26.595
R206 X.n3 X.t2 26.595
R207 X.n4 X.t1 26.595
R208 X.n4 X.t0 26.595
R209 X.n1 X.t7 24.923
R210 X.n1 X.t4 24.923
R211 X.n0 X.t6 24.923
R212 X.n0 X.t5 24.923
R213  X.n5 22.603
R214 X  18.921
R215 X.n6 X 15.86
R216 X.n6 X.n2 14.498
R217 X X.n6 3.06
C0 X VGND 0.43fF
C1 VPWR VGND 0.14fF
C2 VPWR VPB 0.15fF
C3 VPWR X 0.68fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__a221oi_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__a221oi_1 Y C1 A1 A2 B2 B1 VGND VPWR VNB VPB
X0 a_465_47.t1 A1.t0 Y.t1 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 a_109_297.t0 B1.t0 a_193_297.t2 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 a_193_297.t3 B2.t0 a_109_297.t2 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 a_204_47.t0 B2.t1 VGND.t1 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 VGND.t0 A2.t0 a_465_47.t0 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 a_193_297.t1 A1.t1 VPWR.t1 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 Y.t0 B1.t1 a_204_47.t1 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 VPWR.t0 A2.t1 a_193_297.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 a_109_297.t1 C1.t0 Y.t2 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 VGND.t2 C1.t1 Y.t3 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
R0 A1.n0 A1.t1 234.801
R1 A1.n0 A1.t0 162.501
R2 A1 A1.n0 78.76
R3 Y Y.t2 489.973
R4 Y.n0 Y.t3 233.312
R5 Y.n0 Y.t0 157.115
R6 Y.n1 Y.t1 157.115
R7 Y Y.n1 65.067
R8 Y.n1 Y.n0 26.624
R9 a_465_47.t0 a_465_47.t1 56.307
R10 VNB VNB.t4 6078.09
R11 VNB.t0 VNB.t2 4545.05
R12 VNB.t4 VNB.t3 2296.7
R13 VNB.t2 VNB.t1 2200
R14 VNB.t3 VNB.t0 1764.83
R15 B1.n0 B1.t0 239.038
R16 B1.n0 B1.t1 166.738
R17 B1 B1.n0 80.951
R18 a_193_297.n1 a_193_297.n0 512.302
R19 a_193_297.t0 a_193_297.n1 33.49
R20 a_193_297.n0 a_193_297.t2 26.595
R21 a_193_297.n0 a_193_297.t3 26.595
R22 a_193_297.n1 a_193_297.t1 26.595
R23 a_109_297.t0 a_109_297.n0 770.533
R24 a_109_297.n0 a_109_297.t2 26.595
R25 a_109_297.n0 a_109_297.t1 26.595
R26 VPB.t2 VPB.t1 556.386
R27 VPB.t1 VPB.t0 269.314
R28 VPB.t4 VPB.t2 248.598
R29 VPB.t3 VPB.t4 248.598
R30 VPB VPB.t3 192.367
R31 B2.n0 B2.t0 241.534
R32 B2.n0 B2.t1 169.234
R33 B2 B2.n0 92.761
R34 VGND.n1 VGND.t0 175.315
R35 VGND.n1 VGND.n0 112.984
R36 VGND.n0 VGND.t1 35.076
R37 VGND.n0 VGND.t2 24.923
R38 VGND VGND.n1 0.143
R39 a_204_47.t0 a_204_47.t1 39.692
R40 A2.n0 A2.t1 241.534
R41 A2.n0 A2.t0 169.234
R42 A2 A2.n0 83.757
R43 VPWR.n0 VPWR.t1 550.772
R44 VPWR.n0 VPWR.t0 205.231
R45 VPWR VPWR.n0 0.586
R46 C1.n0 C1.t0 230.154
R47 C1.n0 C1.t1 157.854
R48 C1 C1.n0 82.4
C0 A1 Y 0.17fF
C1 VGND Y 0.57fF
C2 B1 Y 0.21fF
C3 VPWR Y 0.11fF
C4 A2 Y 0.18fF
C5 B2 Y 0.20fF
C6 C1 Y 0.10fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__a221oi_2.ext - technology: sky130A

.subckt sky130_fd_sc_hd__a221oi_2 B2 C1 A2 A1 B1 Y VGND VPWR VNB VPB
X0 Y.t3 B1.t0 a_383_47.t3 VNB.t7 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 a_301_297.t7 B1.t1 a_27_297.t3 VPB.t7 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 a_301_297.t5 A2.t0 VPWR.t3 VPB.t5 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 VGND.t1 B2.t0 a_383_47.t1 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 Y.t0 A1.t0 a_735_47.t3 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 a_27_297.t1 B2.t1 a_301_297.t1 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 VPWR.t0 A1.t1 a_301_297.t3 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 VGND.t3 A2.t1 a_735_47.t1 VNB.t5 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 a_301_297.t4 A1.t2 VPWR.t1 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 Y.t4 C1.t0 a_27_297.t4 VPB.t8 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 VGND.t4 C1.t1 Y.t5 VNB.t8 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 Y.t6 C1.t2 VGND.t5 VNB.t9 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 VPWR.t2 A2.t2 a_301_297.t2 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13 a_383_47.t0 B2.t2 VGND.t0 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14 a_383_47.t2 B1.t2 Y.t2 VNB.t6 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X15 a_735_47.t0 A2.t3 VGND.t2 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X16 a_27_297.t5 C1.t3 Y.t7 VPB.t9 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17 a_301_297.t0 B2.t3 a_27_297.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X18 a_735_47.t2 A1.t3 Y.t1 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X19 a_27_297.t2 B1.t3 a_301_297.t6 VPB.t6 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
R0 B1.n0 B1.t3 212.079
R1 B1.n1 B1.t1 212.079
R2 B1.n0 B1.t2 139.779
R3 B1.n1 B1.t0 139.779
R4 B1 B1.n2 77.268
R5 B1.n2 B1.n0 30.672
R6 B1.n2 B1.n1 30.672
R7 a_383_47.n1 a_383_47.n0 233.872
R8 a_383_47.n0 a_383_47.t1 24.923
R9 a_383_47.n0 a_383_47.t2 24.923
R10 a_383_47.n1 a_383_47.t3 24.923
R11 a_383_47.t0 a_383_47.n1 24.923
R12 Y.n2 Y.n0 210.434
R13 Y.n4 Y.n3 146.375
R14 Y.n5 Y.n2 110.795
R15  Y.n6 94.292
R16 Y.n2 Y.n1 92.5
R17 Y.n7 Y.n6 92.5
R18 Y.n3 Y.t7 26.595
R19 Y.n3 Y.t4 26.595
R20 Y.n6 Y.t5 24.923
R21 Y.n6 Y.t6 24.923
R22 Y.n1 Y.t2 24.923
R23 Y.n1 Y.t3 24.923
R24 Y.n0 Y.t1 24.923
R25 Y.n0 Y.t0 24.923
R26 Y  17.408
R27 Y.n7  15.616
R28 Y.n5 Y 14.848
R29  Y.n4 13.062
R30 Y.n4  4.228
R31  Y.n5 2.56
R32  Y.n7 1.792
R33 VNB VNB.t9 6102.26
R34 VNB.t8 VNB.t0 4545.05
R35 VNB.t1 VNB.t2 2417.58
R36 VNB.t4 VNB.t5 2030.77
R37 VNB.t3 VNB.t4 2030.77
R38 VNB.t2 VNB.t3 2030.77
R39 VNB.t6 VNB.t1 2030.77
R40 VNB.t7 VNB.t6 2030.77
R41 VNB.t0 VNB.t7 2030.77
R42 VNB.t9 VNB.t8 2030.77
R43 a_27_297.n3 a_27_297.n2 346.333
R44 a_27_297.n2 a_27_297.n0 292.5
R45 a_27_297.n1 a_27_297.t5 264.699
R46 a_27_297.n1 a_27_297.t4 237.884
R47 a_27_297.n2 a_27_297.n1 64.618
R48 a_27_297.n0 a_27_297.t3 26.595
R49 a_27_297.n0 a_27_297.t1 26.595
R50 a_27_297.t0 a_27_297.n3 26.595
R51 a_27_297.n3 a_27_297.t2 26.595
R52 a_301_297.n4 a_301_297.t1 585.006
R53 a_301_297.n5 a_301_297.n4 292.5
R54 a_301_297.n1 a_301_297.t5 179.392
R55 a_301_297.n1 a_301_297.n0 155.085
R56 a_301_297.n3 a_301_297.n2 141.904
R57 a_301_297.n4 a_301_297.n3 64.93
R58 a_301_297.n3 a_301_297.n1 60.225
R59 a_301_297.n2 a_301_297.t2 34.475
R60 a_301_297.n2 a_301_297.t0 34.475
R61 a_301_297.n0 a_301_297.t3 26.595
R62 a_301_297.n0 a_301_297.t4 26.595
R63 a_301_297.t6 a_301_297.n5 26.595
R64 a_301_297.n5 a_301_297.t7 26.595
R65 VPB.t9 VPB.t1 556.386
R66 VPB.t0 VPB.t2 295.95
R67 VPB.t3 VPB.t5 248.598
R68 VPB.t4 VPB.t3 248.598
R69 VPB.t2 VPB.t4 248.598
R70 VPB.t6 VPB.t0 248.598
R71 VPB.t7 VPB.t6 248.598
R72 VPB.t1 VPB.t7 248.598
R73 VPB.t8 VPB.t9 248.598
R74 VPB VPB.t8 195.327
R75 A2.n0 A2.t0 241.534
R76 A2.n1 A2.t2 241.534
R77 A2.n2 A2.n1 184.186
R78 A2.n0 A2.t1 169.234
R79 A2.n1 A2.t3 169.234
R80 A2.n2 A2.n0 76
R81 A2 A2.n2 23.68
R82 VPWR.n2 VPWR.n0 319.467
R83 VPWR.n2 VPWR.n1 317.297
R84 VPWR.n0 VPWR.t3 26.595
R85 VPWR.n0 VPWR.t0 26.595
R86 VPWR.n1 VPWR.t1 26.595
R87 VPWR.n1 VPWR.t2 26.595
R88 VPWR VPWR.n2 1.116
R89 B2.n1 B2.t1 241.534
R90 B2.n0 B2.t3 241.534
R91 B2.n1 B2.t2 169.234
R92 B2.n0 B2.t0 169.234
R93 B2.n2 B2.n0 162.479
R94 B2.n2 B2.n1 76
R95 B2 B2.n2 6.874
R96 VGND.n2 VGND.t3 125.614
R97 VGND.n1 VGND.n0 115.464
R98 VGND.n19 VGND.t5 108.134
R99 VGND.n10 VGND.n9 92.5
R100 VGND.n14 VGND.n13 92.5
R101 VGND.n0 VGND.t1 33.23
R102 VGND.n0 VGND.t2 31.384
R103 VGND.n9 VGND.t0 24.923
R104 VGND.n13 VGND.t4 24.923
R105 VGND.n2 VGND.n1 11.289
R106 VGND.n20 VGND.n19 4.65
R107 VGND.n4 VGND.n3 4.65
R108 VGND.n6 VGND.n5 4.65
R109 VGND.n8 VGND.n7 4.65
R110 VGND.n12 VGND.n11 4.65
R111 VGND.n16 VGND.n15 4.65
R112 VGND.n18 VGND.n17 4.65
R113 VGND.n15 VGND.n14 0.8
R114 VGND.n11 VGND.n10 0.4
R115 VGND.n4 VGND.n2 0.137
R116 VGND.n6 VGND.n4 0.119
R117 VGND.n8 VGND.n6 0.119
R118 VGND.n12 VGND.n8 0.119
R119 VGND.n16 VGND.n12 0.119
R120 VGND.n18 VGND.n16 0.119
R121 VGND.n20 VGND.n18 0.119
R122 VGND VGND.n20 0.02
R123 A1.n0 A1.t1 212.079
R124 A1.n1 A1.t2 212.079
R125 A1.n0 A1.t3 139.779
R126 A1.n1 A1.t0 139.779
R127 A1 A1.n2 81.12
R128 A1.n2 A1.n0 30.672
R129 A1.n2 A1.n1 30.672
R130 a_735_47.n1 a_735_47.n0 187.935
R131 a_735_47.n0 a_735_47.t3 24.923
R132 a_735_47.n0 a_735_47.t0 24.923
R133 a_735_47.t1 a_735_47.n1 24.923
R134 a_735_47.n1 a_735_47.t2 24.923
R135 C1.n0 C1.t3 212.079
R136 C1.n1 C1.t0 212.079
R137 C1.n0 C1.t1 139.779
R138 C1.n1 C1.t2 139.779
R139 C1.n2 C1.n1 108.863
R140 C1.n1 C1.n0 61.345
R141 C1.n2 C1 11.054
R142 C1 C1.n2 2.133
C0 VPB VPWR 0.10fF
C1 B2 A2 0.14fF
C2 B2 B1 0.33fF
C3 VGND VPWR 0.12fF
C4 VGND Y 0.45fF
C5 Y B1 0.12fF
C6 A1 A2 0.31fF
C7 Y B2 0.20fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__a221oi_4.ext - technology: sky130A

.subckt sky130_fd_sc_hd__a221oi_4 A2 Y C1 A1 B2 B1 VPWR VGND VNB VPB
X0 Y.t3 A1.t0 a_1241_47.t4 VNB.t6 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 a_453_47.t7 B2.t0 VGND.t9 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 Y.t8 B1.t0 a_453_47.t0 VNB.t10 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 Y.t2 A1.t1 a_1241_47.t3 VNB.t5 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 Y.t10 C1.t0 a_27_297.t3 VPB.t9 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 a_471_297.t7 A2.t0 VPWR.t7 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 Y.t9 B1.t1 a_453_47.t1 VNB.t11 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 VGND.t1 A2.t1 a_1241_47.t5 VNB.t7 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 Y.t11 C1.t1 VGND.t4 VNB.t12 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 a_27_297.t2 C1.t2 Y.t12 VPB.t8 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 VPWR.t6 A2.t2 a_471_297.t6 VPB.t5 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 a_453_47.t2 B1.t2 Y.t14 VNB.t16 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 a_471_297.t15 B2.t1 a_27_297.t11 VPB.t17 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13 VGND.t8 B2.t2 a_453_47.t6 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14 a_1241_47.t2 A1.t2 Y.t1 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X15 a_27_297.t10 B2.t3 a_471_297.t14 VPB.t16 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16 a_453_47.t3 B1.t3 Y.t15 VNB.t17 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X17 a_1241_47.t1 A1.t3 Y.t0 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X18 VGND.t5 C1.t3 Y.t13 VNB.t13 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X19 a_1241_47.t6 A2.t3 VGND.t10 VNB.t18 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X20 Y.t4 C1.t4 VGND.t2 VNB.t8 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X21 VGND.t3 C1.t5 Y.t5 VNB.t9 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X22 VPWR.t5 A2.t4 a_471_297.t5 VPB.t18 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X23 a_471_297.t13 B2.t4 a_27_297.t9 VPB.t15 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X24 a_471_297.t4 A2.t5 VPWR.t4 VPB.t19 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X25 a_471_297.t11 B1.t4 a_27_297.t7 VPB.t13 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X26 VPWR.t3 A1.t4 a_471_297.t3 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X27 Y.t6 C1.t6 a_27_297.t1 VPB.t7 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X28 a_27_297.t6 B1.t5 a_471_297.t10 VPB.t12 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X29 VGND.t11 A2.t6 a_1241_47.t7 VNB.t19 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X30 a_471_297.t2 A1.t5 VPWR.t2 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X31 a_27_297.t5 B1.t6 a_471_297.t9 VPB.t11 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X32 a_1241_47.t0 A2.t7 VGND.t0 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X33 a_471_297.t8 B1.t7 a_27_297.t4 VPB.t10 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X34 VPWR.t1 A1.t6 a_471_297.t1 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X35 a_27_297.t8 B2.t5 a_471_297.t12 VPB.t14 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X36 a_471_297.t0 A1.t7 VPWR.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X37 a_27_297.t0 C1.t7 Y.t7 VPB.t6 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X38 a_453_47.t5 B2.t6 VGND.t7 VNB.t14 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X39 VGND.t6 B2.t7 a_453_47.t4 VNB.t15 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
R0 A1.n0 A1.t4 212.079
R1 A1.n2 A1.t5 212.079
R2 A1.n7 A1.t6 212.079
R3 A1.n5 A1.t7 212.079
R4 A1.n0 A1.t3 139.779
R5 A1.n2 A1.t1 139.779
R6 A1.n7 A1.t2 139.779
R7 A1.n5 A1.t0 139.779
R8 A1.n9 A1.n6 97.76
R9 A1.n4 A1.n1 97.76
R10 A1.n4 A1.n3 76
R11 A1.n9 A1.n8 76
R12 A1.n1 A1.n0 21.909
R13 A1 A1.n4 16
R14 A1.n6 A1.n5 13.145
R15 A1.n3 A1.n2 10.224
R16 A1 A1.n9 5.76
R17 A1.n8 A1.n7 1.46
R18 a_1241_47.n5 a_1241_47.n4 141.372
R19 a_1241_47.n2 a_1241_47.n0 101.198
R20 a_1241_47.n4 a_1241_47.n3 92.5
R21 a_1241_47.n4 a_1241_47.n2 53.163
R22 a_1241_47.n2 a_1241_47.n1 42.273
R23 a_1241_47.n3 a_1241_47.t3 24.923
R24 a_1241_47.n3 a_1241_47.t2 24.923
R25 a_1241_47.n1 a_1241_47.t5 24.923
R26 a_1241_47.n1 a_1241_47.t1 24.923
R27 a_1241_47.n0 a_1241_47.t7 24.923
R28 a_1241_47.n0 a_1241_47.t6 24.923
R29 a_1241_47.n5 a_1241_47.t4 24.923
R30 a_1241_47.t0 a_1241_47.n5 24.923
R31 Y.n9 Y.n8 208.919
R32 Y.n10 Y.n6 197.313
R33 Y.n2 Y.n0 153.94
R34 Y.n9 Y.n7 150.733
R35 Y.n4 Y.n2 121.911
R36 Y.n2 Y.n1 92.5
R37 Y.n6 Y.n5 92.5
R38 Y.n4 Y.n3 92.5
R39 Y.n13 Y.n11 88.89
R40 Y.n6 Y.n4 61.44
R41 Y.n13 Y.n12 52.624
R42 Y.n8 Y.t12 26.595
R43 Y.n8 Y.t6 26.595
R44 Y.n7 Y.t7 26.595
R45 Y.n7 Y.t10 26.595
R46 Y.n3 Y.t14 24.923
R47 Y.n3 Y.t9 24.923
R48 Y.n5 Y.t15 24.923
R49 Y.n5 Y.t8 24.923
R50 Y.n0 Y.t0 24.923
R51 Y.n0 Y.t2 24.923
R52 Y.n1 Y.t1 24.923
R53 Y.n1 Y.t3 24.923
R54 Y.n12 Y.t5 24.923
R55 Y.n12 Y.t11 24.923
R56 Y.n11 Y.t13 24.923
R57 Y.n11 Y.t4 24.923
R58 Y.n10 Y.n9 21.534
R59 Y Y.n13 16.29
R60 Y Y.n10 5.12
R61 VNB VNB.t8 6150.61
R62 VNB.t0 VNB.t10 4448.35
R63 VNB.t15 VNB.t2 2417.58
R64 VNB.t9 VNB.t14 2127.47
R65 VNB.t18 VNB.t19 2030.77
R66 VNB.t7 VNB.t18 2030.77
R67 VNB.t3 VNB.t7 2030.77
R68 VNB.t5 VNB.t3 2030.77
R69 VNB.t4 VNB.t5 2030.77
R70 VNB.t6 VNB.t4 2030.77
R71 VNB.t2 VNB.t6 2030.77
R72 VNB.t16 VNB.t15 2030.77
R73 VNB.t11 VNB.t16 2030.77
R74 VNB.t17 VNB.t11 2030.77
R75 VNB.t10 VNB.t17 2030.77
R76 VNB.t1 VNB.t0 2030.77
R77 VNB.t14 VNB.t1 2030.77
R78 VNB.t12 VNB.t9 2030.77
R79 VNB.t13 VNB.t12 2030.77
R80 VNB.t8 VNB.t13 2030.77
R81 B2.n0 B2.t4 241.534
R82 B2.n5 B2.t5 216.46
R83 B2.n4 B2.t1 212.079
R84 B2.n2 B2.t3 212.079
R85 B2 B2.n0 211.951
R86 B2.n1 B2.t6 201.124
R87 B2.n0 B2.t7 169.234
R88 B2.n1 B2.t2 139.779
R89 B2.n3 B2.t0 139.779
R90 B2 B2.n5 104.816
R91 B2.n5 B2.n4 56.963
R92 B2.n3 B2.n2 49.66
R93 B2.n4 B2.n3 11.684
R94 B2.n2 B2.n1 11.684
R95 VGND.n33 VGND.n31 151.014
R96 VGND.n2 VGND.t11 124.459
R97 VGND.n1 VGND.n0 115.464
R98 VGND.n14 VGND.n13 115.464
R99 VGND.n40 VGND.n39 115.464
R100 VGND.n45 VGND.t2 106.782
R101 VGND.n33 VGND.n32 92.5
R102 VGND.n13 VGND.t6 39.692
R103 VGND.n32 VGND.t7 28.615
R104 VGND.n0 VGND.t10 24.923
R105 VGND.n0 VGND.t1 24.923
R106 VGND.n13 VGND.t0 24.923
R107 VGND.n32 VGND.t3 24.923
R108 VGND.n31 VGND.t9 24.923
R109 VGND.n31 VGND.t8 24.923
R110 VGND.n39 VGND.t4 24.923
R111 VGND.n39 VGND.t5 24.923
R112 VGND.n34 VGND.n33 22.964
R113 VGND.n15 VGND.n14 12.8
R114 VGND.n2 VGND.n1 9.23
R115 VGND.n35 VGND.n34 8.282
R116 VGND.n46 VGND.n45 4.65
R117 VGND.n4 VGND.n3 4.65
R118 VGND.n6 VGND.n5 4.65
R119 VGND.n8 VGND.n7 4.65
R120 VGND.n10 VGND.n9 4.65
R121 VGND.n12 VGND.n11 4.65
R122 VGND.n16 VGND.n15 4.65
R123 VGND.n18 VGND.n17 4.65
R124 VGND.n20 VGND.n19 4.65
R125 VGND.n22 VGND.n21 4.65
R126 VGND.n24 VGND.n23 4.65
R127 VGND.n26 VGND.n25 4.65
R128 VGND.n28 VGND.n27 4.65
R129 VGND.n30 VGND.n29 4.65
R130 VGND.n36 VGND.n35 4.65
R131 VGND.n38 VGND.n37 4.65
R132 VGND.n42 VGND.n41 4.65
R133 VGND.n44 VGND.n43 4.65
R134 VGND.n41 VGND.n40 2.258
R135 VGND.n4 VGND.n2 0.313
R136 VGND.n6 VGND.n4 0.119
R137 VGND.n8 VGND.n6 0.119
R138 VGND.n10 VGND.n8 0.119
R139 VGND.n12 VGND.n10 0.119
R140 VGND.n16 VGND.n12 0.119
R141 VGND.n18 VGND.n16 0.119
R142 VGND.n20 VGND.n18 0.119
R143 VGND.n22 VGND.n20 0.119
R144 VGND.n24 VGND.n22 0.119
R145 VGND.n26 VGND.n24 0.119
R146 VGND.n28 VGND.n26 0.119
R147 VGND.n30 VGND.n28 0.119
R148 VGND.n36 VGND.n30 0.119
R149 VGND.n38 VGND.n36 0.119
R150 VGND.n42 VGND.n38 0.119
R151 VGND.n44 VGND.n42 0.119
R152 VGND.n46 VGND.n44 0.119
R153 VGND VGND.n46 0.02
R154 a_453_47.n7 a_453_47.n6 148.645
R155 a_453_47.n2 a_453_47.n0 141.372
R156 a_453_47.n2 a_453_47.n1 92.5
R157 a_453_47.n4 a_453_47.n3 92.5
R158 a_453_47.n6 a_453_47.n5 92.5
R159 a_453_47.n4 a_453_47.n2 48.872
R160 a_453_47.n6 a_453_47.n4 29.09
R161 a_453_47.n3 a_453_47.t0 24.923
R162 a_453_47.n5 a_453_47.t7 24.923
R163 a_453_47.n1 a_453_47.t1 24.923
R164 a_453_47.n1 a_453_47.t3 24.923
R165 a_453_47.n0 a_453_47.t4 24.923
R166 a_453_47.n0 a_453_47.t2 24.923
R167 a_453_47.t6 a_453_47.n7 24.923
R168 a_453_47.n7 a_453_47.t5 24.923
R169 B1.n0 B1.t5 212.079
R170 B1.n2 B1.t4 212.079
R171 B1.n5 B1.t6 212.079
R172 B1.n8 B1.t7 212.079
R173 B1.n0 B1.t2 139.779
R174 B1.n2 B1.t1 139.779
R175 B1.n5 B1.t3 139.779
R176 B1.n8 B1.t0 139.779
R177 B1.n4 B1.n1 91.542
R178 B1 B1.n9 85.6
R179 B1.n4 B1.n3 76
R180 B1.n7 B1.n6 76
R181 B1.n9 B1.n8 21.909
R182 B1.n7 B1.n4 15.542
R183 B1.n1 B1.n0 13.145
R184 B1.n6 B1.n5 10.224
R185 B1 B1.n7 5.942
R186 B1.n3 B1.n2 1.46
R187 C1.n3 C1.t6 212.079
R188 C1.n0 C1.t7 212.079
R189 C1.n1 C1.t0 212.079
R190 C1.n4 C1.t2 212.079
R191 C1.n3 C1.t4 139.779
R192 C1.n0 C1.t5 139.779
R193 C1.n1 C1.t1 139.779
R194 C1.n4 C1.t3 139.779
R195 C1 C1.n2 82.4
R196 C1.n1 C1.n0 61.345
R197 C1 C1.n5 48.615
R198 C1.n5 C1.n4 28.577
R199 C1.n2 C1.n1 23.369
R200 C1.n5 C1.n3 21.73
R201 a_27_297.n2 a_27_297.n0 343.7
R202 a_27_297.n2 a_27_297.n1 292.5
R203 a_27_297.n4 a_27_297.n3 292.5
R204 a_27_297.n8 a_27_297.t1 179.121
R205 a_27_297.n9 a_27_297.n8 154.572
R206 a_27_297.n6 a_27_297.n5 143.076
R207 a_27_297.n7 a_27_297.t0 116.829
R208 a_27_297.n7 a_27_297.n6 78.157
R209 a_27_297.n8 a_27_297.n7 67.45
R210 a_27_297.n4 a_27_297.n2 51.2
R211 a_27_297.n6 a_27_297.n4 50.068
R212 a_27_297.n5 a_27_297.t11 26.595
R213 a_27_297.n5 a_27_297.t10 26.595
R214 a_27_297.n3 a_27_297.t4 26.595
R215 a_27_297.n3 a_27_297.t8 26.595
R216 a_27_297.n1 a_27_297.t7 26.595
R217 a_27_297.n1 a_27_297.t5 26.595
R218 a_27_297.n0 a_27_297.t9 26.595
R219 a_27_297.n0 a_27_297.t6 26.595
R220 a_27_297.t3 a_27_297.n9 26.595
R221 a_27_297.n9 a_27_297.t2 26.595
R222 VPB.t6 VPB.t16 556.386
R223 VPB.t15 VPB.t5 295.95
R224 VPB.t18 VPB.t4 248.598
R225 VPB.t19 VPB.t18 248.598
R226 VPB.t3 VPB.t19 248.598
R227 VPB.t2 VPB.t3 248.598
R228 VPB.t1 VPB.t2 248.598
R229 VPB.t0 VPB.t1 248.598
R230 VPB.t5 VPB.t0 248.598
R231 VPB.t12 VPB.t15 248.598
R232 VPB.t13 VPB.t12 248.598
R233 VPB.t11 VPB.t13 248.598
R234 VPB.t10 VPB.t11 248.598
R235 VPB.t14 VPB.t10 248.598
R236 VPB.t17 VPB.t14 248.598
R237 VPB.t16 VPB.t17 248.598
R238 VPB.t9 VPB.t6 248.598
R239 VPB.t8 VPB.t9 248.598
R240 VPB.t7 VPB.t8 248.598
R241 VPB VPB.t7 201.246
R242 A2.n6 A2.n5 254.04
R243 A2.n5 A2.t2 241.534
R244 A2.n0 A2.t0 212.079
R245 A2.n1 A2.t4 212.079
R246 A2.n3 A2.t5 212.079
R247 A2.n5 A2.t7 169.234
R248 A2.n0 A2.t6 139.779
R249 A2.n1 A2.t3 139.779
R250 A2.n3 A2.t1 139.779
R251 A2.n6 A2.n4 76
R252 A2 A2.n2 46.695
R253 A2.n2 A2.n0 31.954
R254 A2.n2 A2.n1 18.353
R255 A2.n4 A2.n3 13.145
R256 A2 A2.n6 8.32
R257 VPWR.n4 VPWR.n3 292.5
R258 VPWR.n9 VPWR.n8 292.5
R259 VPWR.n1 VPWR.n0 292.5
R260 VPWR.n5 VPWR.n2 186.42
R261 VPWR.n0 VPWR.t0 26.595
R262 VPWR.n0 VPWR.t6 26.595
R263 VPWR.n8 VPWR.t2 26.595
R264 VPWR.n8 VPWR.t1 26.595
R265 VPWR.n3 VPWR.t4 26.595
R266 VPWR.n3 VPWR.t3 26.595
R267 VPWR.n2 VPWR.t7 26.595
R268 VPWR.n2 VPWR.t5 26.595
R269 VPWR.n14 VPWR.n1 6.937
R270 VPWR.n7 VPWR.n6 4.65
R271 VPWR.n11 VPWR.n10 4.65
R272 VPWR.n13 VPWR.n12 4.65
R273 VPWR.n5 VPWR.n4 4.518
R274 VPWR VPWR.n14 1.559
R275 VPWR.n10 VPWR.n9 1.084
R276 VPWR.n7 VPWR.n5 0.306
R277 VPWR.n14 VPWR.n13 0.134
R278 VPWR.n11 VPWR.n7 0.119
R279 VPWR.n13 VPWR.n11 0.119
R280 a_471_297.n9 a_471_297.n4 292.5
R281 a_471_297.n8 a_471_297.n5 292.5
R282 a_471_297.n7 a_471_297.n6 292.5
R283 a_471_297.n11 a_471_297.n2 292.5
R284 a_471_297.n13 a_471_297.n12 292.5
R285 a_471_297.n7 a_471_297.t14 219.535
R286 a_471_297.n1 a_471_297.t7 202.417
R287 a_471_297.n1 a_471_297.n0 150.897
R288 a_471_297.n10 a_471_297.n3 144.107
R289 a_471_297.n10 a_471_297.n9 49.345
R290 a_471_297.n11 a_471_297.n10 47.612
R291 a_471_297.n9 a_471_297.n8 43.008
R292 a_471_297.n8 a_471_297.n7 43.008
R293 a_471_297.n12 a_471_297.n1 41.353
R294 a_471_297.n12 a_471_297.n11 41.353
R295 a_471_297.n3 a_471_297.t6 34.475
R296 a_471_297.n3 a_471_297.t13 34.475
R297 a_471_297.n6 a_471_297.t12 26.595
R298 a_471_297.n6 a_471_297.t15 26.595
R299 a_471_297.n5 a_471_297.t9 26.595
R300 a_471_297.n5 a_471_297.t8 26.595
R301 a_471_297.n4 a_471_297.t10 26.595
R302 a_471_297.n4 a_471_297.t11 26.595
R303 a_471_297.n2 a_471_297.t1 26.595
R304 a_471_297.n2 a_471_297.t0 26.595
R305 a_471_297.n0 a_471_297.t5 26.595
R306 a_471_297.n0 a_471_297.t4 26.595
R307 a_471_297.t3 a_471_297.n13 26.595
R308 a_471_297.n13 a_471_297.t2 26.595
C0 A1 Y 0.15fF
C1 A1 A2 0.54fF
C2 Y B1 0.34fF
C3 Y B2 0.23fF
C4 VPWR VPB 0.17fF
C5 Y C1 0.33fF
C6 B2 A2 0.14fF
C7 B2 B1 0.53fF
C8 VPWR VGND 0.20fF
C9 Y VGND 0.85fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__a222oi_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__a222oi_1 VPWR VGND C2 C1 B1 A2 A1 Y B2 VNB VPB
X0 Y.t1 B1.t0 a_393_47.t0 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1 VGND.t1 A2.t0 a_561_47.t0 VNB sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X2 VGND.t2 C2.t0 a_109_47.t1 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X3 Y.t2 C2.t1 a_109_297.t3 VPB.t5 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 VPWR.t0 A1.t0 a_311_297.t2 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 a_311_297.t3 A2.t1 VPWR.t1 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 a_311_297.t0 B1.t1 a_109_297.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 a_109_297.t2 B2.t0 a_311_297.t1 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 a_109_297.t1 C1.t0 Y.t3 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 a_393_47.t1 B2.t1 VGND.t0 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X10 a_109_47.t0 C1.t1 Y.t0 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X11 a_561_47.t1 A1.t1 Y.t4 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
R0 B1.n0 B1.t1 239.927
R1 B1.n0 B1.t0 172.447
R2 B1 B1.n0 79.296
R3 a_393_47.t0 a_393_47.t1 39.375
R4 Y.n0 Y.t2 534.961
R5 Y.n0 Y.t3 193.045
R6 Y.n2 Y.t0 151.436
R7 Y.n2 Y.n1 112.283
R8 Y Y.n0 44.523
R9 Y.n1 Y.t4 32.812
R10 Y.n1 Y.t1 29.062
R11 Y Y.n2 20.48
R12 VNB.n0 VNB 105600
R13 VNB.t4 VNB.t2 4640.8
R14 VNB.t1 VNB.t3 2101.49
R15 VNB.t3 VNB 2101.49
R16 VNB.n0 VNB.t0 2035.82
R17 VNB.t2 VNB.t1 1576.12
R18 VNB.t0 VNB.t4 1576.12
R19 VNB VNB.n0 21.89
R20 A2.n0 A2.t1 239.927
R21 A2.n0 A2.t0 172.447
R22 A2 A2.n0 79.576
R23 a_561_47.t0 a_561_47.t1 61.875
R24 VGND.n2 VGND.t1 107.787
R25 VGND.n1 VGND.n0 92.5
R26 VGND.n4 VGND.n3 92.5
R27 VGND.n0 VGND.t0 81.562
R28 VGND.n3 VGND.t2 25.312
R29 VGND.n2 VGND.n1 9.751
R30 VGND.n6 VGND.n5 4.65
R31 VGND.n5 VGND.n4 2.56
R32 VGND VGND.n7 0.166
R33 VGND.n6 VGND.n2 0.135
R34 VGND.n7 VGND.n6 0.132
R35 C2.n0 C2.t1 239.927
R36 C2.n0 C2.t0 172.447
R37 C2 C2.n0 78.594
R38 a_109_47.t0 a_109_47.t1 39.375
R39 a_109_297.n1 a_109_297.n0 550.741
R40 a_109_297.n0 a_109_297.t3 26.595
R41 a_109_297.n0 a_109_297.t1 26.595
R42 a_109_297.t0 a_109_297.n1 26.595
R43 a_109_297.n1 a_109_297.t2 26.595
R44 VPB.t5 VPB.t3 591.9
R45 VPB.t1 VPB.t4 284.112
R46 VPB VPB.t2 278.193
R47 VPB.t0 VPB.t1 248.598
R48 VPB.t3 VPB.t0 248.598
R49 VPB.t2 VPB.t5 248.598
R50 A1.n0 A1.t0 239.927
R51 A1.n0 A1.t1 172.447
R52 A1 A1.n0 79.296
R53 a_311_297.n0 a_311_297.t1 411.116
R54 a_311_297.n0 a_311_297.t3 190.391
R55 a_311_297.n1 a_311_297.n0 103.867
R56 a_311_297.n1 a_311_297.t2 26.595
R57 a_311_297.t0 a_311_297.n1 26.595
R58 VPWR VPWR.n0 181.246
R59 VPWR.n0 VPWR.t1 38.415
R60 VPWR.n0 VPWR.t0 26.595
R61 B2.n0 B2.t0 236.126
R62 B2.n0 B2.t1 168.646
R63 B2 B2.n0 79.096
R64 C1.n0 C1.t0 228.547
R65 C1.n0 C1.t1 161.067
R66 C1 C1.n0 85.142
C0 C1 C2 0.12fF
C1 Y VGND 0.34fF
C2 B1 B2 0.12fF
C3 Y B2 0.13fF
C4 Y C2 0.21fF
C5 Y C1 0.18fF
C6 A1 A2 0.11fF
C7 B1 A1 0.11fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__a311o_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__a311o_1 A1 A2 X B1 C1 A3 VGND VPWR VNB VPB
X0 a_75_199.t3 C1.t0 VGND.t3 VNB.t5 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 a_208_47.t0 A3.t0 VGND.t1 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 a_315_47.t1 A2.t0 a_208_47.t1 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 VGND.t2 B1.t0 a_75_199.t0 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 a_75_199.t1 A1.t0 a_315_47.t0 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 a_75_199.t2 C1.t1 a_544_297.t1 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 a_544_297.t0 B1.t1 a_201_297.t1 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 VPWR.t0 a_75_199.t4 X.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 a_201_297.t0 A3.t1 VPWR.t1 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 VPWR.t3 A2.t1 a_201_297.t3 VPB.t5 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 a_201_297.t2 A1.t1 VPWR.t2 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 VGND.t0 a_75_199.t5 X.t1 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
R0 C1.n0 C1.t1 230.361
R1 C1.n0 C1.t0 158.061
R2 C1 C1.n0 78.909
R3 VGND.n2 VGND.n0 111.984
R4 VGND.n2 VGND.n1 110.622
R5 VGND.n0 VGND.t2 38.769
R6 VGND.n1 VGND.t0 38.769
R7 VGND.n0 VGND.t3 37.846
R8 VGND.n1 VGND.t1 24.923
R9 VGND VGND.n2 0.15
R10 a_75_199.t2 a_75_199.n3 429.366
R11 a_75_199.n2 a_75_199.t3 268.173
R12 a_75_199.n0 a_75_199.t4 241.534
R13 a_75_199.n3 a_75_199.n2 169.446
R14 a_75_199.n0 a_75_199.t5 169.234
R15 a_75_199.n2 a_75_199.n1 92.5
R16 a_75_199.n3 a_75_199.n0 76
R17 a_75_199.n1 a_75_199.t1 30.461
R18 a_75_199.n1 a_75_199.t0 29.538
R19 VNB VNB.t0 6078.09
R20 VNB.t3 VNB.t4 3239.56
R21 VNB.t2 VNB.t5 2731.87
R22 VNB.t1 VNB.t3 2586.81
R23 VNB.t0 VNB.t1 2393.41
R24 VNB.t4 VNB.t2 2296.7
R25 A3.n0 A3.t1 241.534
R26 A3.n0 A3.t0 169.234
R27 A3 A3.n0 78.909
R28 a_208_47.t0 a_208_47.t1 71.076
R29 A2.n0 A2.t1 231.014
R30 A2.n0 A2.t0 158.714
R31 A2 A2.n0 79.61
R32 a_315_47.t0 a_315_47.t1 96
R33 B1.n0 B1.t1 241.534
R34 B1.n0 B1.t0 169.234
R35 B1 B1.n0 83.757
R36 A1.n0 A1.t1 241.534
R37 A1.n0 A1.t0 169.234
R38 A1.n1 A1.n0 82.4
R39 A1.n1 A1 15.494
R40 A1 A1.n1 2.909
R41 a_544_297.t0 a_544_297.t1 81.755
R42 VPB.t5 VPB.t4 449.844
R43 VPB.t2 VPB.t3 334.423
R44 VPB.t1 VPB.t5 284.112
R45 VPB.t4 VPB.t2 281.152
R46 VPB.t0 VPB.t1 257.476
R47 VPB VPB.t0 207.165
R48 a_201_297.n1 a_201_297.n0 381.728
R49 a_201_297.t0 a_201_297.n1 34.475
R50 a_201_297.n0 a_201_297.t2 32.505
R51 a_201_297.n0 a_201_297.t1 31.52
R52 a_201_297.n1 a_201_297.t3 30.535
R53 X X.t1 251.389
R54 X.n0 X.t0 178.6
R55 X X.n0 10.397
R56 X.n0 X 2.366
R57 VPWR.n9 VPWR.n8 312.353
R58 VPWR.n3 VPWR.n2 292.5
R59 VPWR.n1 VPWR.n0 292.5
R60 VPWR.n8 VPWR.t1 29.55
R61 VPWR.n0 VPWR.t2 26.595
R62 VPWR.n2 VPWR.t3 26.595
R63 VPWR.n8 VPWR.t0 26.595
R64 VPWR.n5 VPWR.n1 6.798
R65 VPWR.n5 VPWR.n4 4.65
R66 VPWR.n7 VPWR.n6 4.65
R67 VPWR.n10 VPWR.n9 4.05
R68 VPWR.n4 VPWR.n3 0.232
R69 VPWR.n10 VPWR.n7 0.134
R70 VPWR VPWR.n10 0.126
R71 VPWR.n7 VPWR.n5 0.119
.ends

* NGSPICE file created from sky130_fd_sc_hd__a311o_2.ext - technology: sky130A

.subckt sky130_fd_sc_hd__a311o_2 VGND VPWR X C1 B1 A1 A2 A3 VNB VPB
X0 a_79_21.t0 C1.t0 a_635_297.t1 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 VPWR.t1 A2.t0 a_319_297.t2 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 VGND.t2 B1.t0 a_79_21.t2 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 a_417_47.t0 A2.t1 a_319_47.t1 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 a_79_21.t3 A1.t0 a_417_47.t1 VNB.t6 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 a_319_47.t0 A3.t0 VGND.t0 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 VPWR.t3 a_79_21.t4 X.t3 VPB.t5 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 a_319_297.t3 A1.t1 VPWR.t4 VPB.t6 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 VGND.t4 a_79_21.t5 X.t1 VNB.t5 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 a_319_297.t0 A3.t1 VPWR.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 a_79_21.t1 C1.t1 VGND.t1 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 a_635_297.t0 B1.t1 a_319_297.t1 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 X.t2 a_79_21.t6 VPWR.t2 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13 X.t0 a_79_21.t7 VGND.t3 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
R0 C1.n0 C1.t0 236.932
R1 C1.n0 C1.t1 164.632
R2 C1 C1.n0 78.27
R3 a_635_297.t0 a_635_297.t1 82.74
R4 a_79_21.t0 a_79_21.n4 435.729
R5 a_79_21.n3 a_79_21.t1 256.879
R6 a_79_21.n1 a_79_21.t4 212.079
R7 a_79_21.n0 a_79_21.t6 212.079
R8 a_79_21.n4 a_79_21.n3 187.104
R9 a_79_21.n1 a_79_21.t5 139.779
R10 a_79_21.n0 a_79_21.t7 139.779
R11 a_79_21.n4 a_79_21.n1 106.672
R12 a_79_21.n3 a_79_21.n2 92.5
R13 a_79_21.n1 a_79_21.n0 61.345
R14 a_79_21.n2 a_79_21.t3 49.846
R15 a_79_21.n2 a_79_21.t2 25.846
R16 VPB.t5 VPB.t0 372.897
R17 VPB.t1 VPB.t2 337.383
R18 VPB.t6 VPB.t1 337.383
R19 VPB.t3 VPB.t6 307.788
R20 VPB.t0 VPB.t3 290.031
R21 VPB.t4 VPB.t5 248.598
R22 VPB VPB.t4 189.408
R23 A2.n0 A2.t0 241.534
R24 A2.n0 A2.t1 169.234
R25 A2 A2.n0 77.422
R26 a_319_297.n1 a_319_297.n0 366.911
R27 a_319_297.n0 a_319_297.t3 50.235
R28 a_319_297.n1 a_319_297.t2 35.46
R29 a_319_297.n0 a_319_297.t1 32.505
R30 a_319_297.t0 a_319_297.n1 31.52
R31 VPWR.n1 VPWR.n0 311.585
R32 VPWR.n3 VPWR.n2 173.143
R33 VPWR.n8 VPWR.t2 152.162
R34 VPWR.n2 VPWR.t3 55.16
R35 VPWR.n0 VPWR.t1 40.385
R36 VPWR.n2 VPWR.t0 39.4
R37 VPWR.n0 VPWR.t4 32.505
R38 VPWR.n5 VPWR.n4 4.65
R39 VPWR.n7 VPWR.n6 4.65
R40 VPWR.n9 VPWR.n8 4.65
R41 VPWR.n4 VPWR.n3 0.752
R42 VPWR.n5 VPWR.n1 0.4
R43 VPWR.n7 VPWR.n5 0.119
R44 VPWR.n9 VPWR.n7 0.119
R45 VPWR VPWR.n9 0.02
R46 B1.n0 B1.t1 241.534
R47 B1.n0 B1.t0 169.234
R48 B1 B1.n0 85.309
R49 VGND.n3 VGND.n0 111.965
R50 VGND.n6 VGND.t3 108.779
R51 VGND.n2 VGND.n1 107.239
R52 VGND.n1 VGND.t0 48.923
R53 VGND.n0 VGND.t2 40.615
R54 VGND.n1 VGND.t4 39.692
R55 VGND.n0 VGND.t1 38.769
R56 VGND.n7 VGND.n6 4.65
R57 VGND.n5 VGND.n4 4.65
R58 VGND.n3 VGND.n2 3.88
R59 VGND.n5 VGND.n3 0.141
R60 VGND.n7 VGND.n5 0.119
R61 VGND VGND.n7 0.02
R62 VNB VNB.t4 6053.91
R63 VNB.t5 VNB.t0 3046.15
R64 VNB.t3 VNB.t1 2804.4
R65 VNB.t6 VNB.t3 2707.69
R66 VNB.t2 VNB.t6 2514.28
R67 VNB.t0 VNB.t2 2369.23
R68 VNB.t4 VNB.t5 2030.77
R69 a_319_47.t0 a_319_47.t1 62.769
R70 a_417_47.t0 a_417_47.t1 68.307
R71 A1.n0 A1.t1 241.534
R72 A1.n0 A1.t0 169.234
R73 A1 A1.n0 78.995
R74 A3.n0 A3.t1 241.534
R75 A3.n0 A3.t0 169.234
R76 A3 A3.n0 79.274
R77 X.n1 X.n0 147.104
R78 X X.n2 94.245
R79 X.n3 X.n2 92.5
R80 X.n0 X.t3 26.595
R81 X.n0 X.t2 26.595
R82 X.n2 X.t1 24.923
R83 X.n2 X.t0 24.923
R84 X.n3 X 11.442
R85 X X.n1 10.71
R86 X.n4 X 8.339
R87 X X.n4 4.848
R88 X.n1 X 2.439
R89 X X.n3 1.745
C0 X VGND 0.18fF
C1 VPWR VGND 0.11fF
C2 VPWR X 0.26fF
C3 A2 A1 0.12fF
C4 A2 A3 0.10fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__a311o_4.ext - technology: sky130A

.subckt sky130_fd_sc_hd__a311o_4 VGND VPWR C1 A1 A2 A3 X B1 VNB VPB
X0 VPWR.t7 a_109_47.t8 X.t7 VPB.t8 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_277_297.t7 A1.t0 VPWR.t9 VPB.t11 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 X.t6 a_109_47.t9 VPWR.t6 VPB.t7 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 a_861_47.t3 A3.t0 VGND.t8 VNB.t10 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 a_27_297.t2 B1.t0 a_277_297.t4 VPB.t12 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 a_1059_47.t1 A2.t0 a_861_47.t0 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 a_1059_47.t3 A1.t1 a_109_47.t4 VNB.t13 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 a_277_297.t5 B1.t1 a_27_297.t1 VPB.t13 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 VGND.t5 a_109_47.t10 X.t5 VNB.t7 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 a_27_297.t3 C1.t0 a_109_47.t3 VPB.t9 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 VGND.t4 a_109_47.t11 X.t4 VNB.t6 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 VGND.t7 A3.t1 a_861_47.t2 VNB.t9 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 VGND.t0 C1.t1 a_109_47.t0 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 VGND.t9 B1.t2 a_109_47.t7 VNB.t11 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14 VPWR.t5 a_109_47.t12 X.t1 VPB.t6 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 a_109_47.t5 A1.t2 a_1059_47.t2 VNB.t12 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X16 X.t0 a_109_47.t13 VPWR.t4 VPB.t5 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17 X.t3 a_109_47.t14 VGND.t3 VNB.t5 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X18 a_109_47.t6 B1.t3 VGND.t6 VNB.t8 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X19 X.t2 a_109_47.t15 VGND.t2 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X20 VPWR.t0 A3.t2 a_277_297.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X21 VPWR.t2 A2.t1 a_277_297.t2 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X22 a_109_47.t1 C1.t2 a_27_297.t0 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X23 VPWR.t8 A1.t3 a_277_297.t6 VPB.t10 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X24 a_277_297.t1 A3.t3 VPWR.t1 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X25 a_277_297.t3 A2.t2 VPWR.t3 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X26 a_109_47.t2 C1.t3 VGND.t1 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X27 a_861_47.t1 A2.t3 a_1059_47.t0 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
R0 a_109_47.n3 a_109_47.n2 371.37
R1 a_109_47.n6 a_109_47.t12 221.719
R2 a_109_47.n8 a_109_47.t13 221.719
R3 a_109_47.n15 a_109_47.n14 213.032
R4 a_109_47.n0 a_109_47.t8 204.171
R5 a_109_47.n1 a_109_47.t9 191.624
R6 a_109_47.n10 a_109_47.t15 174.741
R7 a_109_47.n5 a_109_47.t11 147.989
R8 a_109_47.n9 a_109_47.t10 139.779
R9 a_109_47.n7 a_109_47.t14 139.779
R10 a_109_47.n4 a_109_47.n3 101.6
R11 a_109_47.n12 a_109_47.n10 96.256
R12 a_109_47.n14 a_109_47.n12 63.247
R13 a_109_47.n8 a_109_47.n7 54.626
R14 a_109_47.n14 a_109_47.n13 51.189
R15 a_109_47.n12 a_109_47.n11 51.189
R16 a_109_47.n6 a_109_47.n5 50.182
R17 a_109_47.n4 a_109_47.n1 42.17
R18 a_109_47.n10 a_109_47.n9 35.121
R19 a_109_47.n1 a_109_47.n0 29.993
R20 a_109_47.n15 a_109_47.t3 26.595
R21 a_109_47.t1 a_109_47.n15 26.595
R22 a_109_47.n11 a_109_47.t7 24.923
R23 a_109_47.n11 a_109_47.t6 24.923
R24 a_109_47.n13 a_109_47.t0 24.923
R25 a_109_47.n13 a_109_47.t2 24.923
R26 a_109_47.n2 a_109_47.t4 24.923
R27 a_109_47.n2 a_109_47.t5 24.923
R28 a_109_47.n5 a_109_47.n4 15.348
R29 a_109_47.n7 a_109_47.n6 12.853
R30 a_109_47.n9 a_109_47.n8 12.853
R31 X.n4 X.n3 338.805
R32 X.n4 X.n2 294.758
R33 X.n5 X.n0 91.057
R34 X.n5 X.n1 59.847
R35 X.n5 X 42.338
R36 X.n0 X.t2 28.615
R37 X.n3 X.t7 26.595
R38 X.n3 X.t6 26.595
R39 X.n2 X.t1 26.595
R40 X.n2 X.t0 26.595
R41 X.n1 X.t4 24.923
R42 X.n1 X.t3 24.923
R43 X.n0 X.t5 24.923
R44 X X.n4 12.143
R45 X X.n5 2.297
R46 VPWR.n19 VPWR.t4 576.219
R47 VPWR.n1 VPWR.n0 307.239
R48 VPWR.n11 VPWR.n10 307.239
R49 VPWR.n15 VPWR.n14 307.239
R50 VPWR.n6 VPWR.n5 306.011
R51 VPWR.n2 VPWR.t8 195.802
R52 VPWR.n0 VPWR.t9 101.455
R53 VPWR.n5 VPWR.t3 38.415
R54 VPWR.n0 VPWR.t2 26.595
R55 VPWR.n5 VPWR.t0 26.595
R56 VPWR.n10 VPWR.t1 26.595
R57 VPWR.n10 VPWR.t7 26.595
R58 VPWR.n14 VPWR.t6 26.595
R59 VPWR.n14 VPWR.t5 26.595
R60 VPWR.n12 VPWR.n11 4.894
R61 VPWR.n4 VPWR.n3 4.65
R62 VPWR.n7 VPWR.n6 4.65
R63 VPWR.n9 VPWR.n8 4.65
R64 VPWR.n13 VPWR.n12 4.65
R65 VPWR.n16 VPWR.n15 4.65
R66 VPWR.n18 VPWR.n17 4.65
R67 VPWR.n20 VPWR.n19 3.79
R68 VPWR.n2 VPWR.n1 3.591
R69 VPWR VPWR.n20 0.593
R70 VPWR.n4 VPWR.n2 0.166
R71 VPWR.n20 VPWR.n18 0.144
R72 VPWR.n7 VPWR.n4 0.119
R73 VPWR.n9 VPWR.n7 0.119
R74 VPWR.n13 VPWR.n9 0.119
R75 VPWR.n16 VPWR.n13 0.119
R76 VPWR.n18 VPWR.n16 0.119
R77 VPB.t12 VPB.t5 556.386
R78 VPB.t3 VPB.t11 473.52
R79 VPB.t0 VPB.t4 284.112
R80 VPB.t11 VPB.t10 248.598
R81 VPB.t4 VPB.t3 248.598
R82 VPB.t1 VPB.t0 248.598
R83 VPB.t8 VPB.t1 248.598
R84 VPB.t7 VPB.t8 248.598
R85 VPB.t6 VPB.t7 248.598
R86 VPB.t5 VPB.t6 248.598
R87 VPB.t13 VPB.t12 248.598
R88 VPB.t9 VPB.t13 248.598
R89 VPB.t2 VPB.t9 248.598
R90 VPB VPB.t2 189.408
R91 A1.n1 A1.t3 212.079
R92 A1.n0 A1.t0 212.079
R93 A1.n1 A1.t1 139.779
R94 A1.n0 A1.t2 139.779
R95 A1.n2 A1.n1 108.133
R96 A1.n1 A1.n0 61.345
R97  A1.n2 11.054
R98 A1.n2 A1 2.133
R99 a_277_297.n3 a_277_297.n2 563.299
R100 a_277_297.n5 a_277_297.n4 242.048
R101 a_277_297.n4 a_277_297.n0 150.188
R102 a_277_297.n3 a_277_297.n1 150.188
R103 a_277_297.n4 a_277_297.n3 67.764
R104 a_277_297.n1 a_277_297.t0 26.595
R105 a_277_297.n1 a_277_297.t1 26.595
R106 a_277_297.n0 a_277_297.t2 26.595
R107 a_277_297.n0 a_277_297.t3 26.595
R108 a_277_297.n2 a_277_297.t4 26.595
R109 a_277_297.n2 a_277_297.t5 26.595
R110 a_277_297.t6 a_277_297.n5 26.595
R111 a_277_297.n5 a_277_297.t7 26.595
R112 A3.n2 A3.t2 194.406
R113 A3.n0 A3.t3 184.766
R114 A3.n0 A3.t0 149.517
R115 A3.n1 A3.t1 128.533
R116 A3 A3.n2 81.485
R117 A3.n1 A3.n0 32.133
R118 A3.n2 A3.n1 3.213
R119 VGND.n0 VGND.t7 202.917
R120 VGND.n27 VGND.t1 186.826
R121 VGND.n10 VGND.n9 114.711
R122 VGND.n16 VGND.n15 114.711
R123 VGND.n22 VGND.n21 114.711
R124 VGND.n2 VGND.n1 92.5
R125 VGND.n4 VGND.n3 92.5
R126 VGND.n1 VGND.t8 32.307
R127 VGND.n3 VGND.t4 24.923
R128 VGND.n9 VGND.t3 24.923
R129 VGND.n9 VGND.t5 24.923
R130 VGND.n15 VGND.t2 24.923
R131 VGND.n15 VGND.t9 24.923
R132 VGND.n21 VGND.t6 24.923
R133 VGND.n21 VGND.t0 24.923
R134 VGND.n11 VGND.n10 14.305
R135 VGND.n17 VGND.n16 9.788
R136 VGND.n5 VGND.n4 5.485
R137 VGND.n28 VGND.n27 4.65
R138 VGND.n6 VGND.n5 4.65
R139 VGND.n8 VGND.n7 4.65
R140 VGND.n12 VGND.n11 4.65
R141 VGND.n14 VGND.n13 4.65
R142 VGND.n18 VGND.n17 4.65
R143 VGND.n20 VGND.n19 4.65
R144 VGND.n24 VGND.n23 4.65
R145 VGND.n26 VGND.n25 4.65
R146 VGND.n23 VGND.n22 3.764
R147 VGND.n5 VGND.n2 1.422
R148 VGND.n6 VGND.n0 0.55
R149 VGND.n8 VGND.n6 0.119
R150 VGND.n12 VGND.n8 0.119
R151 VGND.n14 VGND.n12 0.119
R152 VGND.n18 VGND.n14 0.119
R153 VGND.n20 VGND.n18 0.119
R154 VGND.n24 VGND.n20 0.119
R155 VGND.n26 VGND.n24 0.119
R156 VGND.n28 VGND.n26 0.119
R157 VGND VGND.n28 0.02
R158 a_861_47.n1 a_861_47.n0 245.478
R159 a_861_47.n0 a_861_47.t0 24.923
R160 a_861_47.n0 a_861_47.t1 24.923
R161 a_861_47.t2 a_861_47.n1 24.923
R162 a_861_47.n1 a_861_47.t3 24.923
R163 VNB VNB.t1 6053.91
R164 VNB.t9 VNB.t3 4738.46
R165 VNB.t6 VNB.t10 3868.13
R166 VNB.t4 VNB.t7 2127.47
R167 VNB.t12 VNB.t13 2030.77
R168 VNB.t2 VNB.t12 2030.77
R169 VNB.t3 VNB.t2 2030.77
R170 VNB.t10 VNB.t9 2030.77
R171 VNB.t5 VNB.t6 2030.77
R172 VNB.t7 VNB.t5 2030.77
R173 VNB.t11 VNB.t4 2030.77
R174 VNB.t8 VNB.t11 2030.77
R175 VNB.t0 VNB.t8 2030.77
R176 VNB.t1 VNB.t0 2030.77
R177 B1.n0 B1.t0 221.719
R178 B1.n1 B1.t1 221.719
R179 B1.n0 B1.t2 133.353
R180 B1.n1 B1.t3 133.353
R181 B1.n3 B1.n2 87.276
R182 B1.n2 B1.n0 58.743
R183  B1.n3 10.502
R184 B1.n3 B1 5.18
R185 B1.n2 B1.n1 4.518
R186 a_27_297.t2 a_27_297.n1 242.139
R187 a_27_297.n1 a_27_297.t0 242.137
R188 a_27_297.n1 a_27_297.n0 152.295
R189 a_27_297.n0 a_27_297.t1 26.595
R190 a_27_297.n0 a_27_297.t3 26.595
R191 A2.n3 A2.t2 252.067
R192 A2.n1 A2.t1 221.719
R193 A2.n0 A2.t0 180.659
R194 A2.n2 A2.t3 149.419
R195 A2.n0 A2 83.619
R196 A2.n4 A2.n3 76
R197 A2.n3 A2.n2 37.488
R198 A2.n1 A2.n0 36.596
R199 A2.n4 A2 20.114
R200 A2 A2.n4 7.923
R201 A2.n2 A2.n1 7.14
R202 a_1059_47.n0 a_1059_47.t0 226.776
R203 a_1059_47.n0 a_1059_47.t3 146.118
R204 a_1059_47.n1 a_1059_47.n0 50.6
R205 a_1059_47.n1 a_1059_47.t2 24.923
R206 a_1059_47.t1 a_1059_47.n1 24.923
R207 C1.n0 C1.t0 212.079
R208 C1.n1 C1.t2 212.079
R209 C1.n0 C1.t1 139.779
R210 C1.n1 C1.t3 139.779
R211 C1.n2 C1.n1 108.863
R212 C1.n1 C1.n0 61.345
R213  C1 20.241
R214 C1.n2  16.967
R215 C1 C1.n2 3.274
C0 X VGND 0.31fF
C1 VPWR VGND 0.16fF
C2 VPB VPWR 0.14fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__a311oi_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__a311oi_1 A3 Y C1 B1 A2 A1 VPWR VGND VNB VPB
X0 Y.t0 A1.t0 a_194_47.t0 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 a_194_47.t1 A2.t0 a_109_47.t1 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 Y.t2 C1.t0 a_376_297.t1 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 VPWR.t1 A2.t1 a_109_297.t1 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 Y.t3 C1.t1 VGND.t2 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 VGND.t1 B1.t0 Y.t1 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 a_109_297.t0 A1.t1 VPWR.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 a_376_297.t0 B1.t1 a_109_297.t2 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 a_109_297.t3 A3.t0 VPWR.t2 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 a_109_47.t0 A3.t1 VGND.t0 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
R0 A1.n0 A1.t1 241.534
R1 A1.n0 A1.t0 169.234
R2 A1 A1.n0 116.866
R3 a_194_47.t0 a_194_47.t1 51.692
R4 Y.n5 Y.n1 292.5
R5 Y.n4 Y.n3 153.111
R6 Y.n2 Y.t3 117.423
R7 Y.n5 Y.n4 75.544
R8 Y.n3 Y.t0 40.615
R9 Y.n1 Y.t2 26.595
R10 Y.n4 Y.n2 25.592
R11 Y.n3 Y.t1 24.923
R12 Y Y.n0 15.733
R13 Y.n2 Y 7.053
R14 Y.n0 Y 2.4
R15 Y Y.n5 2.4
R16 VNB VNB.t0 6029.73
R17 VNB.t1 VNB.t2 2441.76
R18 VNB.t2 VNB.t4 2393.41
R19 VNB.t3 VNB.t1 2079.12
R20 VNB.t0 VNB.t3 2054.95
R21 A2.n0 A2.t1 241.534
R22 A2.n0 A2.t0 169.234
R23 A2.n1 A2.n0 83.563
R24 A2 A2.n1 15.097
R25 A2.n1 A2 3.49
R26 a_109_47.t0 a_109_47.t1 50.769
R27 C1.n0 C1.t0 230.154
R28 C1.n0 C1.t1 157.854
R29 C1 C1.n0 78.909
R30 a_376_297.t0 a_376_297.t1 67.965
R31 VPB.t2 VPB.t3 292.99
R32 VPB.t0 VPB.t2 284.112
R33 VPB.t1 VPB.t0 254.517
R34 VPB.t4 VPB.t1 251.557
R35 VPB VPB.t4 186.448
R36 a_109_297.n1 a_109_297.n0 542.672
R37 a_109_297.n1 a_109_297.t2 38.415
R38 a_109_297.n0 a_109_297.t3 27.58
R39 a_109_297.n0 a_109_297.t1 26.595
R40 a_109_297.t0 a_109_297.n1 26.595
R41 VPWR.n1 VPWR.n0 327.551
R42 VPWR.n1 VPWR.t2 149.626
R43 VPWR.n0 VPWR.t0 28.565
R44 VPWR.n0 VPWR.t1 26.595
R45 VPWR VPWR.n1 0.154
R46 VGND.n1 VGND.n0 111.878
R47 VGND.n1 VGND.t0 107.385
R48 VGND.n0 VGND.t2 33.23
R49 VGND.n0 VGND.t1 30.461
R50 VGND VGND.n1 0.042
R51 B1.n0 B1.t1 241.534
R52 B1.n0 B1.t0 169.234
R53 B1 B1.n0 129.735
R54 A3.n0 A3.t0 212.152
R55 A3.n0 A3.t1 157.854
R56 A3 A3.n0 79.474
C0 C1 Y 0.13fF
C1 B1 Y 0.24fF
C2 Y VGND 0.19fF
C3 A1 A2 0.21fF
C4 A3 A2 0.11fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__a311oi_2.ext - technology: sky130A

.subckt sky130_fd_sc_hd__a311oi_2 C1 A3 Y B1 A1 A2 VGND VPWR VNB VPB
X0 Y.t2 A1.t0 a_277_47.t3 VNB.t5 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 a_641_297.t3 B1.t0 a_109_297.t7 VPB.t9 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 VPWR.t5 A1.t1 a_109_297.t5 VPB.t6 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 a_109_297.t6 B1.t1 a_641_297.t2 VPB.t8 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 a_109_297.t4 A1.t2 VPWR.t4 VPB.t5 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 a_277_47.t2 A1.t3 Y.t1 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 a_109_297.t0 A2.t0 VPWR.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 VPWR.t2 A3.t0 a_109_297.t2 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 a_27_47.t3 A3.t1 VGND.t1 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 a_27_47.t1 A2.t1 a_277_47.t0 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 VGND.t2 C1.t0 Y.t5 VNB.t8 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 VPWR.t1 A2.t2 a_109_297.t1 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 a_641_297.t1 C1.t1 Y.t6 VPB.t7 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13 a_277_47.t1 A2.t3 a_27_47.t0 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14 VGND.t5 B1.t2 Y.t3 VNB.t6 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X15 Y.t7 C1.t2 VGND.t3 VNB.t9 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X16 a_109_297.t3 A3.t2 VPWR.t3 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17 Y.t0 C1.t3 a_641_297.t0 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X18 VGND.t0 A3.t3 a_27_47.t2 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X19 Y.t4 B1.t3 VGND.t4 VNB.t7 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
R0 A1.n6 A1.t2 220.842
R1 A1.n2 A1.t1 212.079
R2 A1.n0 A1.t0 164.609
R3 A1.n1 A1.t3 139.779
R4 A1.n5 A1.n4 76
R5 A1.n7 A1.n6 76
R6 A1.n6 A1.n5 49.66
R7 A1.n1 A1.n0 36.515
R8 A1.n4 A1.n3 13.187
R9 A1.n2 A1.n1 10.224
R10 A1.n7 A1 8.921
R11 A1 A1.n7 8.921
R12 A1.n4 A1 4.266
R13 A1.n5 A1.n2 2.921
R14 A1.n3 A1 0.387
R15 a_277_47.n1 a_277_47.n0 287.4
R16 a_277_47.n0 a_277_47.t3 24.923
R17 a_277_47.n0 a_277_47.t2 24.923
R18 a_277_47.t0 a_277_47.n1 24.923
R19 a_277_47.n1 a_277_47.t1 24.923
R20 Y.n4 Y.t1 240.328
R21 Y.n6 Y.t7 233.914
R22 Y.n1 Y.n0 147.104
R23 Y.n4 Y.n3 110.194
R24 Y.n5 Y.n2 110.194
R25 Y.n2 Y.t5 71.076
R26 Y.n5 Y.n4 64
R27 Y.n3 Y.t2 28.615
R28 Y Y.n1 27.751
R29 Y.n3 Y.t3 26.769
R30 Y.n0 Y.t6 26.595
R31 Y.n0 Y.t0 26.595
R32 Y.n2 Y.t4 24.923
R33 Y.n6 Y.n5 6.776
R34 Y.n1 Y 2.439
R35 Y Y.n6 1.488
R36 VNB VNB.t3 6053.91
R37 VNB.t0 VNB.t4 4545.05
R38 VNB.t7 VNB.t8 3239.56
R39 VNB.t5 VNB.t6 2175.82
R40 VNB.t8 VNB.t9 2030.77
R41 VNB.t6 VNB.t7 2030.77
R42 VNB.t4 VNB.t5 2030.77
R43 VNB.t1 VNB.t0 2030.77
R44 VNB.t2 VNB.t1 2030.77
R45 VNB.t3 VNB.t2 2030.77
R46 B1.n0 B1.t0 212.079
R47 B1.n2 B1.t1 212.079
R48 B1.n0 B1.t3 139.779
R49 B1.n2 B1.t2 139.779
R50 B1.n1 B1 76.775
R51 B1.n4 B1.n3 76
R52 B1.n3 B1.n1 49.66
R53 B1.n4 B1 12.412
R54 B1.n1 B1.n0 10.224
R55 B1 B1.n4 5.43
R56 B1.n3 B1.n2 1.46
R57 a_109_297.n2 a_109_297.n1 239.451
R58 a_109_297.n4 a_109_297.n3 231.818
R59 a_109_297.n2 a_109_297.n0 168.571
R60 a_109_297.n5 a_109_297.n4 168.57
R61 a_109_297.n4 a_109_297.n2 65.505
R62 a_109_297.n5 a_109_297.t1 28.565
R63 a_109_297.n1 a_109_297.t7 26.595
R64 a_109_297.n1 a_109_297.t6 26.595
R65 a_109_297.n0 a_109_297.t5 26.595
R66 a_109_297.n0 a_109_297.t4 26.595
R67 a_109_297.n3 a_109_297.t2 26.595
R68 a_109_297.n3 a_109_297.t3 26.595
R69 a_109_297.t0 a_109_297.n5 26.595
R70 a_641_297.t2 a_641_297.n1 620.209
R71 a_641_297.n1 a_641_297.t1 239.936
R72 a_641_297.n1 a_641_297.n0 149.475
R73 a_641_297.n0 a_641_297.t0 55.16
R74 a_641_297.n0 a_641_297.t3 47.28
R75 VPB.t6 VPB.t8 556.386
R76 VPB.t9 VPB.t4 396.573
R77 VPB.t1 VPB.t5 260.436
R78 VPB.t0 VPB.t1 254.517
R79 VPB.t4 VPB.t7 248.598
R80 VPB.t8 VPB.t9 248.598
R81 VPB.t5 VPB.t6 248.598
R82 VPB.t2 VPB.t0 248.598
R83 VPB.t3 VPB.t2 248.598
R84 VPB VPB.t3 189.408
R85 VPWR.n2 VPWR.t5 194.537
R86 VPWR.n6 VPWR.n5 164.214
R87 VPWR.n1 VPWR.n0 163.192
R88 VPWR.n10 VPWR.t3 152.715
R89 VPWR.n0 VPWR.t4 30.535
R90 VPWR.n5 VPWR.t0 26.595
R91 VPWR.n5 VPWR.t2 26.595
R92 VPWR.n0 VPWR.t1 26.595
R93 VPWR.n4 VPWR.n3 4.65
R94 VPWR.n7 VPWR.n6 4.65
R95 VPWR.n9 VPWR.n8 4.65
R96 VPWR.n11 VPWR.n10 4.65
R97 VPWR.n2 VPWR.n1 3.903
R98 VPWR.n4 VPWR.n2 0.298
R99 VPWR.n7 VPWR.n4 0.119
R100 VPWR.n9 VPWR.n7 0.119
R101 VPWR.n11 VPWR.n9 0.119
R102 VPWR VPWR.n11 0.02
R103 A2.n0 A2.t2 213.539
R104 A2.n2 A2.t0 212.079
R105 A2.n2 A2.t3 139.779
R106 A2.n0 A2.t1 139.779
R107 A2 A2.n1 82.981
R108 A2.n4 A2.n3 76
R109 A2.n4 A2 11.636
R110 A2.n3 A2.n2 8.763
R111 A2 A2.n4 6.206
R112 A2.n1 A2.n0 2.921
R113 A3.n0 A3.t0 212.079
R114 A3.n1 A3.t2 212.079
R115 A3.n0 A3.t1 139.779
R116 A3.n1 A3.t3 139.779
R117 A3.n4 A3.n2 76
R118 A3.n2 A3.n0 43.087
R119 A3.n2 A3.n1 18.257
R120 A3.n4 A3.n3 13.187
R121 A3.n3 A3 4.072
R122 A3 A3.n4 0.581
R123 VGND.n3 VGND.n0 110.817
R124 VGND.n2 VGND.n1 107.239
R125 VGND.n17 VGND.n16 107.239
R126 VGND.n0 VGND.t3 24.923
R127 VGND.n0 VGND.t2 24.923
R128 VGND.n1 VGND.t4 24.923
R129 VGND.n1 VGND.t5 24.923
R130 VGND.n16 VGND.t1 24.923
R131 VGND.n16 VGND.t0 24.923
R132 VGND.n5 VGND.n4 4.65
R133 VGND.n7 VGND.n6 4.65
R134 VGND.n9 VGND.n8 4.65
R135 VGND.n11 VGND.n10 4.65
R136 VGND.n13 VGND.n12 4.65
R137 VGND.n15 VGND.n14 4.65
R138 VGND.n3 VGND.n2 4.07
R139 VGND.n18 VGND.n17 3.932
R140 VGND.n5 VGND.n3 0.197
R141 VGND.n18 VGND.n15 0.137
R142 VGND VGND.n18 0.121
R143 VGND.n7 VGND.n5 0.119
R144 VGND.n9 VGND.n7 0.119
R145 VGND.n11 VGND.n9 0.119
R146 VGND.n13 VGND.n11 0.119
R147 VGND.n15 VGND.n13 0.119
R148 a_27_47.t1 a_27_47.n1 238.823
R149 a_27_47.n1 a_27_47.t2 238.056
R150 a_27_47.n1 a_27_47.n0 110.194
R151 a_27_47.n0 a_27_47.t0 24.923
R152 a_27_47.n0 a_27_47.t3 24.923
R153 C1.n3 C1.t1 212.079
R154 C1.n0 C1.t3 212.079
R155 C1.n3 C1.t2 139.779
R156 C1.n0 C1.t0 139.779
R157 C1.n4 C1.n3 106.898
R158 C1.n2 C1.n1 76
R159 C1.n1 C1.n0 40.166
R160 C1.n5 C1.n2 15.709
R161 C1 C1.n5 14.161
R162 C1.n2 C1 9.6
R163 C1.n4 C1 2.995
R164 C1.n5 C1.n4 1.361
C0 VPB VPWR 0.11fF
C1 Y VGND 0.38fF
C2 VPWR VGND 0.12fF
C3 C1 Y 0.17fF
C4 B1 Y 0.20fF
C5 A1 Y 0.15fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__a311oi_4.ext - technology: sky130A

.subckt sky130_fd_sc_hd__a311oi_4 Y B1 A1 A3 C1 A2 VPWR VGND VNB VPB
X0 a_27_47.t7 A2.t0 a_445_47.t5 VNB.t19 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 a_27_47.t6 A2.t1 a_445_47.t4 VNB.t18 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 VGND.t11 C1.t0 Y.t15 VNB.t9 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 a_1139_297.t3 B1.t0 a_109_297.t9 VPB.t9 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 a_109_297.t15 A2.t2 VPWR.t11 VPB.t15 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 VPWR.t0 A3.t0 a_109_297.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 a_109_297.t8 B1.t1 a_1139_297.t2 VPB.t8 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 Y.t14 C1.t1 VGND.t10 VNB.t10 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 Y.t13 C1.t2 VGND.t9 VNB.t11 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 a_1139_297.t1 B1.t2 a_109_297.t7 VPB.t7 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 a_445_47.t0 A1.t0 Y.t0 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 a_109_297.t3 A3.t1 VPWR.t3 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 VPWR.t1 A1.t1 a_109_297.t1 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13 a_109_297.t2 A1.t2 VPWR.t2 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14 a_109_297.t6 B1.t3 a_1139_297.t0 VPB.t6 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 a_445_47.t1 A1.t3 Y.t5 VNB.t13 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X16 VGND.t3 B1.t4 Y.t1 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X17 VPWR.t4 A3.t2 a_109_297.t4 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X18 VPWR.t6 A1.t4 a_109_297.t10 VPB.t10 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X19 a_1139_297.t7 C1.t3 Y.t11 VPB.t19 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X20 a_27_47.t0 A3.t3 VGND.t0 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X21 a_27_47.t1 A3.t4 VGND.t1 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X22 VGND.t8 C1.t4 Y.t12 VNB.t12 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X23 a_109_297.t11 A1.t5 VPWR.t7 VPB.t11 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X24 Y.t10 C1.t5 a_1139_297.t6 VPB.t18 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X25 Y.t6 A1.t6 a_445_47.t2 VNB.t14 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X26 VPWR.t10 A2.t3 a_109_297.t14 VPB.t14 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X27 a_1139_297.t5 C1.t6 Y.t9 VPB.t17 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X28 Y.t7 A1.t7 a_445_47.t3 VNB.t15 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X29 Y.t2 B1.t5 VGND.t4 VNB.t5 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X30 Y.t3 B1.t6 VGND.t5 VNB.t6 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X31 VGND.t2 A3.t5 a_27_47.t2 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X32 a_445_47.t7 A2.t4 a_27_47.t5 VNB.t17 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X33 a_109_297.t13 A2.t5 VPWR.t9 VPB.t13 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X34 Y.t8 C1.t7 a_1139_297.t4 VPB.t16 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X35 a_445_47.t6 A2.t6 a_27_47.t4 VNB.t16 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X36 VPWR.t8 A2.t7 a_109_297.t12 VPB.t12 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X37 VGND.t6 B1.t7 Y.t4 VNB.t7 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X38 a_109_297.t5 A3.t6 VPWR.t5 VPB.t5 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X39 VGND.t7 A3.t7 a_27_47.t3 VNB.t8 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
R0 A2.n0 A2.t3 212.079
R1 A2.n2 A2.t5 212.079
R2 A2.n3 A2.t7 212.079
R3 A2.n4 A2.t2 212.079
R4 A2.n0 A2.t1 139.779
R5 A2.n2 A2.t6 139.779
R6 A2.n3 A2.t0 139.779
R7 A2.n4 A2.t4 139.779
R8 A2.n11 A2.n1 76
R9 A2.n10 A2.n9 76
R10 A2.n8 A2.n7 76
R11 A2.n6 A2.n5 76
R12 A2.n9 A2.n8 54.042
R13 A2.n5 A2.n3 52.581
R14 A2.n11 A2.n10 14.351
R15 A2.n1 A2.n0 13.145
R16 A2.n7 A2 12.8
R17 A2 A2.n6 9.309
R18 A2.n5 A2.n4 8.763
R19 A2.n6 A2 8.533
R20 A2.n9 A2.n2 5.842
R21 A2.n7 A2 5.042
R22 A2 A2.n11 1.939
R23 A2.n10 A2 1.551
R24 A2.n8 A2.n3 1.46
R25 a_445_47.n5 a_445_47.n4 155.747
R26 a_445_47.n3 a_445_47.n2 155.747
R27 a_445_47.n4 a_445_47.n3 102.4
R28 a_445_47.n4 a_445_47.n0 92.5
R29 a_445_47.n3 a_445_47.n1 92.5
R30 a_445_47.n2 a_445_47.t5 24.923
R31 a_445_47.n2 a_445_47.t7 24.923
R32 a_445_47.n1 a_445_47.t4 24.923
R33 a_445_47.n1 a_445_47.t6 24.923
R34 a_445_47.n0 a_445_47.t3 24.923
R35 a_445_47.n0 a_445_47.t1 24.923
R36 a_445_47.n5 a_445_47.t2 24.923
R37 a_445_47.t0 a_445_47.n5 24.923
R38 a_27_47.n3 a_27_47.t3 236.55
R39 a_27_47.t6 a_27_47.n5 229.593
R40 a_27_47.n3 a_27_47.n2 108.688
R41 a_27_47.n4 a_27_47.n1 108.688
R42 a_27_47.n5 a_27_47.n0 92.5
R43 a_27_47.n5 a_27_47.n4 63.247
R44 a_27_47.n4 a_27_47.n3 63.247
R45 a_27_47.n0 a_27_47.t4 24.923
R46 a_27_47.n0 a_27_47.t7 24.923
R47 a_27_47.n2 a_27_47.t2 24.923
R48 a_27_47.n2 a_27_47.t0 24.923
R49 a_27_47.n1 a_27_47.t5 24.923
R50 a_27_47.n1 a_27_47.t1 24.923
R51 VNB VNB.t8 6053.91
R52 VNB.t18 VNB.t13 4545.05
R53 VNB.t6 VNB.t9 3094.5
R54 VNB.t12 VNB.t11 2030.77
R55 VNB.t10 VNB.t12 2030.77
R56 VNB.t9 VNB.t10 2030.77
R57 VNB.t7 VNB.t6 2030.77
R58 VNB.t5 VNB.t7 2030.77
R59 VNB.t4 VNB.t5 2030.77
R60 VNB.t14 VNB.t4 2030.77
R61 VNB.t0 VNB.t14 2030.77
R62 VNB.t15 VNB.t0 2030.77
R63 VNB.t13 VNB.t15 2030.77
R64 VNB.t16 VNB.t18 2030.77
R65 VNB.t19 VNB.t16 2030.77
R66 VNB.t17 VNB.t19 2030.77
R67 VNB.t2 VNB.t17 2030.77
R68 VNB.t3 VNB.t2 2030.77
R69 VNB.t1 VNB.t3 2030.77
R70 VNB.t8 VNB.t1 2030.77
R71 C1.n0 C1.t3 212.079
R72 C1.n7 C1.t5 212.079
R73 C1.n1 C1.t6 212.079
R74 C1.n2 C1.t7 212.079
R75 C1.n0 C1.t2 139.779
R76 C1.n7 C1.t4 139.779
R77 C1.n1 C1.t1 139.779
R78 C1.n2 C1.t0 139.779
R79 C1.n9 C1.n8 76
R80 C1.n6 C1.n5 76
R81 C1.n4 C1.n3 76
R82 C1.n3 C1.n2 54.772
R83 C1.n6 C1.n1 47.469
R84 C1.n8 C1.n7 40.166
R85 C1.n8 C1.n0 21.178
R86 C1.n7 C1.n6 13.875
R87 C1.n4 C1 13.381
R88 C1 C1.n9 11.442
R89 C1.n5 C1 9.89
R90 C1.n5 C1 7.951
R91 C1.n3 C1.n1 6.572
R92 C1.n9 C1 6.4
R93 C1 C1.n4 4.46
R94 Y.n11 Y.t13 236.55
R95 Y.n7 Y.t5 229.593
R96 Y.n2 Y.n0 188.153
R97 Y.n2 Y.n1 149.753
R98 Y.n13 Y.n12 112.088
R99 Y.n11 Y.n10 108.688
R100 Y.n9 Y.n4 108.688
R101 Y.n7 Y.n6 92.5
R102 Y.n8 Y.n5 92.5
R103 Y.n12 Y.t15 65.538
R104 Y.n9 Y.n8 63.247
R105 Y.n8 Y.n7 63.247
R106 Y.n13 Y.n11 62.117
R107 Y.n13 Y.n9 56.847
R108 Y.n0 Y.t11 26.595
R109 Y.n0 Y.t10 26.595
R110 Y.n1 Y.t9 26.595
R111 Y.n1 Y.t8 26.595
R112 Y.n10 Y.t12 24.923
R113 Y.n10 Y.t14 24.923
R114 Y.n5 Y.t1 24.923
R115 Y.n5 Y.t6 24.923
R116 Y.n6 Y.t0 24.923
R117 Y.n6 Y.t7 24.923
R118 Y.n4 Y.t4 24.923
R119 Y.n4 Y.t2 24.923
R120 Y.n12 Y.t3 24.923
R121 Y.n3 Y.n2 18.07
R122 Y Y.n3 7.4
R123 Y.n3 Y 6.2
R124 Y Y.n13 1.8
R125 VGND.n3 VGND.n0 110.747
R126 VGND.n2 VGND.n1 107.239
R127 VGND.n7 VGND.n6 107.239
R128 VGND.n12 VGND.n11 107.239
R129 VGND.n33 VGND.n32 107.239
R130 VGND.n38 VGND.n37 107.239
R131 VGND.n0 VGND.t9 24.923
R132 VGND.n0 VGND.t8 24.923
R133 VGND.n1 VGND.t10 24.923
R134 VGND.n1 VGND.t11 24.923
R135 VGND.n6 VGND.t5 24.923
R136 VGND.n6 VGND.t6 24.923
R137 VGND.n11 VGND.t4 24.923
R138 VGND.n11 VGND.t3 24.923
R139 VGND.n32 VGND.t1 24.923
R140 VGND.n32 VGND.t2 24.923
R141 VGND.n37 VGND.t0 24.923
R142 VGND.n37 VGND.t7 24.923
R143 VGND.n5 VGND.n4 4.65
R144 VGND.n8 VGND.n7 4.65
R145 VGND.n10 VGND.n9 4.65
R146 VGND.n13 VGND.n12 4.65
R147 VGND.n15 VGND.n14 4.65
R148 VGND.n17 VGND.n16 4.65
R149 VGND.n19 VGND.n18 4.65
R150 VGND.n21 VGND.n20 4.65
R151 VGND.n23 VGND.n22 4.65
R152 VGND.n25 VGND.n24 4.65
R153 VGND.n27 VGND.n26 4.65
R154 VGND.n29 VGND.n28 4.65
R155 VGND.n31 VGND.n30 4.65
R156 VGND.n34 VGND.n33 4.65
R157 VGND.n36 VGND.n35 4.65
R158 VGND.n39 VGND.n38 3.932
R159 VGND.n3 VGND.n2 3.618
R160 VGND.n5 VGND.n3 0.257
R161 VGND.n39 VGND.n36 0.137
R162 VGND VGND.n39 0.121
R163 VGND.n8 VGND.n5 0.119
R164 VGND.n10 VGND.n8 0.119
R165 VGND.n13 VGND.n10 0.119
R166 VGND.n15 VGND.n13 0.119
R167 VGND.n17 VGND.n15 0.119
R168 VGND.n19 VGND.n17 0.119
R169 VGND.n21 VGND.n19 0.119
R170 VGND.n23 VGND.n21 0.119
R171 VGND.n25 VGND.n23 0.119
R172 VGND.n27 VGND.n25 0.119
R173 VGND.n29 VGND.n27 0.119
R174 VGND.n31 VGND.n29 0.119
R175 VGND.n34 VGND.n31 0.119
R176 VGND.n36 VGND.n34 0.119
R177 B1.n6 B1.t3 212.079
R178 B1.n1 B1.t0 212.079
R179 B1.n2 B1.t1 212.079
R180 B1.n0 B1.t2 212.079
R181 B1.n6 B1.t4 139.779
R182 B1.n1 B1.t6 139.779
R183 B1.n2 B1.t7 139.779
R184 B1.n0 B1.t5 139.779
R185 B1 B1.n3 79.225
R186 B1.n5 B1.n4 76
R187 B1.n7 B1.n6 76
R188 B1.n2 B1.n1 61.345
R189 B1.n6 B1.n5 54.042
R190 B1.n3 B1.n0 46.739
R191 B1.n3 B1.n2 14.606
R192 B1.n5 B1.n0 7.303
R193 B1 B1.n7 6.853
R194 B1.n4 B1 5.039
R195 B1.n4 B1 4.233
R196 B1.n7 B1 2.418
R197 a_109_297.n5 a_109_297.n3 355.747
R198 a_109_297.n5 a_109_297.n4 292.5
R199 a_109_297.n12 a_109_297.n11 237.841
R200 a_109_297.n8 a_109_297.n2 174.594
R201 a_109_297.n9 a_109_297.n1 174.594
R202 a_109_297.n10 a_109_297.n0 174.594
R203 a_109_297.n13 a_109_297.n12 174.593
R204 a_109_297.n7 a_109_297.n6 150.188
R205 a_109_297.n7 a_109_297.n5 102.4
R206 a_109_297.n8 a_109_297.n7 82.07
R207 a_109_297.n9 a_109_297.n8 63.247
R208 a_109_297.n10 a_109_297.n9 63.247
R209 a_109_297.n12 a_109_297.n10 63.247
R210 a_109_297.n6 a_109_297.t1 26.595
R211 a_109_297.n6 a_109_297.t2 26.595
R212 a_109_297.n4 a_109_297.t7 26.595
R213 a_109_297.n4 a_109_297.t6 26.595
R214 a_109_297.n3 a_109_297.t9 26.595
R215 a_109_297.n3 a_109_297.t8 26.595
R216 a_109_297.n2 a_109_297.t10 26.595
R217 a_109_297.n2 a_109_297.t11 26.595
R218 a_109_297.n1 a_109_297.t14 26.595
R219 a_109_297.n1 a_109_297.t13 26.595
R220 a_109_297.n0 a_109_297.t12 26.595
R221 a_109_297.n0 a_109_297.t15 26.595
R222 a_109_297.n11 a_109_297.t4 26.595
R223 a_109_297.n11 a_109_297.t5 26.595
R224 a_109_297.t0 a_109_297.n13 26.595
R225 a_109_297.n13 a_109_297.t3 26.595
R226 a_1139_297.n3 a_1139_297.t0 624.727
R227 a_1139_297.n1 a_1139_297.n0 292.5
R228 a_1139_297.n3 a_1139_297.n2 292.5
R229 a_1139_297.n5 a_1139_297.n4 292.5
R230 a_1139_297.n1 a_1139_297.t7 233.919
R231 a_1139_297.n4 a_1139_297.n1 79.811
R232 a_1139_297.n5 a_1139_297.t4 69.935
R233 a_1139_297.n4 a_1139_297.n3 63.247
R234 a_1139_297.n2 a_1139_297.t2 26.595
R235 a_1139_297.n2 a_1139_297.t1 26.595
R236 a_1139_297.n0 a_1139_297.t6 26.595
R237 a_1139_297.n0 a_1139_297.t5 26.595
R238 a_1139_297.t3 a_1139_297.n5 26.595
R239 VPB.t1 VPB.t6 556.386
R240 VPB.t9 VPB.t16 378.816
R241 VPB.t18 VPB.t19 248.598
R242 VPB.t17 VPB.t18 248.598
R243 VPB.t16 VPB.t17 248.598
R244 VPB.t8 VPB.t9 248.598
R245 VPB.t7 VPB.t8 248.598
R246 VPB.t6 VPB.t7 248.598
R247 VPB.t2 VPB.t1 248.598
R248 VPB.t10 VPB.t2 248.598
R249 VPB.t11 VPB.t10 248.598
R250 VPB.t14 VPB.t11 248.598
R251 VPB.t13 VPB.t14 248.598
R252 VPB.t12 VPB.t13 248.598
R253 VPB.t15 VPB.t12 248.598
R254 VPB.t0 VPB.t15 248.598
R255 VPB.t3 VPB.t0 248.598
R256 VPB.t4 VPB.t3 248.598
R257 VPB.t5 VPB.t4 248.598
R258 VPB VPB.t5 189.408
R259 VPWR.n2 VPWR.t1 579.719
R260 VPWR.n21 VPWR.n20 164.214
R261 VPWR.n16 VPWR.n15 164.214
R262 VPWR.n10 VPWR.n9 164.214
R263 VPWR.n6 VPWR.n5 164.214
R264 VPWR.n1 VPWR.n0 164.214
R265 VPWR.n25 VPWR.t5 145.867
R266 VPWR.n20 VPWR.t3 26.595
R267 VPWR.n20 VPWR.t4 26.595
R268 VPWR.n15 VPWR.t11 26.595
R269 VPWR.n15 VPWR.t0 26.595
R270 VPWR.n9 VPWR.t9 26.595
R271 VPWR.n9 VPWR.t8 26.595
R272 VPWR.n5 VPWR.t7 26.595
R273 VPWR.n5 VPWR.t10 26.595
R274 VPWR.n0 VPWR.t2 26.595
R275 VPWR.n0 VPWR.t6 26.595
R276 VPWR.n4 VPWR.n3 4.65
R277 VPWR.n8 VPWR.n7 4.65
R278 VPWR.n12 VPWR.n11 4.65
R279 VPWR.n14 VPWR.n13 4.65
R280 VPWR.n17 VPWR.n16 4.65
R281 VPWR.n19 VPWR.n18 4.65
R282 VPWR.n22 VPWR.n21 4.65
R283 VPWR.n24 VPWR.n23 4.65
R284 VPWR.n26 VPWR.n25 4.65
R285 VPWR.n2 VPWR.n1 3.618
R286 VPWR.n11 VPWR.n10 3.388
R287 VPWR.n7 VPWR.n6 0.376
R288 VPWR.n4 VPWR.n2 0.257
R289 VPWR.n8 VPWR.n4 0.119
R290 VPWR.n12 VPWR.n8 0.119
R291 VPWR.n14 VPWR.n12 0.119
R292 VPWR.n17 VPWR.n14 0.119
R293 VPWR.n19 VPWR.n17 0.119
R294 VPWR.n22 VPWR.n19 0.119
R295 VPWR.n24 VPWR.n22 0.119
R296 VPWR.n26 VPWR.n24 0.119
R297 VPWR VPWR.n26 0.02
R298 A3.n1 A3.t0 212.079
R299 A3.n3 A3.t1 212.079
R300 A3.n0 A3.t2 212.079
R301 A3.n9 A3.t6 212.079
R302 A3.n1 A3.t4 139.779
R303 A3.n3 A3.t5 139.779
R304 A3.n0 A3.t3 139.779
R305 A3.n9 A3.t7 139.779
R306 A3.n10 A3.n9 103.021
R307 A3.n5 A3.n4 76
R308 A3.n8 A3.n7 76
R309 A3.n4 A3.n1 48.93
R310 A3.n3 A3.n2 41.627
R311 A3.n8 A3.n0 34.324
R312 A3.n9 A3.n8 27.021
R313 A3.n2 A3.n0 19.718
R314 A3.n7 A3.n6 14.351
R315 A3 A3.n5 12.606
R316 A3.n10 A3 12.606
R317 A3.n4 A3.n3 12.415
R318 A3.n5 A3 5.236
R319 A3 A3.n10 5.236
R320 A3.n6 A3 1.745
R321 A3.n7 A3 1.745
R322 A1.n8 A1.t5 213.914
R323 A1.n1 A1.t1 205.652
R324 A1.n5 A1.t2 205.652
R325 A1.n11 A1.t4 205.652
R326 A1.n0 A1.t6 200.628
R327 A1.n10 A1.t3 139.779
R328 A1.n4 A1.t7 139.779
R329 A1.n0 A1.t0 137.677
R330 A1.n3 A1.n2 76
R331 A1.n7 A1.n6 76
R332 A1.n13 A1.n12 76
R333 A1.n9 A1.n8 76
R334 A1.n4 A1.n3 31.674
R335 A1.n13 A1.n9 14.351
R336 A1.n5 A1.n4 13.771
R337 A1.n1 A1.n0 13.196
R338 A1 A1.n7 13.187
R339 A1.n3 A1.n1 12.394
R340 A1.n12 A1.n10 12.394
R341 A1.n2 A1 9.696
R342 A1.n2 A1 8.145
R343 A1.n6 A1.n5 5.508
R344 A1.n7 A1 4.654
R345 A1.n9 A1 2.327
R346 A1.n12 A1.n11 1.377
R347 A1 A1.n13 1.163
C0 Y VGND 0.67fF
C1 VPWR VGND 0.20fF
C2 VPWR VPB 0.19fF
C3 A3 A2 0.10fF
C4 Y C1 0.50fF
C5 Y B1 0.22fF
C6 Y A1 0.24fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__a2111o_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__a2111o_1 VGND VPWR B1 X D1 A1 A2 C1 VNB VPB
X0 VGND.t3 A2.t0 a_660_47.t1 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 VGND.t1 C1.t0 a_85_193.t0 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 a_414_297.t0 C1.t1 a_334_297.t0 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 VGND.t0 a_85_193.t5 X.t1 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 a_334_297.t1 D1.t0 a_85_193.t3 VPB.t5 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 a_516_297.t1 B1.t0 a_414_297.t1 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 a_516_297.t2 A2.t1 VPWR.t2 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 a_660_47.t0 A1.t0 a_85_193.t2 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 a_85_193.t4 D1.t1 VGND.t4 VNB.t5 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 VPWR.t1 A1.t1 a_516_297.t0 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 a_85_193.t1 B1.t1 VGND.t2 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 VPWR.t0 a_85_193.t6 X.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
R0 A2.n0 A2.t1 235.47
R1 A2.n0 A2.t0 157.783
R2 A2 A2.n0 81.554
R3 a_660_47.t0 a_660_47.t1 47.076
R4 VGND.n0 VGND.t3 147.874
R5 VGND.n2 VGND.n1 107.34
R6 VGND.n8 VGND.n7 92.5
R7 VGND.n12 VGND.n11 92.5
R8 VGND.n7 VGND.t4 58.153
R9 VGND.n11 VGND.t0 34.153
R10 VGND.n1 VGND.t2 33.23
R11 VGND.n1 VGND.t1 33.23
R12 VGND.n13 VGND.n12 6.648
R13 VGND.n10 VGND.n9 4.65
R14 VGND.n4 VGND.n3 4.65
R15 VGND.n6 VGND.n5 4.65
R16 VGND.n3 VGND.n2 1.129
R17 VGND.n4 VGND.n0 0.142
R18 VGND.n13 VGND.n10 0.133
R19 VGND VGND.n13 0.128
R20 VGND.n6 VGND.n4 0.119
R21 VGND.n10 VGND.n6 0.119
R22 VGND.n9 VGND.n8 0.115
R23 VNB VNB.t0 6416.55
R24 VNB.n0 VNB 4917.65
R25 VNB.t0 VNB.t5 4810.99
R26 VNB.t2 VNB.t3 3481.32
R27 VNB.t5 VNB.t1 2224.18
R28 VNB.n0 VNB.t2 2103.3
R29 VNB.t3 VNB.t4 1958.24
R30 VNB.t1 VNB.n0 362.637
R31 C1.n0 C1.t1 229.752
R32 C1.n0 C1.t0 166.289
R33 C1.n1 C1.n0 76
R34 C1 C1.n1 11.054
R35 C1.n1 C1 2.133
R36 a_85_193.n0 a_85_193.t5 1784.9
R37 a_85_193.t3 a_85_193.n4 284.569
R38 a_85_193.n0 a_85_193.t6 223.475
R39 a_85_193.n3 a_85_193.n1 159.254
R40 a_85_193.n1 a_85_193.t2 79.384
R41 a_85_193.n4 a_85_193.n0 76
R42 a_85_193.n4 a_85_193.n3 73.732
R43 a_85_193.n3 a_85_193.n2 49.521
R44 a_85_193.n2 a_85_193.t0 31.384
R45 a_85_193.n2 a_85_193.t4 25.846
R46 a_85_193.n1 a_85_193.t1 25.846
R47 a_334_297.t0 a_334_297.t1 49.25
R48 a_414_297.t0 a_414_297.t1 70.92
R49 VPB.t0 VPB.t5 648.13
R50 VPB.t3 VPB.t2 420.249
R51 VPB.t1 VPB.t3 301.869
R52 VPB.t2 VPB.t4 248.598
R53 VPB.t5 VPB.t1 236.76
R54 VPB VPB.t0 210.124
R55 X.n2 X.n1 292.5
R56 X.n1 X.n0 146.251
R57 X X.n4 93.469
R58 X.n4 X.t1 30.461
R59 X.n1 X.t0 28.565
R60 X.n0 X 12.679
R61 X X.n3 12.218
R62 X.n2 X 8.669
R63 X X.n2 6.4
R64 X.n0 X 4.267
R65 X.n3 X 0.969
R66 D1.n0 D1.t0 234.801
R67 D1.n0 D1.t1 162.501
R68 D1.n1 D1.n0 76
R69 D1 D1.n1 13.547
R70 D1.n1 D1 1.637
R71 B1.n0 B1.t0 235.302
R72 B1.n0 B1.t1 157.745
R73 B1.n1 B1.n0 76
R74 B1.n1 B1 13.028
R75 B1 B1.n1 2.514
R76 a_516_297.n0 a_516_297.t2 395.414
R77 a_516_297.n0 a_516_297.t1 83.725
R78 a_516_297.t0 a_516_297.n0 26.595
R79 VPWR.n1 VPWR.t0 195.974
R80 VPWR.n1 VPWR.n0 177.727
R81 VPWR.n0 VPWR.t2 26.595
R82 VPWR.n0 VPWR.t1 26.595
R83 VPWR VPWR.n1 0.147
R84 A1.n0 A1.t1 1053.26
R85 A1.n0 A1.t0 157.783
R86 A1.n1 A1.n0 76.387
R87 A1.n1 A1 15.981
R88 A1 A1.n1 8.921
C0 A1 VGND 0.16fF
C1 C1 B1 0.27fF
C2 X VPWR 0.14fF
C3 C1 D1 0.19fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__a2111o_2.ext - technology: sky130A

.subckt sky130_fd_sc_hd__a2111o_2 D1 A1 B1 C1 X A2 VGND VPWR VNB VPB
X0 VPWR.t3 a_86_235.t5 X.t1 VPB.t6 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 VGND.t5 C1.t0 a_86_235.t0 VNB.t6 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 X.t0 a_86_235.t6 VPWR.t2 VPB.t5 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 a_86_235.t3 D1.t0 VGND.t2 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 X.t3 a_86_235.t7 VGND.t4 VNB.t5 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 a_715_47.t0 A1.t0 a_86_235.t2 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 VGND.t1 A2.t0 a_715_47.t1 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 a_499_297.t1 C1.t1 a_427_297.t1 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 VGND.t3 a_86_235.t8 X.t2 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 a_86_235.t1 B1.t0 VGND.t0 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 a_607_297.t1 B1.t1 a_499_297.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 a_427_297.t0 D1.t1 a_86_235.t4 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 VPWR.t1 A1.t1 a_607_297.t0 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13 a_607_297.t2 A2.t1 VPWR.t0 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
R0 a_86_235.t4 a_86_235.n6 247.685
R1 a_86_235.n3 a_86_235.t6 227.544
R2 a_86_235.n4 a_86_235.t5 212.079
R3 a_86_235.n2 a_86_235.n0 157.575
R4 a_86_235.n3 a_86_235.t7 139.779
R5 a_86_235.n5 a_86_235.t8 139.779
R6 a_86_235.n6 a_86_235.n5 128.244
R7 a_86_235.n2 a_86_235.n1 107.433
R8 a_86_235.n6 a_86_235.n2 58.621
R9 a_86_235.n4 a_86_235.n3 51.121
R10 a_86_235.n0 a_86_235.t2 36
R11 a_86_235.n0 a_86_235.t1 25.846
R12 a_86_235.n1 a_86_235.t0 25.846
R13 a_86_235.n1 a_86_235.t3 25.846
R14 a_86_235.n5 a_86_235.n4 11.684
R15 X.n3 X.n0 292.5
R16 X.n4 X.n0 292.5
R17 X X.n1 92.72
R18 X.n2 X.n1 92.5
R19 X.n0 X.t1 27.58
R20 X.n0 X.t0 27.58
R21 X.n1 X.t2 25.846
R22 X.n1 X.t3 25.846
R23 X.n2 X 14.786
R24 X.n4 X 11.696
R25 X.n3 X 11.696
R26 X X.n4 3.31
R27 X X.n3 3.31
R28 X X.n2 0.22
R29 VPWR.n2 VPWR.n0 311.121
R30 VPWR.n5 VPWR.t2 257.773
R31 VPWR.n1 VPWR.t3 153.701
R32 VPWR.n0 VPWR.t0 41.37
R33 VPWR.n0 VPWR.t1 35.46
R34 VPWR.n4 VPWR.n3 4.65
R35 VPWR.n6 VPWR.n5 4.65
R36 VPWR.n2 VPWR.n1 3.936
R37 VPWR.n4 VPWR.n2 0.14
R38 VPWR.n6 VPWR.n4 0.119
R39 VPWR VPWR.n6 0.022
R40 VPB.t6 VPB.t4 665.887
R41 VPB.t3 VPB.t2 319.626
R42 VPB.t0 VPB.t3 319.626
R43 VPB.t1 VPB.t0 319.626
R44 VPB.t5 VPB.t6 254.517
R45 VPB.t4 VPB.t1 213.084
R46 VPB VPB.t5 213.084
R47 C1.n0 C1.t1 236.179
R48 C1.n0 C1.t0 163.879
R49 C1.n1 C1.n0 76
R50 C1 C1.n1 11.767
R51 C1.n1 C1 2.27
R52 VGND.n0 VGND.t1 106.926
R53 VGND.n2 VGND.n1 106.463
R54 VGND.n17 VGND.t4 92.599
R55 VGND.n8 VGND.n7 92.5
R56 VGND.n12 VGND.n11 48.98
R57 VGND.n1 VGND.t5 35.076
R58 VGND.n1 VGND.t0 34.153
R59 VGND.n7 VGND.t2 25.846
R60 VGND.n11 VGND.t3 25.846
R61 VGND.n9 VGND.n8 5.675
R62 VGND.n18 VGND.n17 4.65
R63 VGND.n4 VGND.n3 4.65
R64 VGND.n6 VGND.n5 4.65
R65 VGND.n10 VGND.n9 4.65
R66 VGND.n14 VGND.n13 4.65
R67 VGND.n16 VGND.n15 4.65
R68 VGND.n3 VGND.n2 4.517
R69 VGND.n13 VGND.n12 1.534
R70 VGND.n4 VGND.n0 0.143
R71 VGND.n6 VGND.n4 0.119
R72 VGND.n10 VGND.n6 0.119
R73 VGND.n14 VGND.n10 0.119
R74 VGND.n16 VGND.n14 0.119
R75 VGND.n18 VGND.n16 0.119
R76 VGND VGND.n18 0.022
R77 VNB VNB.t5 6634.13
R78 VNB.t4 VNB.t3 5052.75
R79 VNB.t1 VNB.t2 2610.99
R80 VNB.t6 VNB.t0 2538.46
R81 VNB.t0 VNB.t1 2345.05
R82 VNB.t3 VNB.t6 2079.12
R83 VNB.t5 VNB.t4 2079.12
R84 D1.n0 D1.t1 236.179
R85 D1.n0 D1.t0 163.879
R86 D1.n1 D1.n0 76
R87 D1 D1.n1 10.914
R88 D1.n1 D1 1.902
R89 A1.n0 A1.t1 236.179
R90 A1.n0 A1.t0 161.249
R91 A1.n1 A1.n0 76
R92 A1 A1.n1 8.897
R93 A1.n1 A1 1.717
R94 a_715_47.t0 a_715_47.t1 72
R95 A2.n0 A2.t1 236.179
R96 A2.n0 A2.t0 163.879
R97 A2.n1 A2.n0 76
R98 A2.n1 A2 6.4
R99 A2 A2.n1 1.235
R100 a_427_297.t0 a_427_297.t1 41.37
R101 a_499_297.t0 a_499_297.t1 76.83
R102 B1.n0 B1.t1 236.179
R103 B1.n0 B1.t0 163.879
R104 B1.n1 B1.n0 76
R105 B1.n1 B1 12.579
R106 B1 B1.n1 2.427
R107 a_607_297.n0 a_607_297.t2 377.774
R108 a_607_297.n0 a_607_297.t1 39.4
R109 a_607_297.t0 a_607_297.n0 37.43
C0 VPWR X 0.25fF
C1 A1 A2 0.18fF
C2 B1 A1 0.17fF
C3 C1 B1 0.17fF
C4 C1 D1 0.20fF
C5 VGND X 0.22fF
C6 VGND VPWR 0.12fF
C7 A1 VGND 0.17fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__a2111o_4.ext - technology: sky130A

.subckt sky130_fd_sc_hd__a2111o_4 C1 B1 A1 A2 X D1 VGND VPWR VNB VPB
X0 a_30_297.t3 C1.t0 a_285_297.t3 VPB.t12 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 VGND.t10 C1.t1 a_44_47.t8 VNB.t12 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 a_44_47.t2 B1.t0 VGND.t0 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 VGND.t5 a_44_47.t10 X.t7 VNB.t7 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 VPWR.t7 A1.t0 a_477_297.t5 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 VPWR.t3 a_44_47.t11 X.t3 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 X.t6 a_44_47.t12 VGND.t4 VNB.t6 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 VGND.t1 B1.t1 a_44_47.t3 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 X.t5 a_44_47.t13 VGND.t3 VNB.t5 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 a_477_297.t4 A1.t1 VPWR.t6 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 a_285_297.t0 B1.t2 a_477_297.t3 VPB.t5 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 VGND.t7 D1.t0 a_44_47.t4 VNB.t9 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 a_770_47.t3 A2.t0 VGND.t11 VNB.t13 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 X.t2 a_44_47.t14 VPWR.t2 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14 a_30_297.t0 D1.t1 a_44_47.t5 VPB.t9 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 VGND.t6 A2.t1 a_770_47.t2 VNB.t8 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X16 a_44_47.t6 D1.t2 a_30_297.t1 VPB.t10 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17 a_477_297.t2 B1.t3 a_285_297.t1 VPB.t6 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X18 a_770_47.t1 A1.t2 a_44_47.t0 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X19 a_477_297.t0 A2.t2 VPWR.t4 VPB.t7 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X20 VPWR.t1 a_44_47.t15 X.t1 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X21 a_285_297.t2 C1.t2 a_30_297.t2 VPB.t11 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X22 a_44_47.t7 D1.t3 VGND.t8 VNB.t10 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X23 a_44_47.t1 A1.t3 a_770_47.t0 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X24 VGND.t2 a_44_47.t16 X.t4 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X25 VPWR.t5 A2.t3 a_477_297.t1 VPB.t8 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X26 X.t0 a_44_47.t17 VPWR.t0 VPB.t13 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X27 a_44_47.t9 C1.t3 VGND.t9 VNB.t11 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
R0 C1.n2 C1.t2 224.067
R1 C1.n1 C1.t0 213.686
R2 C1.n0 C1.t3 144.969
R3 C1.n2 C1.t1 139.779
R4 C1.n5 C1.n0 76
R5 C1.n4 C1.n3 76
R6 C1.n3 C1.n1 40.043
R7 C1.n4 C1 18.374
R8 C1.n5 C1 13.419
R9 C1.n3 C1.n2 13.347
R10 C1.n1 C1.n0 10.381
R11 C1 C1.n5 5.574
R12 C1 C1.n4 0.619
R13 a_285_297.n1 a_285_297.n0 392.88
R14 a_285_297.n0 a_285_297.t3 27.58
R15 a_285_297.n0 a_285_297.t2 27.58
R16 a_285_297.n1 a_285_297.t1 27.58
R17 a_285_297.t0 a_285_297.n1 27.58
R18 a_30_297.n0 a_30_297.t1 232.284
R19 a_30_297.n0 a_30_297.t3 231.299
R20 a_30_297.n1 a_30_297.n0 114.752
R21 a_30_297.t2 a_30_297.n1 27.58
R22 a_30_297.n1 a_30_297.t0 27.58
R23 VPB.t4 VPB.t7 556.386
R24 VPB.t12 VPB.t5 556.386
R25 VPB.t6 VPB.t3 393.613
R26 VPB.t1 VPB.t2 254.517
R27 VPB.t0 VPB.t1 254.517
R28 VPB.t13 VPB.t0 254.517
R29 VPB.t8 VPB.t13 254.517
R30 VPB.t7 VPB.t8 254.517
R31 VPB.t3 VPB.t4 254.517
R32 VPB.t5 VPB.t6 254.517
R33 VPB.t11 VPB.t12 254.517
R34 VPB.t9 VPB.t11 254.517
R35 VPB.t10 VPB.t9 254.517
R36 VPB VPB.t10 204.205
R37 a_44_47.n11 a_44_47.t1 241.207
R38 a_44_47.n12 a_44_47.n9 240.068
R39 a_44_47.n5 a_44_47.t11 212.079
R40 a_44_47.n0 a_44_47.t15 212.079
R41 a_44_47.n2 a_44_47.t14 212.079
R42 a_44_47.n7 a_44_47.t17 212.079
R43 a_44_47.n18 a_44_47.n17 186.324
R44 a_44_47.n17 a_44_47.t4 140.644
R45 a_44_47.n5 a_44_47.t10 139.779
R46 a_44_47.n0 a_44_47.t16 139.779
R47 a_44_47.n2 a_44_47.t12 139.779
R48 a_44_47.n7 a_44_47.t13 139.779
R49 a_44_47.n14 a_44_47.n13 108.997
R50 a_44_47.n16 a_44_47.n15 108.639
R51 a_44_47.n4 a_44_47.n1 101.6
R52 a_44_47.n14 a_44_47.n12 88.926
R53 a_44_47.n4 a_44_47.n3 76
R54 a_44_47.n6 a_44_47.n5 76
R55 a_44_47.n9 a_44_47.n8 76
R56 a_44_47.n16 a_44_47.n14 45.473
R57 a_44_47.n11 a_44_47.n10 43.555
R58 a_44_47.n13 a_44_47.t3 36
R59 a_44_47.t5 a_44_47.n18 27.58
R60 a_44_47.n18 a_44_47.t6 27.58
R61 a_44_47.n10 a_44_47.t2 26.769
R62 a_44_47.n1 a_44_47.n0 26.29
R63 a_44_47.n15 a_44_47.t8 25.846
R64 a_44_47.n15 a_44_47.t7 25.846
R65 a_44_47.n10 a_44_47.t0 25.846
R66 a_44_47.n13 a_44_47.t9 25.846
R67 a_44_47.n6 a_44_47.n4 25.6
R68 a_44_47.n9 a_44_47.n6 25.6
R69 a_44_47.n17 a_44_47.n16 18.626
R70 a_44_47.n3 a_44_47.n2 13.145
R71 a_44_47.n8 a_44_47.n7 13.145
R72 a_44_47.n12 a_44_47.n11 5.393
R73 VGND.n2 VGND.t2 192.675
R74 VGND.n10 VGND.t11 191.969
R75 VGND.n34 VGND.n33 107.239
R76 VGND.n1 VGND.n0 106.463
R77 VGND.n6 VGND.n5 106.463
R78 VGND.n29 VGND.n28 106.463
R79 VGND.n19 VGND.n18 92.5
R80 VGND.n23 VGND.n22 92.5
R81 VGND.n28 VGND.t10 33.23
R82 VGND.n18 VGND.t0 29.538
R83 VGND.n22 VGND.t1 25.846
R84 VGND.n0 VGND.t4 25.846
R85 VGND.n0 VGND.t5 25.846
R86 VGND.n5 VGND.t3 25.846
R87 VGND.n5 VGND.t6 25.846
R88 VGND.n33 VGND.t8 25.846
R89 VGND.n33 VGND.t7 25.846
R90 VGND.n28 VGND.t9 24.923
R91 VGND.n4 VGND.n3 4.65
R92 VGND.n7 VGND.n6 4.65
R93 VGND.n9 VGND.n8 4.65
R94 VGND.n11 VGND.n10 4.65
R95 VGND.n13 VGND.n12 4.65
R96 VGND.n15 VGND.n14 4.65
R97 VGND.n17 VGND.n16 4.65
R98 VGND.n21 VGND.n20 4.65
R99 VGND.n25 VGND.n24 4.65
R100 VGND.n27 VGND.n26 4.65
R101 VGND.n30 VGND.n29 4.65
R102 VGND.n32 VGND.n31 4.65
R103 VGND.n35 VGND.n34 4.067
R104 VGND.n2 VGND.n1 3.773
R105 VGND.n20 VGND.n19 2.777
R106 VGND.n24 VGND.n23 1.328
R107 VGND.n4 VGND.n2 0.261
R108 VGND.n35 VGND.n32 0.134
R109 VGND VGND.n35 0.127
R110 VGND.n7 VGND.n4 0.119
R111 VGND.n9 VGND.n7 0.119
R112 VGND.n11 VGND.n9 0.119
R113 VGND.n13 VGND.n11 0.119
R114 VGND.n15 VGND.n13 0.119
R115 VGND.n17 VGND.n15 0.119
R116 VGND.n21 VGND.n17 0.119
R117 VGND.n25 VGND.n21 0.119
R118 VGND.n27 VGND.n25 0.119
R119 VGND.n30 VGND.n27 0.119
R120 VGND.n32 VGND.n30 0.119
R121 VNB VNB.t9 6513.25
R122 VNB.t1 VNB.t13 4738.46
R123 VNB.t3 VNB.t2 4690.11
R124 VNB.t11 VNB.t3 2345.05
R125 VNB.t12 VNB.t11 2248.35
R126 VNB.t2 VNB.t0 2103.3
R127 VNB.t6 VNB.t4 2079.12
R128 VNB.t7 VNB.t6 2079.12
R129 VNB.t5 VNB.t7 2079.12
R130 VNB.t8 VNB.t5 2079.12
R131 VNB.t13 VNB.t8 2079.12
R132 VNB.t0 VNB.t1 2079.12
R133 VNB.t10 VNB.t12 2079.12
R134 VNB.t9 VNB.t10 2079.12
R135 B1.n0 B1.t3 213.686
R136 B1.n2 B1.t2 213.686
R137 B1.n3 B1.t1 176.114
R138 B1.n0 B1.t0 167.957
R139 B1.n1 B1 83.225
R140 B1.n4 B1.n3 76
R141 B1.n2 B1.n1 54.873
R142 B1.n3 B1.n2 15.572
R143 B1.n4 B1 12.387
R144 B1.n1 B1.n0 8.898
R145 B1 B1.n4 6.606
R146 X.n2 X.n1 205.8
R147 X.n5 X.n3 163.157
R148 X.n2 X.n0 161.768
R149 X.n5 X.n4 112.71
R150 X X.n2 31.054
R151 X.n0 X.t1 27.58
R152 X.n0 X.t2 27.58
R153 X.n1 X.t3 27.58
R154 X.n1 X.t0 27.58
R155 X.n3 X.t7 25.846
R156 X.n3 X.t5 25.846
R157 X.n4 X.t4 25.846
R158 X.n4 X.t6 25.846
R159 X X.n5 23.056
R160 A1.n0 A1.t1 208.866
R161 A1.n2 A1.t0 208.866
R162 A1.n2 A1.t2 145.449
R163 A1.n1 A1.t3 139.779
R164 A1.n0 A1 90.29
R165 A1.n4 A1.n3 76
R166 A1.n3 A1.n1 30.479
R167 A1.n3 A1.n2 24.808
R168 A1.n4 A1 19.52
R169 A1 A1.n4 9.92
R170 A1.n1 A1.n0 5.67
R171 a_477_297.t3 a_477_297.n3 241.706
R172 a_477_297.n1 a_477_297.n0 200.942
R173 a_477_297.n1 a_477_297.t4 177.652
R174 a_477_297.n3 a_477_297.n2 143.026
R175 a_477_297.n3 a_477_297.n1 52.402
R176 a_477_297.n2 a_477_297.t2 51.22
R177 a_477_297.n2 a_477_297.t5 50.235
R178 a_477_297.n0 a_477_297.t1 27.58
R179 a_477_297.n0 a_477_297.t0 27.58
R180 VPWR.n12 VPWR.t4 575.999
R181 VPWR.n1 VPWR.n0 310.73
R182 VPWR.n4 VPWR.t1 195.999
R183 VPWR.n8 VPWR.n7 165.273
R184 VPWR.n3 VPWR.n2 164.492
R185 VPWR.n2 VPWR.t2 27.58
R186 VPWR.n2 VPWR.t3 27.58
R187 VPWR.n7 VPWR.t0 27.58
R188 VPWR.n7 VPWR.t5 27.58
R189 VPWR.n0 VPWR.t6 27.58
R190 VPWR.n0 VPWR.t7 27.58
R191 VPWR.n6 VPWR.n5 4.65
R192 VPWR.n9 VPWR.n8 4.65
R193 VPWR.n11 VPWR.n10 4.65
R194 VPWR.n13 VPWR.n12 4.65
R195 VPWR.n15 VPWR.n14 4.65
R196 VPWR.n16 VPWR.n1 4.097
R197 VPWR.n4 VPWR.n3 3.773
R198 VPWR VPWR.n16 0.963
R199 VPWR.n6 VPWR.n4 0.261
R200 VPWR.n16 VPWR.n15 0.135
R201 VPWR.n9 VPWR.n6 0.119
R202 VPWR.n11 VPWR.n9 0.119
R203 VPWR.n13 VPWR.n11 0.119
R204 VPWR.n15 VPWR.n13 0.119
R205 D1.n0 D1.t1 212.079
R206 D1.n2 D1.t2 212.079
R207 D1.n0 D1.t3 151.81
R208 D1.n1 D1.t0 139.779
R209 D1.n3 D1.n2 108.133
R210 D1.n1 D1.n0 52.581
R211 D1.n3 D1 12.8
R212 D1.n2 D1.n1 10.224
R213 D1 D1.n3 2.47
R214 A2.n0 A2.t3 212.079
R215 A2.n2 A2.t2 212.079
R216 A2.n0 A2.t1 139.779
R217 A2.n2 A2.t0 139.779
R218 A2.n1 A2 91.04
R219 A2.n3 A2.n2 85.493
R220 A2.n2 A2.n1 40.166
R221 A2 A2.n3 23.36
R222 A2.n1 A2.n0 22.639
R223 A2.n3 A2 6.72
R224 a_770_47.n1 a_770_47.n0 303.76
R225 a_770_47.n0 a_770_47.t2 25.846
R226 a_770_47.n0 a_770_47.t3 25.846
R227 a_770_47.n1 a_770_47.t0 25.846
R228 a_770_47.t1 a_770_47.n1 25.846
C0 X VGND 0.33fF
C1 VPWR VGND 0.17fF
C2 VPWR X 0.55fF
C3 VPWR VPB 0.15fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__a2111oi_0.ext - technology: sky130A

.subckt sky130_fd_sc_hd__a2111oi_0 A2 A1 B1 C1 Y D1 VPWR VGND VNB VPB
X0 Y.t4 B1.t0 VGND.t3 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1 VPWR.t1 A1.t0 a_313_369.t2 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X2 a_427_47.t1 A1.t1 Y.t0 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3 a_241_369.t0 C1.t0 a_169_369.t1 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X4 VGND.t1 C1.t1 Y.t2 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 VGND.t0 A2.t0 a_427_47.t0 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 a_169_369.t0 D1.t0 Y.t1 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X7 Y.t3 D1.t1 VGND.t2 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 a_313_369.t1 B1.t1 a_241_369.t1 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X9 a_313_369.t0 A2.t1 VPWR.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
R0 B1.n0 B1.t1 271.526
R1 B1.n0 B1.t0 218.735
R2 B1.n1 B1.n0 76
R3 B1.n1 B1 8.228
R4 B1 B1.n1 4.205
R5 VGND.n7 VGND.t2 157.239
R6 VGND.n0 VGND.t0 149.986
R7 VGND.n2 VGND.n1 106.463
R8 VGND.n1 VGND.t3 51.428
R9 VGND.n1 VGND.t1 48.571
R10 VGND.n8 VGND.n7 8.791
R11 VGND.n4 VGND.n3 4.65
R12 VGND.n6 VGND.n5 4.65
R13 VGND.n3 VGND.n2 4.517
R14 VGND.n4 VGND.n0 0.182
R15 VGND.n6 VGND.n4 0.119
R16 VGND.n8 VGND.n6 0.119
R17 VGND VGND.n8 0.022
R18 Y.n0 Y.t1 199.097
R19 Y.n4 Y.n3 142.255
R20 Y.n4 Y.n2 102.288
R21 Y.n3 Y.t0 40
R22 Y.n3 Y.t4 40
R23 Y.n2 Y.t2 40
R24 Y.n2 Y.t3 40
R25 Y.n1 Y.n0 6.967
R26 Y Y.n4 6.28
R27 Y Y.n1 2.844
R28 Y.n0 Y 2.04
R29 Y.n1 Y 1.204
R30 VNB VNB.t3 8012.74
R31 VNB.t2 VNB.t4 3235.29
R32 VNB.t4 VNB.t0 2782.35
R33 VNB.t3 VNB.t2 2782.35
R34 VNB.t0 VNB.t1 2329.41
R35 A1.n1 A1.t1 208.815
R36 A1.n1 A1.t0 200.216
R37 A1.n2 A1.n1 59.619
R38 A1.n0 A1 14.459
R39 A1.n0 A1 1.719
R40 A1.n2 A1.n0 1.505
R41 A1 A1.n2 0.238
R42 a_313_369.t0 a_313_369.n0 402.009
R43 a_313_369.n0 a_313_369.t2 43.093
R44 a_313_369.n0 a_313_369.t1 43.093
R45 VPWR VPWR.n0 311.009
R46 VPWR.n0 VPWR.t1 64.64
R47 VPWR.n0 VPWR.t0 52.328
R48 VPB VPB.t1 369.937
R49 VPB.t4 VPB.t0 313.707
R50 VPB.t3 VPB.t4 254.517
R51 VPB.t2 VPB.t3 213.084
R52 VPB.t1 VPB.t2 213.084
R53 a_427_47.t0 a_427_47.t1 60
R54 C1.n0 C1.t0 270.357
R55 C1.n0 C1.t1 221.865
R56 C1.n1 C1.n0 76
R57 C1 C1.n1 7.783
R58 C1.n1 C1 3.978
R59 a_169_369.t0 a_169_369.t1 64.64
R60 a_241_369.t0 a_241_369.t1 64.64
R61 A2.n1 A2.t0 285.183
R62 A2.n0 A2.t1 285.067
R63 A2 A2.n0 77.882
R64 A2.n2 A2.n1 76
R65 A2 A2.n2 10.917
R66 A2.n2 A2 1.882
R67 D1.n1 D1.t0 286.343
R68 D1.n2 D1.t1 182.98
R69 D1.n3 D1.n2 76
R70 D1.n1 D1.n0 76
R71 D1.n2 D1.n1 68.729
R72 D1.n0 D1 7.68
R73 D1.n3 D1 6.4
R74 D1 D1.n3 6.034
R75 D1.n0 D1 4.754
C0 A1 A2 0.29fF
C1 B1 A1 0.16fF
C2 C1 Y 0.27fF
C3 D1 Y 0.13fF
C4 Y VGND 0.30fF
C5 C1 B1 0.19fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__a2111oi_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__a2111oi_1 B1 D1 C1 Y A2 A1 VPWR VGND VNB VPB
X0 a_316_297.t1 C1.t0 a_217_297.t0 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 Y.t0 D1.t0 VGND.t0 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 VGND.t3 C1.t1 Y.t4 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 a_420_297.t0 B1.t0 a_316_297.t0 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 VPWR.t1 A1.t0 a_420_297.t2 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 VGND.t1 A2.t0 a_568_47.t0 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 Y.t3 B1.t1 VGND.t2 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 a_420_297.t1 A2.t1 VPWR.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 a_217_297.t1 D1.t1 Y.t1 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 a_568_47.t1 A1.t1 Y.t2 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
R0 C1.n0 C1.t0 228.612
R1 C1.n0 C1.t1 161.287
R2 C1.n1 C1.n0 76
R3 C1.n1 C1 10.889
R4 C1 C1.n1 2.101
R5 a_217_297.t0 a_217_297.t1 67.965
R6 a_316_297.t0 a_316_297.t1 72.89
R7 VPB VPB.t4 511.993
R8 VPB.t2 VPB.t1 432.087
R9 VPB.t3 VPB.t2 307.788
R10 VPB.t4 VPB.t3 292.99
R11 VPB.t1 VPB.t0 251.557
R12 D1.n0 D1.t1 238.589
R13 D1.n0 D1.t0 166.289
R14 D1.n1 D1.n0 76
R15 D1.n1 D1 8.106
R16 D1 D1.n1 1.564
R17 VGND.n5 VGND.t0 183.743
R18 VGND.n2 VGND.t1 148.94
R19 VGND.n1 VGND.n0 106.851
R20 VGND.n0 VGND.t2 43.384
R21 VGND.n0 VGND.t3 24.923
R22 VGND.n4 VGND.n3 4.65
R23 VGND.n7 VGND.n6 4.65
R24 VGND.n6 VGND.n5 4.517
R25 VGND.n2 VGND.n1 3.691
R26 VGND.n4 VGND.n2 0.148
R27 VGND.n7 VGND.n4 0.119
R28 VGND.n8 VGND.n7 0.119
R29 VGND VGND.n8 0.022
R30 Y.n5 Y.n4 292.5
R31 Y.n6 Y.n5 146.251
R32 Y.n2 Y.n0 106.864
R33 Y.n5 Y.t1 96.53
R34 Y.n0 Y.t2 80.307
R35 Y.n2 Y.n1 51.426
R36 Y.n1 Y.t4 41.105
R37 Y.n3 Y.n2 36.622
R38 Y.n1 Y.t0 29.967
R39 Y.n0 Y.t3 28.615
R40 Y Y.n3 10.472
R41 Y.n6 Y 8.423
R42 Y.n4 Y 5.818
R43 Y.n4 Y 5.485
R44 Y Y.n6 2.826
R45 Y.n3 Y 0.831
R46 VNB.t0 VNB 8495.67
R47 VNB VNB.n0 4400
R48 VNB.n0 VNB.t2 3408.79
R49 VNB.t4 VNB.t0 2586.81
R50 VNB.t3 VNB.t4 2514.28
R51 VNB.t2 VNB.t1 1982.42
R52 VNB.n0 VNB.t3 169.23
R53 B1.n0 B1.t0 238.248
R54 B1.n0 B1.t1 161.21
R55 B1.n1 B1.n0 76
R56 B1 B1.n1 11.403
R57 B1.n1 B1 2.133
R58 a_420_297.n0 a_420_297.t1 406.123
R59 a_420_297.t0 a_420_297.n0 86.68
R60 a_420_297.n0 a_420_297.t2 27.58
R61 A1.n0 A1.t0 327.612
R62 A1.n0 A1.t1 154.551
R63 A1 A1.n0 81.53
R64 VPWR VPWR.n0 168.167
R65 VPWR.n0 VPWR.t0 27.58
R66 VPWR.n0 VPWR.t1 26.595
R67 A2.n0 A2.t1 235.47
R68 A2.n0 A2.t0 157.783
R69 A2.n1 A2.n0 76
R70 A2 A2.n1 30.205
R71 A2.n1 A2 4.977
R72 a_568_47.t0 a_568_47.t1 48
C0 A2 A1 0.10fF
C1 B1 A1 0.10fF
C2 C1 B1 0.29fF
C3 Y VGND 0.40fF
C4 A2 VGND 0.14fF
C5 Y D1 0.23fF
C6 D1 C1 0.24fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__a2111oi_2.ext - technology: sky130A

.subckt sky130_fd_sc_hd__a2111oi_2 D1 C1 A2 A1 Y B1 VGND VPWR VNB VPB
X0 a_467_297.t2 B1.t0 a_28_297.t3 VPB.t6 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_287_297.t0 D1.t0 Y.t4 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 VPWR.t1 A2.t0 a_467_297.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 a_923_47.t0 A2.t1 VGND.t4 VNB.t6 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 Y.t8 B1.t1 VGND.t7 VNB.t8 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 a_28_297.t2 B1.t2 a_467_297.t1 VPB.t5 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 VGND.t2 C1.t0 Y.t5 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 a_28_297.t0 C1.t1 a_287_297.t1 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 Y.t9 A1.t0 a_923_47.t1 VNB.t9 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 VGND.t5 A2.t2 a_684_47.t0 VNB.t5 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 Y.t3 D1.t1 VGND.t1 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 VGND.t6 B1.t3 Y.t7 VNB.t7 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 Y.t1 D1.t2 a_115_297.t0 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13 a_467_297.t4 A1.t1 VPWR.t2 VPB.t8 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14 VGND.t0 D1.t3 Y.t2 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X15 Y.t6 C1.t2 VGND.t3 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X16 VPWR.t3 A1.t2 a_467_297.t5 VPB.t9 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17 a_115_297.t1 C1.t3 a_28_297.t1 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X18 a_467_297.t3 A2.t3 VPWR.t0 VPB.t7 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X19 a_684_47.t1 A1.t3 Y.t0 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
R0 B1.n2 B1.t0 225.224
R1 B1.n0 B1.t2 212.079
R2 B1.n0 B1.t1 172.642
R3 B1.n1 B1.t3 139.779
R4 B1 B1.n0 88.8
R5 B1 B1.n2 80.963
R6 B1.n2 B1.n1 3.651
R7 a_28_297.n0 a_28_297.t2 597.134
R8 a_28_297.n1 a_28_297.n0 292.5
R9 a_28_297.n0 a_28_297.t1 281.231
R10 a_28_297.n1 a_28_297.t3 35.46
R11 a_28_297.t0 a_28_297.n1 27.58
R12 a_467_297.n3 a_467_297.n2 365.164
R13 a_467_297.n1 a_467_297.t4 227.054
R14 a_467_297.n2 a_467_297.t5 172.358
R15 a_467_297.n1 a_467_297.n0 149.04
R16 a_467_297.n2 a_467_297.n1 45.389
R17 a_467_297.n0 a_467_297.t0 27.58
R18 a_467_297.n0 a_467_297.t3 27.58
R19 a_467_297.n3 a_467_297.t1 27.58
R20 a_467_297.t2 a_467_297.n3 27.58
R21 VPB.t5 VPB.t9 562.305
R22 VPB.t0 VPB.t8 278.193
R23 VPB.t3 VPB.t6 278.193
R24 VPB.t7 VPB.t0 254.517
R25 VPB.t9 VPB.t7 254.517
R26 VPB.t6 VPB.t5 254.517
R27 VPB.t1 VPB.t3 254.517
R28 VPB.t2 VPB.t1 254.517
R29 VPB.t4 VPB.t2 254.517
R30 VPB VPB.t4 210.124
R31 D1.n0 D1.t0 212.079
R32 D1.n1 D1.t2 212.079
R33 D1.n0 D1.t3 139.779
R34 D1.n1 D1.t1 139.779
R35 D1 D1.n2 34.352
R36 D1.n2 D1.n0 33.695
R37 D1.n2 D1.n1 18.714
R38 Y Y.n0 415.563
R39 Y.n6 Y.t9 258.277
R40 Y.n3 Y.t5 113.332
R41 Y.n8 Y.n1 92.5
R42 Y.n3 Y.n2 50.428
R43 Y.n5 Y.n4 49.353
R44 Y Y.n8 38.025
R45 Y.n5 Y.n3 37.286
R46 Y.n7 Y.n5 37.286
R47 Y.n4 Y.t7 31.384
R48 Y.n4 Y.t6 28.615
R49 Y.n0 Y.t4 27.58
R50 Y.n0 Y.t1 27.58
R51 Y.n1 Y.t0 25.846
R52 Y.n1 Y.t8 25.846
R53 Y.n2 Y.t2 25.846
R54 Y.n2 Y.t3 25.846
R55 Y.n7 Y.n6 8.386
R56 Y.n8 Y.n7 0.441
R57 a_287_297.t0 a_287_297.t1 55.16
R58 A2.n0 A2.t0 212.079
R59 A2.n2 A2.t3 212.079
R60 A2.n2 A2.t2 141.77
R61 A2.n1 A2.t1 141.05
R62 A2 A2.n1 87.569
R63 A2 A2.n3 81.169
R64 A2.n3 A2.n2 15.826
R65 A2.n1 A2.n0 2.877
R66 VPWR.n2 VPWR.n0 309.943
R67 VPWR.n2 VPWR.n1 309.752
R68 VPWR.n0 VPWR.t2 31.52
R69 VPWR.n0 VPWR.t1 31.52
R70 VPWR.n1 VPWR.t0 27.58
R71 VPWR.n1 VPWR.t3 27.58
R72 VPWR VPWR.n2 1.063
R73 VGND.n3 VGND.n0 110.262
R74 VGND.n2 VGND.n1 106.463
R75 VGND.n7 VGND.n6 106.463
R76 VGND.n12 VGND.n11 106.463
R77 VGND.n1 VGND.t7 38.769
R78 VGND.n6 VGND.t3 36
R79 VGND.n6 VGND.t0 36
R80 VGND.n1 VGND.t6 33.23
R81 VGND.n0 VGND.t4 32.307
R82 VGND.n0 VGND.t5 31.384
R83 VGND.n11 VGND.t1 25.846
R84 VGND.n11 VGND.t2 25.846
R85 VGND.n5 VGND.n4 4.65
R86 VGND.n8 VGND.n7 4.65
R87 VGND.n10 VGND.n9 4.65
R88 VGND.n13 VGND.n12 3.989
R89 VGND.n3 VGND.n2 3.706
R90 VGND.n5 VGND.n3 0.148
R91 VGND.n13 VGND.n10 0.136
R92 VGND VGND.n13 0.125
R93 VGND.n8 VGND.n5 0.119
R94 VGND.n10 VGND.n8 0.119
R95 a_923_47.t0 a_923_47.t1 51.692
R96 VNB VNB.t3 6223.14
R97 VNB.t0 VNB.t5 3384.61
R98 VNB.t7 VNB.t8 2610.99
R99 VNB.t1 VNB.t4 2610.99
R100 VNB.t5 VNB.t6 2393.41
R101 VNB.t4 VNB.t7 2296.7
R102 VNB.t6 VNB.t9 2079.12
R103 VNB.t8 VNB.t0 2079.12
R104 VNB.t2 VNB.t1 2079.12
R105 VNB.t3 VNB.t2 2079.12
R106 C1.n0 C1.t1 236.179
R107 C1.n1 C1.t3 229.752
R108 C1.n0 C1.t2 163.879
R109 C1.n1 C1.t0 157.452
R110 C1 C1.n1 149.795
R111 C1 C1.n0 101.654
R112 A1.n0 A1.t1 236.179
R113 A1.n1 A1.t2 229.95
R114 A1.n0 A1.t0 163.879
R115 A1.n1 A1.t3 157.65
R116 A1 A1.n0 148.509
R117 A1 A1.n1 102.601
R118 a_684_47.t0 a_684_47.t1 101.538
R119 a_115_297.t0 a_115_297.t1 55.16
C0 A2 Y 0.16fF
C1 A1 Y 0.23fF
C2 B1 Y 0.36fF
C3 VPWR VGND 0.11fF
C4 Y VGND 0.81fF
C5 D1 Y 0.11fF
C6 C1 Y 0.37fF
C7 VPB VPWR 0.10fF
C8 C1 D1 0.34fF
C9 A1 A2 0.37fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__a2111oi_4.ext - technology: sky130A

.subckt sky130_fd_sc_hd__a2111oi_4 D1 C1 B1 A2 A1 Y VGND VPWR VNB VPB
X0 Y.t3 D1.t0 VGND.t7 VNB.t7 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 a_455_297.t7 B1.t0 a_821_297.t8 VPB.t16 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 a_28_297.t3 D1.t1 Y.t5 VPB.t7 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 a_821_297.t1 A2.t0 VPWR.t3 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 a_28_297.t6 C1.t0 a_455_297.t2 VPB.t10 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 a_455_297.t3 C1.t1 a_28_297.t7 VPB.t11 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 VGND.t6 D1.t2 Y.t2 VNB.t6 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 VGND.t13 B1.t1 Y.t15 VNB.t15 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 VPWR.t2 A2.t1 a_821_297.t2 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 Y.t4 D1.t3 a_28_297.t2 VPB.t6 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 Y.t12 C1.t2 VGND.t12 VNB.t12 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 VGND.t5 D1.t4 Y.t1 VNB.t5 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 Y.t0 D1.t5 VGND.t4 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 a_821_297.t7 B1.t2 a_455_297.t6 VPB.t15 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14 Y.t16 B1.t3 VGND.t14 VNB.t16 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X15 Y.t7 D1.t6 a_28_297.t1 VPB.t5 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16 Y.t9 C1.t3 VGND.t9 VNB.t9 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X17 a_1205_47.t3 A2.t2 VGND.t1 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X18 a_28_297.t4 C1.t4 a_455_297.t0 VPB.t8 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X19 Y.t17 B1.t4 VGND.t15 VNB.t17 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X20 a_1205_47.t2 A2.t3 VGND.t2 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X21 a_821_297.t3 A2.t4 VPWR.t1 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X22 VGND.t10 C1.t5 Y.t10 VNB.t10 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X23 Y.t13 A1.t0 a_1205_47.t4 VNB.t13 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X24 VGND.t11 C1.t6 Y.t11 VNB.t11 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X25 VPWR.t4 A1.t1 a_821_297.t4 VPB.t12 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X26 Y.t14 A1.t2 a_1205_47.t5 VNB.t14 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X27 a_1205_47.t6 A1.t3 Y.t18 VNB.t18 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X28 a_28_297.t0 D1.t7 Y.t6 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X29 VGND.t3 A2.t5 a_1205_47.t1 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X30 a_455_297.t5 B1.t5 a_821_297.t6 VPB.t14 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X31 a_821_297.t9 A1.t4 VPWR.t5 VPB.t17 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X32 a_1205_47.t7 A1.t5 Y.t19 VNB.t19 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X33 VGND.t0 A2.t6 a_1205_47.t0 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X34 VPWR.t6 A1.t6 a_821_297.t10 VPB.t18 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X35 a_821_297.t11 A1.t7 VPWR.t7 VPB.t19 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X36 VPWR.t0 A2.t7 a_821_297.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X37 a_455_297.t1 C1.t7 a_28_297.t5 VPB.t9 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X38 a_821_297.t5 B1.t6 a_455_297.t4 VPB.t13 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X39 VGND.t8 B1.t7 Y.t8 VNB.t8 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
R0 D1.n6 D1.t3 213.539
R1 D1.n1 D1.t6 212.079
R2 D1.n0 D1.t7 212.079
R3 D1.n3 D1.t1 212.079
R4 D1.n1 D1.t0 139.779
R5 D1.n0 D1.t2 139.779
R6 D1.n3 D1.t4 139.779
R7 D1.n6 D1.t5 139.779
R8 D1.n5 D1.n4 76
R9 D1.n8 D1.n7 76
R10 D1.n5 D1.n2 49.404
R11 D1.n2 D1.n0 34.276
R12 D1.n7 D1.n6 24.83
R13 D1.n2 D1.n1 17.256
R14 D1.n8 D1.n5 17.066
R15 D1.n4 D1.n3 13.145
R16 D1 D1.n8 2.509
R17 VGND.n44 VGND.t4 192.177
R18 VGND.n14 VGND.t8 191.969
R19 VGND.n3 VGND.n0 109.724
R20 VGND.n2 VGND.n1 106.463
R21 VGND.n19 VGND.n18 106.463
R22 VGND.n24 VGND.n23 106.463
R23 VGND.n29 VGND.n28 106.463
R24 VGND.n40 VGND.n39 106.463
R25 VGND.n34 VGND.n33 92.5
R26 VGND.n33 VGND.t6 40.615
R27 VGND.n23 VGND.t10 36.923
R28 VGND.n23 VGND.t15 35.076
R29 VGND.n33 VGND.t9 25.846
R30 VGND.n0 VGND.t1 25.846
R31 VGND.n0 VGND.t3 25.846
R32 VGND.n1 VGND.t2 25.846
R33 VGND.n1 VGND.t0 25.846
R34 VGND.n18 VGND.t14 25.846
R35 VGND.n18 VGND.t13 25.846
R36 VGND.n28 VGND.t12 25.846
R37 VGND.n28 VGND.t11 25.846
R38 VGND.n39 VGND.t7 25.846
R39 VGND.n39 VGND.t5 25.846
R40 VGND.n45 VGND.n44 4.65
R41 VGND.n5 VGND.n4 4.65
R42 VGND.n7 VGND.n6 4.65
R43 VGND.n9 VGND.n8 4.65
R44 VGND.n11 VGND.n10 4.65
R45 VGND.n13 VGND.n12 4.65
R46 VGND.n15 VGND.n14 4.65
R47 VGND.n17 VGND.n16 4.65
R48 VGND.n20 VGND.n19 4.65
R49 VGND.n22 VGND.n21 4.65
R50 VGND.n25 VGND.n24 4.65
R51 VGND.n27 VGND.n26 4.65
R52 VGND.n30 VGND.n29 4.65
R53 VGND.n32 VGND.n31 4.65
R54 VGND.n36 VGND.n35 4.65
R55 VGND.n38 VGND.n37 4.65
R56 VGND.n41 VGND.n40 4.65
R57 VGND.n43 VGND.n42 4.65
R58 VGND.n3 VGND.n2 3.94
R59 VGND.n5 VGND.n3 0.261
R60 VGND.n35 VGND.n34 0.12
R61 VGND.n7 VGND.n5 0.119
R62 VGND.n9 VGND.n7 0.119
R63 VGND.n11 VGND.n9 0.119
R64 VGND.n13 VGND.n11 0.119
R65 VGND.n15 VGND.n13 0.119
R66 VGND.n17 VGND.n15 0.119
R67 VGND.n20 VGND.n17 0.119
R68 VGND.n22 VGND.n20 0.119
R69 VGND.n25 VGND.n22 0.119
R70 VGND.n27 VGND.n25 0.119
R71 VGND.n30 VGND.n27 0.119
R72 VGND.n32 VGND.n30 0.119
R73 VGND.n36 VGND.n32 0.119
R74 VGND.n38 VGND.n36 0.119
R75 VGND.n41 VGND.n38 0.119
R76 VGND.n43 VGND.n41 0.119
R77 VGND.n45 VGND.n43 0.119
R78 VGND VGND.n45 0.02
R79 Y.n2 Y.n0 184.734
R80 Y.n5 Y.n3 157.252
R81 Y.n2 Y.n1 151.802
R82 Y.n7 Y.n5 102.878
R83 Y.n5 Y.n4 92.5
R84 Y.n7 Y.n6 92.5
R85 Y.n9 Y.n8 92.5
R86 Y.n11 Y.n10 92.5
R87 Y.n13 Y.n12 92.5
R88 Y.n15 Y.n14 92.5
R89 Y.n17 Y.n16 92.5
R90 Y Y.n2 73.845
R91 Y.n15 Y.n13 63.838
R92 Y.n11 Y.n9 62.083
R93 Y.n9 Y.n7 57.815
R94 Y.n13 Y.n11 57.815
R95 Y.n17 Y.n15 57.621
R96 Y Y.n17 30.261
R97 Y.n1 Y.t5 27.58
R98 Y.n1 Y.t4 27.58
R99 Y.n0 Y.t6 27.58
R100 Y.n0 Y.t7 27.58
R101 Y.n14 Y.t2 25.846
R102 Y.n14 Y.t3 25.846
R103 Y.n12 Y.t11 25.846
R104 Y.n12 Y.t9 25.846
R105 Y.n10 Y.t10 25.846
R106 Y.n10 Y.t12 25.846
R107 Y.n8 Y.t15 25.846
R108 Y.n8 Y.t17 25.846
R109 Y.n6 Y.t8 25.846
R110 Y.n6 Y.t16 25.846
R111 Y.n4 Y.t19 25.846
R112 Y.n4 Y.t14 25.846
R113 Y.n3 Y.t18 25.846
R114 Y.n3 Y.t13 25.846
R115 Y.n16 Y.t1 24.923
R116 Y.n16 Y.t0 24.923
R117 VNB VNB.t4 6150.61
R118 VNB.t8 VNB.t14 4738.46
R119 VNB.t10 VNB.t17 2610.99
R120 VNB.t18 VNB.t0 2538.46
R121 VNB.t6 VNB.t9 2465.93
R122 VNB.t3 VNB.t1 2079.12
R123 VNB.t2 VNB.t3 2079.12
R124 VNB.t0 VNB.t2 2079.12
R125 VNB.t13 VNB.t18 2079.12
R126 VNB.t19 VNB.t13 2079.12
R127 VNB.t14 VNB.t19 2079.12
R128 VNB.t16 VNB.t8 2079.12
R129 VNB.t15 VNB.t16 2079.12
R130 VNB.t17 VNB.t15 2079.12
R131 VNB.t12 VNB.t10 2079.12
R132 VNB.t11 VNB.t12 2079.12
R133 VNB.t9 VNB.t11 2079.12
R134 VNB.t7 VNB.t6 2079.12
R135 VNB.t5 VNB.t7 2079.12
R136 VNB.t4 VNB.t5 2030.77
R137 B1.n1 B1.t6 248.594
R138 B1.n2 B1.t5 212.079
R139 B1.n6 B1.t2 212.079
R140 B1.n10 B1.t0 212.079
R141 B1.n13 B1.t4 141.239
R142 B1.n9 B1.t1 139.779
R143 B1.n5 B1.t3 139.779
R144 B1.n0 B1.t7 139.779
R145 B1.n4 B1.n1 93.066
R146 B1 B1.n13 84.533
R147 B1.n4 B1.n3 76
R148 B1.n8 B1.n7 76
R149 B1.n12 B1.n11 76
R150 B1.n3 B1.n2 23.369
R151 B1.n8 B1.n4 17.066
R152 B1.n12 B1.n8 17.066
R153 B1.n6 B1.n5 14.606
R154 B1.n1 B1.n0 11.684
R155 B1.n11 B1.n9 11.684
R156 B1.n7 B1.n6 10.224
R157 B1 B1.n12 8.533
R158 B1.n11 B1.n10 2.921
R159 a_821_297.n2 a_821_297.t8 228.942
R160 a_821_297.n8 a_821_297.t1 226.922
R161 a_821_297.n6 a_821_297.n5 160.496
R162 a_821_297.n9 a_821_297.n8 158.661
R163 a_821_297.n7 a_821_297.n0 151.387
R164 a_821_297.n2 a_821_297.n1 150.103
R165 a_821_297.n4 a_821_297.n3 136.066
R166 a_821_297.n4 a_821_297.n2 83.359
R167 a_821_297.n6 a_821_297.n4 77.553
R168 a_821_297.n7 a_821_297.n6 51.416
R169 a_821_297.n0 a_821_297.t2 46.371
R170 a_821_297.n8 a_821_297.n7 38.981
R171 a_821_297.t0 a_821_297.n9 37.458
R172 a_821_297.n9 a_821_297.t3 35.427
R173 a_821_297.n0 a_821_297.t9 32.273
R174 a_821_297.n3 a_821_297.t5 29.55
R175 a_821_297.n3 a_821_297.t4 27.58
R176 a_821_297.n1 a_821_297.t6 27.58
R177 a_821_297.n1 a_821_297.t7 27.58
R178 a_821_297.n5 a_821_297.t10 27.58
R179 a_821_297.n5 a_821_297.t11 27.58
R180 a_455_297.n3 a_455_297.n1 184.882
R181 a_455_297.n4 a_455_297.n0 184.734
R182 a_455_297.n3 a_455_297.n2 152.43
R183 a_455_297.n5 a_455_297.n4 152.429
R184 a_455_297.n4 a_455_297.n3 75.828
R185 a_455_297.n2 a_455_297.t0 27.58
R186 a_455_297.n2 a_455_297.t3 27.58
R187 a_455_297.n1 a_455_297.t2 27.58
R188 a_455_297.n1 a_455_297.t1 27.58
R189 a_455_297.n0 a_455_297.t4 27.58
R190 a_455_297.n0 a_455_297.t5 27.58
R191 a_455_297.t6 a_455_297.n5 27.58
R192 a_455_297.n5 a_455_297.t7 27.58
R193 VPB.t8 VPB.t16 562.305
R194 VPB.t17 VPB.t2 325.545
R195 VPB.t3 VPB.t0 307.788
R196 VPB.t18 VPB.t17 266.355
R197 VPB.t13 VPB.t12 260.436
R198 VPB.t0 VPB.t1 254.517
R199 VPB.t2 VPB.t3 254.517
R200 VPB.t19 VPB.t18 254.517
R201 VPB.t12 VPB.t19 254.517
R202 VPB.t14 VPB.t13 254.517
R203 VPB.t15 VPB.t14 254.517
R204 VPB.t16 VPB.t15 254.517
R205 VPB.t11 VPB.t8 254.517
R206 VPB.t10 VPB.t11 254.517
R207 VPB.t9 VPB.t10 254.517
R208 VPB.t4 VPB.t9 254.517
R209 VPB.t5 VPB.t4 254.517
R210 VPB.t7 VPB.t5 254.517
R211 VPB.t6 VPB.t7 254.517
R212 VPB VPB.t6 195.327
R213 a_28_297.n4 a_28_297.t2 229.927
R214 a_28_297.n1 a_28_297.t4 228.942
R215 a_28_297.n5 a_28_297.n4 150.104
R216 a_28_297.n1 a_28_297.n0 150.103
R217 a_28_297.n3 a_28_297.n2 150.103
R218 a_28_297.n3 a_28_297.n1 57.936
R219 a_28_297.n4 a_28_297.n3 57.936
R220 a_28_297.n2 a_28_297.t5 27.58
R221 a_28_297.n2 a_28_297.t0 27.58
R222 a_28_297.n0 a_28_297.t7 27.58
R223 a_28_297.n0 a_28_297.t6 27.58
R224 a_28_297.n5 a_28_297.t1 27.58
R225 a_28_297.t3 a_28_297.n5 27.58
R226 A2.n6 A2.t1 225.954
R227 A2.n0 A2.t0 212.079
R228 A2.n10 A2.t7 212.079
R229 A2.n7 A2.t4 212.079
R230 A2.n1 A2.t2 139.779
R231 A2.n5 A2.t6 139.779
R232 A2.n11 A2.t3 139.779
R233 A2.n2 A2.t5 139.779
R234 A2.n9 A2.n6 93.066
R235 A2.n4 A2.n3 76
R236 A2.n13 A2.n12 76
R237 A2.n9 A2.n8 76
R238 A2.n4 A2.n1 66.659
R239 A2.n12 A2.n11 26.29
R240 A2.n12 A2.n10 25.56
R241 A2.n13 A2.n9 17.066
R242 A2.n3 A2.n2 13.145
R243 A2 A2.n4 12.298
R244 A2.n1 A2.n0 10.954
R245 A2.n6 A2.n5 10.224
R246 A2 A2.n13 4.768
R247 A2.n8 A2.n7 0.73
R248 VPWR.n3 VPWR.n2 168.598
R249 VPWR.n11 VPWR.n10 164.634
R250 VPWR.n1 VPWR.n0 164.634
R251 VPWR.n5 VPWR.n4 164.399
R252 VPWR.n10 VPWR.t5 31.52
R253 VPWR.n2 VPWR.t3 27.58
R254 VPWR.n2 VPWR.t0 27.58
R255 VPWR.n4 VPWR.t1 27.58
R256 VPWR.n4 VPWR.t2 27.58
R257 VPWR.n10 VPWR.t6 27.58
R258 VPWR.n0 VPWR.t7 27.58
R259 VPWR.n0 VPWR.t4 27.58
R260 VPWR.n15 VPWR.n1 4.892
R261 VPWR.n7 VPWR.n6 4.65
R262 VPWR.n9 VPWR.n8 4.65
R263 VPWR.n12 VPWR.n11 4.65
R264 VPWR.n14 VPWR.n13 4.65
R265 VPWR.n6 VPWR.n5 2.258
R266 VPWR VPWR.n15 1.56
R267 VPWR.n7 VPWR.n3 0.39
R268 VPWR.n15 VPWR.n14 0.134
R269 VPWR.n9 VPWR.n7 0.119
R270 VPWR.n12 VPWR.n9 0.119
R271 VPWR.n14 VPWR.n12 0.119
R272 C1.n13 C1.t7 215
R273 C1.n0 C1.t4 212.079
R274 C1.n5 C1.t1 212.079
R275 C1.n9 C1.t0 212.079
R276 C1.n12 C1.t3 139.779
R277 C1.n8 C1.t6 139.779
R278 C1.n2 C1.t2 139.779
R279 C1.n1 C1.t5 139.779
R280 C1.n4 C1.n1 94.526
R281 C1 C1.n13 87.545
R282 C1.n4 C1.n3 76
R283 C1.n7 C1.n6 76
R284 C1.n11 C1.n10 76
R285 C1.n6 C1.n5 23.369
R286 C1.n7 C1.n4 17.066
R287 C1.n11 C1.n7 17.066
R288 C1.n3 C1.n2 14.606
R289 C1.n1 C1.n0 11.684
R290 C1.n9 C1.n8 11.684
R291 C1.n10 C1.n9 10.224
R292 C1.n13 C1.n12 8.763
R293 C1 C1.n11 5.521
R294 a_1205_47.n3 a_1205_47.t5 242.59
R295 a_1205_47.t3 a_1205_47.n5 180.653
R296 a_1205_47.n3 a_1205_47.n2 92.5
R297 a_1205_47.n4 a_1205_47.n1 92.5
R298 a_1205_47.n5 a_1205_47.n0 92.5
R299 a_1205_47.n4 a_1205_47.n3 74.857
R300 a_1205_47.n5 a_1205_47.n4 65.754
R301 a_1205_47.n1 a_1205_47.t6 42.461
R302 a_1205_47.n1 a_1205_47.t0 26.769
R303 a_1205_47.n0 a_1205_47.t1 25.846
R304 a_1205_47.n0 a_1205_47.t2 25.846
R305 a_1205_47.n2 a_1205_47.t4 25.846
R306 a_1205_47.n2 a_1205_47.t7 25.846
R307 A1.n10 A1.t1 242.751
R308 A1.n0 A1.t4 212.079
R309 A1.n5 A1.t6 212.079
R310 A1.n9 A1.t7 212.079
R311 A1.n1 A1.t3 157.306
R312 A1.n10 A1.t2 139.779
R313 A1.n6 A1.t5 139.779
R314 A1.n2 A1.t0 139.779
R315 A1.n4 A1.n1 93.066
R316 A1.n4 A1.n3 76
R317 A1.n8 A1.n7 76
R318 A1.n12 A1.n11 76
R319 A1.n7 A1.n5 23.369
R320 A1.n11 A1.n10 21.909
R321 A1 A1.n12 19.576
R322 A1.n8 A1.n4 17.066
R323 A1.n12 A1.n8 17.066
R324 A1.n1 A1.n0 10.224
R325 A1.n11 A1.n9 10.224
R326 A1.n7 A1.n6 8.763
R327 A1.n3 A1.n2 4.381
C0 A1 Y 0.20fF
C1 B1 Y 0.32fF
C2 C1 Y 0.32fF
C3 VPWR VGND 0.21fF
C4 Y VGND 0.70fF
C5 VPB VPWR 0.19fF
C6 D1 Y 0.49fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__and2_0.ext - technology: sky130A

.subckt sky130_fd_sc_hd__and2_0 VPWR VGND X B A VNB VPB
X0 VPWR.t1 B.t0 a_40_47.t1 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1 X.t1 a_40_47.t3 VPWR.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X2 VGND.t1 B.t1 a_123_47.t1 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3 X.t0 a_40_47.t4 VGND.t0 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 a_123_47.t0 A.t0 a_40_47.t0 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 a_40_47.t2 A.t1 VPWR.t2 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
R0 B.n1 B.t1 207.422
R1 B.n0 B.t0 202.132
R2 B.n0 B 78.909
R3 B.n2 B.n1 76
R4 B.n1 B.n0 36.826
R5 B.n2 B 10.278
R6  B.n2 2.909
R7 a_40_47.n2 a_40_47.n0 389.692
R8 a_40_47.n1 a_40_47.t3 277.544
R9 a_40_47.t0 a_40_47.n2 158.025
R10 a_40_47.n1 a_40_47.t4 143.131
R11 a_40_47.n2 a_40_47.n1 81.661
R12 a_40_47.n0 a_40_47.t2 70.357
R13 a_40_47.n0 a_40_47.t1 65.666
R14 VPWR.n1 VPWR.t2 380.004
R15 VPWR.n1 VPWR.n0 120.234
R16 VPWR.n0 VPWR.t1 74.031
R17 VPWR.n0 VPWR.t0 27.821
R18 VPWR VPWR.n1 0.088
R19 VPB.t1 VPB.t0 455.763
R20 VPB.t2 VPB.t1 260.436
R21 VPB VPB.t2 233.8
R22 X.n0 X.t0 219.416
R23 X.n0 X.t1 210.064
R24 X X.n0 1.905
R25 a_123_47.t0 a_123_47.t1 60
R26 VGND VGND.n0 96.634
R27 VGND.n0 VGND.t0 72.857
R28 VGND.n0 VGND.t1 58.571
R29 VNB VNB.t0 6923.53
R30 VNB.t2 VNB.t1 3947.06
R31 VNB.t0 VNB.t2 2329.41
R32 A.n0 A.t0 280.606
R33 A.n0 A.t1 159.362
R34 A A.n0 35.89
C0 X VGND 0.15fF
C1 VPWR X 0.18fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__and2_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__and2_1 VPWR VGND X B A VNB VPB
X0 VPWR.t2 B.t0 a_59_75.t2 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1 X.t1 a_59_75.t3 VPWR.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 VGND.t1 B.t1 a_145_75.t1 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3 a_59_75.t0 A.t0 VPWR.t1 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 X.t0 a_59_75.t4 VGND.t0 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 a_145_75.t0 A.t1 a_59_75.t1 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
R0 B.n0 B.t0 261.886
R1 B.n0 B.t1 155.846
R2 B B.n0 80.864
R3 a_59_75.n2 a_59_75.n1 380.446
R4 a_59_75.n0 a_59_75.t3 236.179
R5 a_59_75.n1 a_59_75.t1 222.061
R6 a_59_75.n0 a_59_75.t4 163.879
R7 a_59_75.n1 a_59_75.n0 76
R8 a_59_75.n2 a_59_75.t2 63.321
R9 a_59_75.t0 a_59_75.n2 63.321
R10 VPWR.n1 VPWR.t1 388.011
R11 VPWR.n1 VPWR.n0 183.665
R12 VPWR.n0 VPWR.t2 116.32
R13 VPWR.n0 VPWR.t0 28.462
R14 VPWR VPWR.n1 0.155
R15 VPB.t2 VPB.t0 319.626
R16 VPB VPB.t1 298.909
R17 VPB.t1 VPB.t2 248.598
R18 X.n0 X.t1 193.162
R19 X X.t0 176.924
R20 X X.n2 11.264
R21 X X.n1 6.656
R22 X.n2 X 6.144
R23 X.n2 X 4.634
R24 X.n1 X.n0 4.077
R25 X.n1 X 3.617
R26 X.n0 X 1.747
R27 a_145_75.t0 a_145_75.t1 77.142
R28 VGND VGND.n0 118.161
R29 VGND.n0 VGND.t1 72.857
R30 VGND.n0 VGND.t0 22.324
R31 VNB VNB.t1 7186.67
R32 VNB.t2 VNB.t0 2650.79
R33 VNB.t1 VNB.t2 2253.66
R34 A.n0 A.t0 256.068
R35 A.n0 A.t1 150.028
R36 A.n1 A.n0 76
R37 A.n2  11.833
R38 A.n1 A 7.68
R39 A.n2 A.n1 4.608
R40 A A.n2 4.588
C0 X VGND 0.15fF
C1 X VPWR 0.16fF
C2 A B 0.12fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__and2_2.ext - technology: sky130A

.subckt sky130_fd_sc_hd__and2_2 VPWR VGND A X B VNB VPB
X0 X.t3 a_61_75.t3 VPWR.t2 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 VPWR.t1 a_61_75.t4 X.t2 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 VPWR.t3 B.t0 a_61_75.t2 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3 VGND.t0 B.t1 a_147_75.t1 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 X.t1 a_61_75.t5 VGND.t2 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 VGND.t1 a_61_75.t6 X.t0 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 a_61_75.t0 A.t0 VPWR.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7 a_147_75.t0 A.t1 a_61_75.t1 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
R0 a_61_75.n4 a_61_75.n3 380.446
R1 a_61_75.n3 a_61_75.t1 222.061
R2 a_61_75.n0 a_61_75.t4 212.079
R3 a_61_75.n1 a_61_75.t3 212.079
R4 a_61_75.n0 a_61_75.t6 139.779
R5 a_61_75.n1 a_61_75.t5 139.779
R6 a_61_75.n3 a_61_75.n2 76
R7 a_61_75.n2 a_61_75.n0 65.727
R8 a_61_75.n4 a_61_75.t2 63.321
R9 a_61_75.t0 a_61_75.n4 63.321
R10 a_61_75.n2 a_61_75.n1 13.145
R11 VPWR.n7 VPWR.t0 382.792
R12 VPWR.n1 VPWR.n0 179.13
R13 VPWR.n2 VPWR.t1 172.63
R14 VPWR.n0 VPWR.t3 116.32
R15 VPWR.n0 VPWR.t2 28.462
R16 VPWR.n8 VPWR.n7 8.791
R17 VPWR.n2 VPWR.n1 6.703
R18 VPWR.n4 VPWR.n3 4.65
R19 VPWR.n6 VPWR.n5 4.65
R20 VPWR.n4 VPWR.n2 0.204
R21 VPWR.n6 VPWR.n4 0.119
R22 VPWR.n8 VPWR.n6 0.119
R23 VPWR VPWR.n8 0.022
R24 X.n1 X.n0 146.88
R25 X X.n3 99.341
R26 X.n3 X.t0 47.076
R27 X.n0 X.t3 46.295
R28 X.n0 X.t2 30.535
R29 X.n3 X.t1 24.923
R30 X X.n4 11.264
R31 X X.n2 6.656
R32 X.n4 X 6.144
R33 X.n4 X 4.634
R34 X.n2 X.n1 4.166
R35 X.n2 X 3.697
R36 X.n1 X 1.786
R37 VPB.t2 VPB.t1 319.626
R38 VPB.t3 VPB.t2 319.626
R39 VPB VPB.t0 304.828
R40 VPB.t0 VPB.t3 248.598
R41 B.n0 B.t0 261.886
R42 B.n0 B.t1 155.846
R43 B B.n0 81.376
R44 a_147_75.t0 a_147_75.t1 77.142
R45 VGND.n1 VGND.n0 117.886
R46 VGND.n1 VGND.t1 114.098
R47 VGND.n0 VGND.t0 72.857
R48 VGND.n0 VGND.t2 22.324
R49 VGND VGND.n1 0.349
R50 VNB VNB.t0 7255.4
R51 VNB.t1 VNB.t3 2650.79
R52 VNB.t3 VNB.t2 2610.99
R53 VNB.t0 VNB.t1 2253.66
R54 A.n0 A.t0 256.068
R55 A.n0 A.t1 150.028
R56 A.n1 A.n0 76
R57 A.n2  9.955
R58 A.n1 A 7.168
R59 A A.n2 3.86
R60 A.n2 A.n1 3.328
C0 X VPWR 0.32fF
C1 B A 0.11fF
C2 X VGND 0.24fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__and2_4.ext - technology: sky130A

.subckt sky130_fd_sc_hd__and2_4 X B A VGND VPWR VNB VPB
X0 VPWR.t0 B.t0 a_27_47.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_27_47.t2 A.t0 VPWR.t5 VPB.t5 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 X.t3 a_27_47.t3 VGND.t4 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 VPWR.t3 a_27_47.t4 X.t7 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 VGND.t0 B.t1 a_110_47.t0 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 X.t6 a_27_47.t5 VPWR.t2 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 a_110_47.t1 A.t1 a_27_47.t1 VNB.t5 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 VPWR.t1 a_27_47.t6 X.t5 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 VGND.t3 a_27_47.t7 X.t2 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 VGND.t2 a_27_47.t8 X.t1 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 X.t4 a_27_47.t9 VPWR.t4 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 X.t0 a_27_47.t10 VGND.t1 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
R0 B.n0 B.t0 241.534
R1 B.n0 B.t1 169.234
R2 B B.n0 87.248
R3 a_27_47.n11 a_27_47.n10 219.41
R4 a_27_47.n5 a_27_47.t4 212.079
R5 a_27_47.n0 a_27_47.t6 212.079
R6 a_27_47.n2 a_27_47.t5 212.079
R7 a_27_47.n7 a_27_47.t9 212.079
R8 a_27_47.n10 a_27_47.t1 155.448
R9 a_27_47.n5 a_27_47.t8 139.779
R10 a_27_47.n0 a_27_47.t7 139.779
R11 a_27_47.n2 a_27_47.t10 139.779
R12 a_27_47.n7 a_27_47.t3 139.779
R13 a_27_47.n4 a_27_47.n1 88.991
R14 a_27_47.n9 a_27_47.n8 76
R15 a_27_47.n4 a_27_47.n3 76
R16 a_27_47.n6 a_27_47.n5 76
R17 a_27_47.t0 a_27_47.n11 27.58
R18 a_27_47.n11 a_27_47.t2 27.58
R19 a_27_47.n1 a_27_47.n0 26.29
R20 a_27_47.n3 a_27_47.n2 13.145
R21 a_27_47.n8 a_27_47.n7 13.145
R22 a_27_47.n6 a_27_47.n4 12.991
R23 a_27_47.n9 a_27_47.n6 12.991
R24 a_27_47.n10 a_27_47.n9 9.361
R25 VPWR.n2 VPWR.t1 194.862
R26 VPWR.n10 VPWR.t5 191.794
R27 VPWR.n6 VPWR.n5 163.438
R28 VPWR.n1 VPWR.n0 163.438
R29 VPWR.n5 VPWR.t4 35.46
R30 VPWR.n5 VPWR.t0 34.475
R31 VPWR.n0 VPWR.t2 27.58
R32 VPWR.n0 VPWR.t3 27.58
R33 VPWR.n4 VPWR.n3 4.65
R34 VPWR.n7 VPWR.n6 4.65
R35 VPWR.n9 VPWR.n8 4.65
R36 VPWR.n11 VPWR.n10 4.65
R37 VPWR.n2 VPWR.n1 3.832
R38 VPWR.n4 VPWR.n2 0.261
R39 VPWR.n7 VPWR.n4 0.119
R40 VPWR.n9 VPWR.n7 0.119
R41 VPWR.n11 VPWR.n9 0.119
R42 VPWR VPWR.n11 0.022
R43 VPB.t0 VPB.t1 298.909
R44 VPB.t3 VPB.t2 254.517
R45 VPB.t4 VPB.t3 254.517
R46 VPB.t1 VPB.t4 254.517
R47 VPB.t5 VPB.t0 254.517
R48 VPB VPB.t5 195.327
R49 A.n0 A.t0 235.819
R50 A.n0 A.t1 163.519
R51 A A.n0 87.767
R52 VGND.n4 VGND.t3 194.517
R53 VGND.n3 VGND.n2 106.463
R54 VGND.n1 VGND.n0 106.463
R55 VGND.n0 VGND.t4 39.692
R56 VGND.n0 VGND.t0 38.769
R57 VGND.n2 VGND.t1 25.846
R58 VGND.n2 VGND.t2 25.846
R59 VGND.n6 VGND.n5 4.65
R60 VGND.n7 VGND.n1 3.881
R61 VGND.n4 VGND.n3 3.832
R62 VGND.n6 VGND.n4 0.261
R63 VGND VGND.n7 0.239
R64 VGND.n7 VGND.n6 0.141
R65 X.n2 X.n1 214.04
R66 X.n5 X.n4 140.36
R67 X.n2 X.n0 105.451
R68 X X.n2 61.048
R69 X.n5 X.n3 49.316
R70 X.n0 X.t5 27.58
R71 X.n0 X.t6 27.58
R72 X.n1 X.t7 27.58
R73 X.n1 X.t4 27.58
R74 X.n4 X.t1 25.846
R75 X.n4 X.t3 25.846
R76 X.n3 X.t2 25.846
R77 X.n3 X.t0 25.846
R78 X X.n5 22.191
R79 VNB VNB.t5 6102.26
R80 VNB.t0 VNB.t4 2780.22
R81 VNB.t1 VNB.t3 2079.12
R82 VNB.t2 VNB.t1 2079.12
R83 VNB.t4 VNB.t2 2079.12
R84 VNB.t5 VNB.t0 1740.66
R85 a_110_47.t0 a_110_47.t1 38.769
C0 VGND X 0.26fF
C1 B A 0.12fF
C2 VPWR X 0.49fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__and2b_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__and2b_1 X A_N B VGND VPWR VNB VPB
X0 VPWR.t0 B.t0 a_207_413.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1 X.t1 a_207_413.t3 VPWR.t1 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 a_297_47.t1 a_27_413.t2 a_207_413.t1 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3 X.t0 a_207_413.t4 VGND.t1 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 a_207_413.t2 a_27_413.t3 VPWR.t3 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 VPWR.t2 A_N.t0 a_27_413.t0 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 VGND.t0 B.t1 a_297_47.t0 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7 a_27_413.t1 A_N.t1 VGND.t2 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
R0 B.n0 B.t1 293.968
R1 B.n0 B.t0 138.336
R2 B.n1 B.n0 76
R3 B B.n1 14.038
R4 B.n1 B 4.954
R5 a_207_413.n2 a_207_413.n1 333.182
R6 a_207_413.n0 a_207_413.t3 240.482
R7 a_207_413.n1 a_207_413.t1 169.75
R8 a_207_413.n0 a_207_413.t4 166.691
R9 a_207_413.n1 a_207_413.n0 98.923
R10 a_207_413.t0 a_207_413.n2 68.011
R11 a_207_413.n2 a_207_413.t2 68.011
R12 VPWR.n9 VPWR.n8 309.954
R13 VPWR.n3 VPWR.n2 292.5
R14 VPWR.n1 VPWR.n0 292.5
R15 VPWR.n8 VPWR.t3 96.154
R16 VPWR.n2 VPWR.t0 86.773
R17 VPWR.n0 VPWR.t1 66.839
R18 VPWR.n8 VPWR.t2 63.321
R19 VPWR.n5 VPWR.n1 5.608
R20 VPWR.n5 VPWR.n4 4.65
R21 VPWR.n7 VPWR.n6 4.65
R22 VPWR.n10 VPWR.n9 3.932
R23 VPWR.n4 VPWR.n3 1
R24 VPWR.n10 VPWR.n7 0.137
R25 VPWR VPWR.n10 0.123
R26 VPWR.n7 VPWR.n5 0.119
R27 VPB.t0 VPB.t1 526.791
R28 VPB.t2 VPB.t3 290.031
R29 VPB.t3 VPB.t0 260.436
R30 VPB VPB.t2 192.367
R31 X.n1 X.t1 212.393
R32 X.n0 X.t0 117.423
R33 X X.n0 79.483
R34 X.n1 X 7.735
R35 X.n0 X 6.666
R36 X X.n1 6.365
R37 a_27_413.t0 a_27_413.n1 433.056
R38 a_27_413.n0 a_27_413.t3 381.656
R39 a_27_413.n0 a_27_413.t2 197.62
R40 a_27_413.n1 a_27_413.t1 151.191
R41 a_27_413.n1 a_27_413.n0 88.993
R42 a_297_47.t0 a_297_47.t1 68.571
R43 VNB VNB.t3 6470.59
R44 VNB.t3 VNB.t2 6082.35
R45 VNB.t2 VNB.t0 2523.53
R46 VNB.t0 VNB.t1 2317.53
R47 VGND.n1 VGND.t2 151.952
R48 VGND.n1 VGND.n0 111.502
R49 VGND.n0 VGND.t0 58.571
R50 VGND.n0 VGND.t1 25.428
R51 VGND VGND.n1 0.045
R52 A_N.n0 A_N.t0 327.988
R53 A_N.n0 A_N.t1 199.455
R54 A_N.n1 A_N.n0 76
R55 A_N.n1 A_N 12.16
R56 A_N A_N.n1 2.346
C0 B VPWR 0.15fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__and2b_2.ext - technology: sky130A

.subckt sky130_fd_sc_hd__and2b_2 VPWR VGND X B A_N VNB VPB
X0 VPWR.t2 a_212_413.t3 X.t2 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_297_47.t1 a_27_413.t2 a_212_413.t1 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 X.t3 a_212_413.t4 VPWR.t1 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 X.t1 a_212_413.t5 VGND.t2 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 a_212_413.t2 a_27_413.t3 VPWR.t4 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 VPWR.t3 A_N.t0 a_27_413.t0 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 VPWR.t0 B.t0 a_212_413.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7 VGND.t0 B.t1 a_297_47.t0 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 VGND.t1 a_212_413.t6 X.t0 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 a_27_413.t1 A_N.t1 VGND.t3 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
R0 a_212_413.n3 a_212_413.n2 333.182
R1 a_212_413.n0 a_212_413.t3 212.079
R2 a_212_413.n1 a_212_413.t4 212.079
R3 a_212_413.n2 a_212_413.t1 171.391
R4 a_212_413.n0 a_212_413.t6 136.566
R5 a_212_413.n1 a_212_413.t5 136.566
R6 a_212_413.n2 a_212_413.n1 109.015
R7 a_212_413.t0 a_212_413.n3 68.011
R8 a_212_413.n3 a_212_413.t2 68.011
R9 a_212_413.n1 a_212_413.n0 59.541
R10 X.n0 X 295.647
R11 X.n3 X.n0 292.5
R12 X.n2 X.n1 92.5
R13 X.n3 X.n2 81.836
R14 X.n0 X.t2 26.595
R15 X.n0 X.t3 26.595
R16 X.n1 X.t0 24.923
R17 X.n1 X.t1 24.923
R18 X.n2 X 2.178
R19 X X.n3 1.468
R20 VPWR.n10 VPWR.n9 309.954
R21 VPWR.n4 VPWR.n3 292.5
R22 VPWR.n1 VPWR.n0 292.5
R23 VPWR.n2 VPWR.t2 205.541
R24 VPWR.n9 VPWR.t4 107.88
R25 VPWR.n3 VPWR.t0 86.773
R26 VPWR.n0 VPWR.t1 69.184
R27 VPWR.n9 VPWR.t3 63.321
R28 VPWR.n2 VPWR.n1 4.862
R29 VPWR.n6 VPWR.n5 4.65
R30 VPWR.n8 VPWR.n7 4.65
R31 VPWR.n11 VPWR.n10 3.932
R32 VPWR.n5 VPWR.n4 1.5
R33 VPWR.n6 VPWR.n2 0.217
R34 VPWR.n11 VPWR.n8 0.137
R35 VPWR VPWR.n11 0.121
R36 VPWR.n8 VPWR.n6 0.119
R37 VPB.t0 VPB.t1 529.75
R38 VPB.t3 VPB.t4 304.828
R39 VPB.t4 VPB.t0 260.436
R40 VPB.t1 VPB.t2 248.598
R41 VPB VPB.t3 189.408
R42 a_27_413.t0 a_27_413.n1 433.334
R43 a_27_413.n0 a_27_413.t3 381.656
R44 a_27_413.n0 a_27_413.t2 189.586
R45 a_27_413.n1 a_27_413.t1 151.588
R46 a_27_413.n1 a_27_413.n0 89.769
R47 a_297_47.t0 a_297_47.t1 77.142
R48 VNB VNB.t3 6438.23
R49 VNB.t3 VNB.t4 6082.35
R50 VNB.t4 VNB.t0 2717.65
R51 VNB.t0 VNB.t2 2327.87
R52 VNB.t2 VNB.t1 2030.77
R53 VGND.n9 VGND.t3 148.331
R54 VGND.n2 VGND.t1 147.584
R55 VGND.n1 VGND.n0 107.54
R56 VGND.n0 VGND.t0 58.571
R57 VGND.n0 VGND.t2 24.923
R58 VGND.n10 VGND.n9 4.65
R59 VGND.n4 VGND.n3 4.65
R60 VGND.n6 VGND.n5 4.65
R61 VGND.n8 VGND.n7 4.65
R62 VGND.n2 VGND.n1 3.752
R63 VGND.n4 VGND.n2 0.246
R64 VGND.n6 VGND.n4 0.119
R65 VGND.n8 VGND.n6 0.119
R66 VGND.n10 VGND.n8 0.119
R67 VGND VGND.n10 0.02
R68 A_N.n0 A_N.t0 328.318
R69 A_N.n0 A_N.t1 199.785
R70 A_N.n1 A_N.n0 76
R71 A_N.n1 A_N 13.226
R72 A_N A_N.n1 1.28
R73 B.n0 B.t1 293.653
R74 B.n0 B.t0 138.336
R75 B.n1 B.n0 76
R76 B.n1 B 17.548
R77 B B.n1 4.954
C0 VGND X 0.16fF
C1 VPWR X 0.17fF
C2 B VPWR 0.15fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__and2b_4.ext - technology: sky130A

.subckt sky130_fd_sc_hd__and2b_4 B X A_N VGND VPWR VNB VPB
X0 X.t3 a_27_47.t3 VGND.t3 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 VGND.t4 B.t0 a_109_47.t1 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 VPWR.t6 B.t1 a_27_47.t0 VPB.t6 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 a_33_199.t0 A_N.t0 VGND.t5 VNB.t6 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 a_33_199.t1 A_N.t1 VPWR.t4 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 VPWR.t3 a_27_47.t4 X.t7 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 VGND.t2 a_27_47.t5 X.t2 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 X.t6 a_27_47.t6 VPWR.t2 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 VGND.t1 a_27_47.t7 X.t1 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 VPWR.t1 a_27_47.t8 X.t5 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 X.t4 a_27_47.t9 VPWR.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 a_27_47.t1 a_33_199.t2 VPWR.t5 VPB.t5 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 X.t0 a_27_47.t10 VGND.t0 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 a_109_47.t0 a_33_199.t3 a_27_47.t2 VNB.t5 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
R0 a_27_47.n12 a_27_47.n11 330.734
R1 a_27_47.n0 a_27_47.t4 212.079
R2 a_27_47.n1 a_27_47.t6 212.079
R3 a_27_47.n4 a_27_47.t8 212.079
R4 a_27_47.n8 a_27_47.t9 212.079
R5 a_27_47.n11 a_27_47.t2 154.281
R6 a_27_47.n0 a_27_47.t5 139.779
R7 a_27_47.n8 a_27_47.t3 139.779
R8 a_27_47.n5 a_27_47.t7 139.779
R9 a_27_47.n2 a_27_47.t10 139.779
R10 a_27_47.n7 a_27_47.n3 88.088
R11 a_27_47.n10 a_27_47.n9 76
R12 a_27_47.n7 a_27_47.n6 76
R13 a_27_47.n1 a_27_47.n0 61.345
R14 a_27_47.t0 a_27_47.n12 26.595
R15 a_27_47.n12 a_27_47.t1 26.595
R16 a_27_47.n3 a_27_47.n2 13.875
R17 a_27_47.n9 a_27_47.n8 12.415
R18 a_27_47.n10 a_27_47.n7 12.088
R19 a_27_47.n11 a_27_47.n10 8.711
R20 a_27_47.n5 a_27_47.n4 2.921
R21 a_27_47.n2 a_27_47.n1 1.46
R22 a_27_47.n6 a_27_47.n5 0.73
R23 VGND.n5 VGND.n2 154.922
R24 VGND.n4 VGND.n3 106.463
R25 VGND.n1 VGND.n0 106.463
R26 VGND.n2 VGND.t5 61.428
R27 VGND.n0 VGND.t3 39.692
R28 VGND.n0 VGND.t4 37.846
R29 VGND.n3 VGND.t0 26.769
R30 VGND.n3 VGND.t1 24.923
R31 VGND.n2 VGND.t2 20.177
R32 VGND.n7 VGND.n6 4.65
R33 VGND.n8 VGND.n1 3.881
R34 VGND.n5 VGND.n4 3.851
R35 VGND.n7 VGND.n5 0.249
R36 VGND VGND.n8 0.239
R37 VGND.n8 VGND.n7 0.141
R38 X.n2 X.n0 341.534
R39 X.n2 X.n1 292.5
R40 X.n5 X.n4 143.362
R41 X.n5 X.n3 92.5
R42 X X.n2 37.737
R43 X.n0 X.t4 32.505
R44 X.n4 X.t1 26.769
R45 X.n1 X.t7 26.595
R46 X.n1 X.t6 26.595
R47 X.n0 X.t5 26.595
R48 X.n3 X.t2 25.846
R49 X.n3 X.t0 25.846
R50 X.n4 X.t3 24.923
R51 X X.n5 1.103
R52 VNB VNB.t5 6078.09
R53 VNB.t4 VNB.t3 2756.04
R54 VNB.t2 VNB.t6 2400.4
R55 VNB.t0 VNB.t2 2079.12
R56 VNB.t1 VNB.t0 2079.12
R57 VNB.t3 VNB.t1 2079.12
R58 VNB.t5 VNB.t4 1789.01
R59 B.n0 B.t1 241.534
R60 B.n0 B.t0 169.234
R61 B B.n0 86.86
R62 a_109_47.t0 a_109_47.t1 40.615
R63 VPWR.n10 VPWR.t5 575.999
R64 VPWR.n2 VPWR.t3 573.754
R65 VPWR.n6 VPWR.n5 306.463
R66 VPWR.n1 VPWR.n0 306.463
R67 VPWR.t3 VPWR.t4 131.152
R68 VPWR.n5 VPWR.t6 37.43
R69 VPWR.n5 VPWR.t0 35.46
R70 VPWR.n0 VPWR.t2 26.595
R71 VPWR.n0 VPWR.t1 26.595
R72 VPWR.n4 VPWR.n3 4.65
R73 VPWR.n7 VPWR.n6 4.65
R74 VPWR.n9 VPWR.n8 4.65
R75 VPWR.n11 VPWR.n10 4.65
R76 VPWR.n2 VPWR.n1 3.812
R77 VPWR.n4 VPWR.n2 0.255
R78 VPWR.n7 VPWR.n4 0.119
R79 VPWR.n9 VPWR.n7 0.119
R80 VPWR.n11 VPWR.n9 0.119
R81 VPWR VPWR.n11 0.022
R82 VPB.t6 VPB.t0 307.788
R83 VPB.t3 VPB.t4 298.909
R84 VPB.t0 VPB.t1 266.355
R85 VPB.t2 VPB.t3 248.598
R86 VPB.t1 VPB.t2 248.598
R87 VPB.t5 VPB.t6 248.598
R88 VPB VPB.t5 192.367
R89 A_N.n0 A_N.t1 143.483
R90 A_N.n0 A_N.t0 129.785
R91 A_N A_N.n0 78.308
R92 a_33_199.n1 a_33_199.n0 383.72
R93 a_33_199.n1 a_33_199.t1 358.166
R94 a_33_199.n0 a_33_199.t2 233.007
R95 a_33_199.t0 a_33_199.n1 202.527
R96 a_33_199.n0 a_33_199.t3 160.707
C0 X VGND 0.12fF
C1 X A_N 0.14fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__and3_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__and3_1 VGND VPWR X B A C VNB VPB
X0 VPWR.t2 A.t0 a_27_47.t2 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1 VPWR.t3 C.t0 a_27_47.t3 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 a_181_47.t0 B.t0 a_109_47.t1 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3 VGND.t1 C.t1 a_181_47.t1 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 a_27_47.t0 B.t1 VPWR.t1 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 X.t1 a_27_47.t4 VPWR.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 X.t0 a_27_47.t5 VGND.t0 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 a_109_47.t0 A.t1 a_27_47.t1 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
R0 A.n0 A.t0 183.503
R1 A.n0 A.t1 114.532
R2 A A.n0 79.84
R3 a_27_47.n1 a_27_47.t2 406.82
R4 a_27_47.n2 a_27_47.n1 374.391
R5 a_27_47.n3 a_27_47.n2 292.5
R6 a_27_47.n1 a_27_47.t1 242.882
R7 a_27_47.n0 a_27_47.t4 241.534
R8 a_27_47.n0 a_27_47.t5 169.234
R9 a_27_47.n2 a_27_47.n0 106.72
R10 a_27_47.t0 a_27_47.n3 84.428
R11 a_27_47.n3 a_27_47.t3 63.321
R12 VPWR.n2 VPWR.n0 428.987
R13 VPWR.n2 VPWR.n1 320.806
R14 VPWR.n0 VPWR.t3 93.809
R15 VPWR.n1 VPWR.t1 63.321
R16 VPWR.n1 VPWR.t2 63.321
R17 VPWR.n0 VPWR.t0 26.972
R18 VPWR VPWR.n2 0.121
R19 VPB.t3 VPB.t0 281.152
R20 VPB.t1 VPB.t3 275.233
R21 VPB.t2 VPB.t1 248.598
R22 VPB VPB.t2 192.367
R23 C.n0 C.t1 173.339
R24 C.n0 C.t0 162.808
R25 C.n1 C.n0 89.187
R26 C.n1 C 2.111
R27 C C.n1 0.969
R28 B.t1 B.t0 395.01
R29 B B.t1 244.948
R30 a_109_47.t0 a_109_47.t1 60
R31 a_181_47.t0 a_181_47.t1 60
R32 VNB VNB.t1 6470.59
R33 VNB.t3 VNB.t0 3397.06
R34 VNB.t2 VNB.t3 2329.41
R35 VNB.t1 VNB.t2 2329.41
R36 VGND VGND.n0 119.936
R37 VGND.n0 VGND.t1 101.428
R38 VGND.n0 VGND.t0 25.934
R39 X.n0 X.t1 172.279
R40 X.n1 X.t0 117.423
R41 X.n1 X.n0 100.727
R42 X.n0 X 4.521
R43 X X.n1 4.184
C0 X VPWR 0.11fF
C1 X VGND 0.10fF
C2 B VPWR 0.19fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__and3_2.ext - technology: sky130A

.subckt sky130_fd_sc_hd__and3_2 B X A C VPWR VGND VNB VPB
X0 VPWR.t3 a_29_311.t4 X.t1 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 X.t0 a_29_311.t5 VPWR.t2 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 VPWR.t1 A.t0 a_29_311.t1 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3 VGND.t1 a_29_311.t6 X.t3 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 a_184_53.t0 B.t0 a_112_53.t0 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 VPWR.t4 C.t0 a_29_311.t3 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 X.t2 a_29_311.t7 VGND.t0 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 a_112_53.t1 A.t1 a_29_311.t2 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 a_29_311.t0 B.t1 VPWR.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9 VGND.t2 C.t1 a_184_53.t1 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
R0 a_29_311.n3 a_29_311.t1 389.828
R1 a_29_311.n5 a_29_311.n4 292.5
R2 a_29_311.n0 a_29_311.t4 214.269
R3 a_29_311.n1 a_29_311.t5 212.079
R4 a_29_311.n3 a_29_311.t2 201.922
R5 a_29_311.n2 a_29_311.t7 139.779
R6 a_29_311.n0 a_29_311.t6 139.779
R7 a_29_311.n4 a_29_311.n2 132.169
R8 a_29_311.n1 a_29_311.n0 59.154
R9 a_29_311.n5 a_29_311.t3 48.587
R10 a_29_311.n6 a_29_311.t0 42.959
R11 a_29_311.n6 a_29_311.n5 36.585
R12 a_29_311.n7 a_29_311.n6 27.58
R13 a_29_311.n4 a_29_311.n3 16.268
R14 a_29_311.n2 a_29_311.n1 2.19
R15 X.n1 X.n0 146.364
R16 X.n3 X.n2 92.5
R17 X X.n1 44.847
R18 X X.n3 29.029
R19 X.n0 X.t1 26.595
R20 X.n0 X.t0 26.595
R21 X.n2 X.t3 24.923
R22 X.n2 X.t2 24.923
R23 X.n3 X 5.376
R24 X.n1 X 3.843
R25 VPWR.n8 VPWR.n1 308.361
R26 VPWR.n4 VPWR.t3 201.71
R27 VPWR.n3 VPWR.n2 176.216
R28 VPWR.n2 VPWR.t4 98.5
R29 VPWR.n1 VPWR.t0 63.321
R30 VPWR.n1 VPWR.t1 63.321
R31 VPWR.n7 VPWR.n6 33.226
R32 VPWR.n6 VPWR.n3 30.494
R33 VPWR.n2 VPWR.t2 26.595
R34 VPWR VPWR.n8 12.045
R35 VPWR.n6 VPWR.n5 4.65
R36 VPWR.n7 VPWR.n0 4.65
R37 VPWR.n4 VPWR.n3 3.851
R38 VPWR.n8 VPWR.n7 1.327
R39 VPWR.n5 VPWR.n4 0.23
R40 VPWR.n5 VPWR.n0 0.119
R41 VPWR VPWR.n0 0.119
R42 VPB.t4 VPB.t2 292.99
R43 VPB.t0 VPB.t4 281.152
R44 VPB.t2 VPB.t3 248.598
R45 VPB.t1 VPB.t0 248.598
R46 VPB VPB.t1 198.286
R47 A.n0 A.t1 186.028
R48 A.n0 A.t0 160.321
R49 A A.n0 89.132
R50 VGND.n1 VGND.t1 145.505
R51 VGND.n1 VGND.n0 116.283
R52 VGND.n0 VGND.t2 88.593
R53 VGND.n0 VGND.t0 21.907
R54 VGND VGND.n1 0.452
R55 VNB.t4 VNB.t2 32341.4
R56 VNB VNB.t1 7344.12
R57 VNB.t0 VNB.t4 2620.59
R58 VNB.t1 VNB.t0 2329.41
R59 VNB.t2 VNB.t3 2030.77
R60 B.t1 B.t0 398.279
R61 B B.t1 227.032
R62 a_112_53.t0 a_112_53.t1 60
R63 a_184_53.t0 a_184_53.t1 72.857
R64 C.n0 C.t1 194.998
R65 C.n0 C.t0 146.798
R66 C C.n0 88.331
R67  C 18.554
C0 VPWR B 0.18fF
C1 X VPWR 0.32fF
C2 X VGND 0.20fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__and3_4.ext - technology: sky130A

.subckt sky130_fd_sc_hd__and3_4 A B C X VGND VPWR VNB VPB
X0 VPWR.t1 A.t0 a_94_47.t1 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_294_47.t1 B.t0 a_185_47.t1 VNB sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 a_185_47.t0 A.t1 a_94_47.t2 VNB sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 VPWR.t5 a_94_47.t4 X.t3 VPB.t5 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 VGND.t4 C.t0 a_294_47.t0 VNB sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 a_94_47.t3 B.t1 VPWR.t6 VPB.t6 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 X.t2 a_94_47.t5 VPWR.t4 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 X.t7 a_94_47.t6 VGND.t3 VNB sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 VPWR.t0 C.t1 a_94_47.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 X.t6 a_94_47.t7 VGND.t2 VNB sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 VGND.t1 a_94_47.t8 X.t5 VNB sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 VPWR.t3 a_94_47.t9 X.t1 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 VGND.t0 a_94_47.t10 X.t4 VNB sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 X.t0 a_94_47.t11 VPWR.t2 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
R0 A.n0 A.t0 241.534
R1 A.n0 A.t1 169.234
R2 A A.n0 82.863
R3 A.n1 A 13.542
R4 A.n1  5.376
R5  A.n1 3.524
R6 a_94_47.n11 a_94_47.t1 260.47
R7 a_94_47.n5 a_94_47.t9 212.079
R8 a_94_47.n0 a_94_47.t4 212.079
R9 a_94_47.n2 a_94_47.t11 212.079
R10 a_94_47.n7 a_94_47.t5 212.079
R11 a_94_47.n10 a_94_47.t2 190.758
R12 a_94_47.n12 a_94_47.n11 173.033
R13 a_94_47.n5 a_94_47.t10 139.779
R14 a_94_47.n0 a_94_47.t8 139.779
R15 a_94_47.n2 a_94_47.t6 139.779
R16 a_94_47.n7 a_94_47.t7 139.779
R17 a_94_47.n4 a_94_47.n1 88.991
R18 a_94_47.n9 a_94_47.n8 76
R19 a_94_47.n4 a_94_47.n3 76
R20 a_94_47.n6 a_94_47.n5 76
R21 a_94_47.n11 a_94_47.n10 46.753
R22 a_94_47.t0 a_94_47.n12 27.58
R23 a_94_47.n12 a_94_47.t3 27.58
R24 a_94_47.n1 a_94_47.n0 26.29
R25 a_94_47.n3 a_94_47.n2 13.145
R26 a_94_47.n8 a_94_47.n7 13.145
R27 a_94_47.n6 a_94_47.n4 12.991
R28 a_94_47.n9 a_94_47.n6 12.991
R29 a_94_47.n10 a_94_47.n9 9.361
R30 VPWR.n2 VPWR.t5 194.862
R31 VPWR.n1 VPWR.n0 163.438
R32 VPWR.n6 VPWR.n5 163.438
R33 VPWR.n11 VPWR.n10 158.869
R34 VPWR.n10 VPWR.t1 40.385
R35 VPWR.n10 VPWR.t6 37.43
R36 VPWR.n5 VPWR.t4 35.46
R37 VPWR.n5 VPWR.t0 34.475
R38 VPWR.n0 VPWR.t2 27.58
R39 VPWR.n0 VPWR.t3 27.58
R40 VPWR.n4 VPWR.n3 4.65
R41 VPWR.n7 VPWR.n6 4.65
R42 VPWR.n9 VPWR.n8 4.65
R43 VPWR.n2 VPWR.n1 3.832
R44 VPWR.n12 VPWR.n11 3.738
R45 VPWR.n4 VPWR.n2 0.261
R46 VPWR VPWR.n12 0.235
R47 VPWR.n12 VPWR.n9 0.145
R48 VPWR.n7 VPWR.n4 0.119
R49 VPWR.n9 VPWR.n7 0.119
R50 VPB VPB.t1 417.289
R51 VPB.t1 VPB.t6 322.585
R52 VPB.t0 VPB.t4 298.909
R53 VPB.t2 VPB.t5 254.517
R54 VPB.t3 VPB.t2 254.517
R55 VPB.t4 VPB.t3 254.517
R56 VPB.t6 VPB.t0 254.517
R57 B.n0 B.t1 235.819
R58 B.n0 B.t0 163.519
R59 B B.n0 78.427
R60  B 15.006
R61 a_185_47.t0 a_185_47.t1 72.923
R62 a_294_47.t0 a_294_47.t1 38.769
R63 X.n2 X.n1 214.04
R64 X.n5 X.n4 140.36
R65 X.n2 X.n0 105.451
R66 X X.n2 61.048
R67 X.n5 X.n3 49.316
R68 X.n0 X.t3 27.58
R69 X.n0 X.t0 27.58
R70 X.n1 X.t1 27.58
R71 X.n1 X.t2 27.58
R72 X.n4 X.t4 25.846
R73 X.n4 X.t6 25.846
R74 X.n3 X.t5 25.846
R75 X.n3 X.t7 25.846
R76 X X.n5 22.191
R77 C.n0 C.t1 241.534
R78 C.n0 C.t0 169.234
R79 C C.n0 87.248
R80 VGND.n4 VGND.t1 194.517
R81 VGND.n3 VGND.n2 106.463
R82 VGND.n1 VGND.n0 106.463
R83 VGND.n0 VGND.t4 44.307
R84 VGND.n0 VGND.t2 34.153
R85 VGND.n2 VGND.t3 25.846
R86 VGND.n2 VGND.t0 25.846
R87 VGND.n6 VGND.n5 4.65
R88 VGND.n7 VGND.n1 3.936
R89 VGND.n4 VGND.n3 3.832
R90 VGND VGND.n7 0.48
R91 VGND.n6 VGND.n4 0.261
R92 VGND.n7 VGND.n6 0.139
C0 X VGND 0.26fF
C1 A B 0.10fF
C2 B C 0.12fF
C3 VPWR X 0.49fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__and3b_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__and3b_1 A_N B X C VGND VPWR VNB VPB
X0 a_109_93.t0 A_N.t0 VGND.t2 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1 X.t1 a_209_311.t4 VPWR.t3 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 a_109_93.t1 A_N.t1 VPWR.t1 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3 a_296_53.t0 a_109_93.t2 a_209_311.t1 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 VPWR.t0 C.t0 a_209_311.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 a_368_53.t0 B.t0 a_296_53.t1 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 X.t0 a_209_311.t5 VGND.t0 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 a_209_311.t3 B.t1 VPWR.t4 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 VPWR.t2 a_109_93.t3 a_209_311.t2 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9 VGND.t1 C.t1 a_368_53.t1 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
R0 A_N.n0 A_N.t1 204.655
R1 A_N.n2 A_N.t0 121.108
R2 A_N.n3 A_N.n2 76
R3 A_N.n1 A_N.n0 76
R4 A_N A_N.n3 10.729
R5 A_N.n1 A_N 9.6
R6 A_N A_N.n1 3.2
R7 A_N.n3 A_N 2.07
R8 VGND.n1 VGND.t2 171.022
R9 VGND.n1 VGND.n0 114.709
R10 VGND.n0 VGND.t1 83.898
R11 VGND.n0 VGND.t0 21.794
R12 VGND VGND.n1 0.038
R13 a_109_93.n1 a_109_93.t1 419.855
R14 a_109_93.n0 a_109_93.t2 186.028
R15 a_109_93.n0 a_109_93.t3 160.321
R16 a_109_93.n2 a_109_93.n1 103.508
R17 a_109_93.n1 a_109_93.n0 100.32
R18 a_109_93.n2 a_109_93.t0 30
R19 VNB.t1 VNB.t0 32220.6
R20 VNB VNB.t2 6869.12
R21 VNB.t2 VNB.t3 5366.18
R22 VNB.t4 VNB.t1 2620.59
R23 VNB.t3 VNB.t4 2329.41
R24 a_209_311.n1 a_209_311.t2 376.851
R25 a_209_311.n3 a_209_311.n2 292.5
R26 a_209_311.n0 a_209_311.t4 241.534
R27 a_209_311.n1 a_209_311.t1 210.234
R28 a_209_311.n0 a_209_311.t5 169.234
R29 a_209_311.n2 a_209_311.n0 111.636
R30 a_209_311.n3 a_209_311.t3 76.731
R31 a_209_311.n4 a_209_311.t0 42.959
R32 a_209_311.n5 a_209_311.n4 27.58
R33 a_209_311.n2 a_209_311.n1 14.386
R34 a_209_311.n4 a_209_311.n3 8.442
R35 VPWR.n3 VPWR.n0 432.494
R36 VPWR.n8 VPWR.t1 376.99
R37 VPWR.n2 VPWR.n1 310.879
R38 VPWR.n0 VPWR.t0 93.809
R39 VPWR.n1 VPWR.t4 63.321
R40 VPWR.n1 VPWR.t2 63.321
R41 VPWR.n0 VPWR.t3 28.516
R42 VPWR.n3 VPWR.n2 5.782
R43 VPWR.n5 VPWR.n4 4.65
R44 VPWR.n7 VPWR.n6 4.65
R45 VPWR.n9 VPWR.n8 4.65
R46 VPWR.n5 VPWR.n3 0.19
R47 VPWR.n7 VPWR.n5 0.119
R48 VPWR.n9 VPWR.n7 0.119
R49 VPWR VPWR.n9 0.02
R50 X.n0 X.t1 172.279
R51 X.n1 X.t0 117.423
R52 X.n1 X.n0 100.727
R53 X.n0 X 4.521
R54 X X.n1 4.184
R55 VPB.t1 VPB.t2 538.629
R56 VPB.t0 VPB.t3 281.152
R57 VPB.t4 VPB.t0 281.152
R58 VPB.t2 VPB.t4 248.598
R59 VPB VPB.t1 189.408
R60 a_296_53.t0 a_296_53.t1 60
R61 C.n0 C.t1 196.548
R62 C.n0 C.t0 148.348
R63 C C.n0 88.331
R64  C 20.448
R65 B.t1 B.t0 403.273
R66 B B.t1 227.513
R67 a_368_53.t0 a_368_53.t1 72.857
C0 VPWR B 0.18fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__and3b_2.ext - technology: sky130A

.subckt sky130_fd_sc_hd__and3b_2 VGND VPWR B X A_N C VNB VPB
X0 a_109_53.t0 A_N.t0 VPWR.t0 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1 X.t3 a_215_311.t4 VGND.t1 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 a_109_53.t1 A_N.t1 VGND.t2 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3 VGND.t3 C.t0 a_373_53.t0 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 VGND.t0 a_215_311.t5 X.t2 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 VPWR.t1 C.t1 a_215_311.t2 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 VPWR.t3 a_215_311.t6 X.t1 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 X.t0 a_215_311.t7 VPWR.t4 VPB.t5 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 a_301_53.t0 a_109_53.t2 a_215_311.t1 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9 a_215_311.t3 B.t0 VPWR.t2 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10 a_373_53.t1 B.t1 a_301_53.t1 VNB.t5 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11 VPWR.t5 a_109_53.t3 a_215_311.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
R0 A_N.n0 A_N.t1 167.093
R1 A_N.n0 A_N.t0 141.386
R2 A_N A_N.n0 107.868
R3  A_N 16.422
R4 VPWR.n13 VPWR.t0 395.643
R5 VPWR.n6 VPWR.n5 308.361
R6 VPWR.n2 VPWR.t3 201.241
R7 VPWR.n1 VPWR.n0 177.914
R8 VPWR.n0 VPWR.t1 96.154
R9 VPWR.n5 VPWR.t2 63.321
R10 VPWR.n5 VPWR.t5 63.321
R11 VPWR.n0 VPWR.t4 25.61
R12 VPWR.n4 VPWR.n3 4.65
R13 VPWR.n8 VPWR.n7 4.65
R14 VPWR.n10 VPWR.n9 4.65
R15 VPWR.n12 VPWR.n11 4.65
R16 VPWR.n14 VPWR.n13 4.65
R17 VPWR.n2 VPWR.n1 3.878
R18 VPWR.n7 VPWR.n6 1.137
R19 VPWR.n4 VPWR.n2 0.227
R20 VPWR.n8 VPWR.n4 0.119
R21 VPWR.n10 VPWR.n8 0.119
R22 VPWR.n12 VPWR.n10 0.119
R23 VPWR.n14 VPWR.n12 0.119
R24 VPWR VPWR.n14 0.022
R25 a_109_53.t0 a_109_53.n1 384.213
R26 a_109_53.n0 a_109_53.t2 186.028
R27 a_109_53.n1 a_109_53.t1 167.505
R28 a_109_53.n0 a_109_53.t3 160.321
R29 a_109_53.n1 a_109_53.n0 96.313
R30 VPB.t1 VPB.t0 556.386
R31 VPB.t2 VPB.t5 287.071
R32 VPB.t3 VPB.t2 281.152
R33 VPB.t5 VPB.t4 248.598
R34 VPB.t0 VPB.t3 248.598
R35 VPB VPB.t1 192.367
R36 a_215_311.t0 a_215_311.n4 392.026
R37 a_215_311.n3 a_215_311.n2 306.984
R38 a_215_311.n0 a_215_311.t6 212.079
R39 a_215_311.n1 a_215_311.t7 212.079
R40 a_215_311.n4 a_215_311.t1 201.922
R41 a_215_311.n0 a_215_311.t5 139.779
R42 a_215_311.n1 a_215_311.t4 139.779
R43 a_215_311.n3 a_215_311.n1 132.875
R44 a_215_311.n2 a_215_311.t3 79.545
R45 a_215_311.n1 a_215_311.n0 61.345
R46 a_215_311.n2 a_215_311.t2 48.587
R47 a_215_311.n4 a_215_311.n3 12.8
R48 VGND.n11 VGND.t2 150.508
R49 VGND.n2 VGND.t0 146.392
R50 VGND.n1 VGND.n0 112.405
R51 VGND.n0 VGND.t3 86.373
R52 VGND.n0 VGND.t1 22.191
R53 VGND.n12 VGND.n11 4.65
R54 VGND.n4 VGND.n3 4.65
R55 VGND.n6 VGND.n5 4.65
R56 VGND.n8 VGND.n7 4.65
R57 VGND.n10 VGND.n9 4.65
R58 VGND.n2 VGND.n1 3.741
R59 VGND.n4 VGND.n2 0.246
R60 VGND.n6 VGND.n4 0.119
R61 VGND.n8 VGND.n6 0.119
R62 VGND.n10 VGND.n8 0.119
R63 VGND.n12 VGND.n10 0.119
R64 VGND VGND.n12 0.022
R65 X.n1 X.n0 146.36
R66 X.n3 X.n2 92.5
R67 X X.n1 44.566
R68 X X.n3 29.284
R69 X.n0 X.t1 26.595
R70 X.n0 X.t0 26.595
R71 X.n2 X.t2 24.923
R72 X.n2 X.t3 24.923
R73 X.n3 X 5.485
R74 X.n1 X 3.708
R75 VNB.t4 VNB.t1 32293.1
R76 VNB VNB.t3 7247.06
R77 VNB.t3 VNB.t2 6211.76
R78 VNB.t5 VNB.t4 2620.59
R79 VNB.t2 VNB.t5 2329.41
R80 VNB.t1 VNB.t0 2030.77
R81 C.n0 C.t0 196.548
R82 C.n0 C.t1 148.348
R83 C C.n0 88.331
R84 C  20.723
R85 a_373_53.t0 a_373_53.t1 72.857
R86 a_301_53.t0 a_301_53.t1 60
R87 B.t0 B.t1 402.004
R88 B B.t0 228.011
C0 X VGND 0.20fF
C1 B VPWR 0.19fF
C2 VPB VPWR 0.10fF
C3 X VPWR 0.33fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__and3b_4.ext - technology: sky130A

.subckt sky130_fd_sc_hd__and3b_4 A_N X C B VGND VPWR VNB VPB
X0 a_98_199.t1 A_N.t0 VGND.t2 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1 X.t7 a_56_297.t4 VGND.t3 VNB.t5 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 VPWR.t7 a_56_297.t5 X.t3 VPB.t7 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 VGND.t4 a_56_297.t6 X.t6 VNB.t6 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 VPWR.t2 a_98_199.t2 a_56_297.t2 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 VPWR.t6 a_56_297.t7 X.t2 VPB.t6 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 VGND.t5 a_56_297.t8 X.t5 VNB.t7 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 a_257_47.t1 B.t0 a_152_47.t1 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 X.t4 a_56_297.t9 VGND.t0 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 X.t1 a_56_297.t10 VPWR.t5 VPB.t5 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 a_152_47.t0 a_98_199.t3 a_56_297.t3 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 VPWR.t0 C.t0 a_56_297.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 a_98_199.t0 A_N.t1 VPWR.t3 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13 a_56_297.t1 B.t1 VPWR.t1 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14 VGND.t1 C.t1 a_257_47.t0 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X15 X.t0 a_56_297.t11 VPWR.t4 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
R0 A_N.n0 A_N.t1 224.933
R1 A_N.n0 A_N.t0 131.746
R2 A_N.n1 A_N.n0 76
R3  A_N.n1 13.028
R4 A_N.n1 A_N 2.514
R5 VGND.n5 VGND.n4 110.811
R6 VGND.n3 VGND.n2 106.463
R7 VGND.n1 VGND.n0 106.463
R8 VGND.n4 VGND.t2 62.857
R9 VGND.n0 VGND.t1 51.692
R10 VGND.n0 VGND.t0 26.769
R11 VGND.n4 VGND.t4 25.846
R12 VGND.n2 VGND.t3 25.846
R13 VGND.n2 VGND.t5 25.846
R14 VGND.n5 VGND.n3 4.995
R15 VGND.n7 VGND.n6 4.65
R16 VGND.n8 VGND.n1 3.627
R17 VGND VGND.n8 0.471
R18 VGND.n7 VGND.n5 0.4
R19 VGND.n8 VGND.n7 0.148
R20 a_98_199.t0 a_98_199.n1 359.537
R21 a_98_199.n1 a_98_199.n0 313.44
R22 a_98_199.n0 a_98_199.t2 241.534
R23 a_98_199.n1 a_98_199.t1 216.5
R24 a_98_199.n0 a_98_199.t3 169.234
R25 VNB VNB.t3 7156.04
R26 VNB.t1 VNB.t0 2780.22
R27 VNB.t3 VNB.t2 2538.46
R28 VNB.t6 VNB.t4 2424.58
R29 VNB.t5 VNB.t6 2079.12
R30 VNB.t7 VNB.t5 2079.12
R31 VNB.t0 VNB.t7 2079.12
R32 VNB.t2 VNB.t1 1837.36
R33 a_56_297.n11 a_56_297.n10 345.975
R34 a_56_297.n0 a_56_297.t2 237.291
R35 a_56_297.n1 a_56_297.t5 212.079
R36 a_56_297.n2 a_56_297.t11 212.079
R37 a_56_297.n4 a_56_297.t7 212.079
R38 a_56_297.n7 a_56_297.t10 212.079
R39 a_56_297.n5 a_56_297.t8 139.779
R40 a_56_297.n1 a_56_297.t6 139.779
R41 a_56_297.n2 a_56_297.t4 139.779
R42 a_56_297.n7 a_56_297.t9 139.779
R43 a_56_297.n10 a_56_297.n0 110.03
R44 a_56_297.n6 a_56_297.n3 88.991
R45 a_56_297.n0 a_56_297.t3 78.34
R46 a_56_297.n6 a_56_297.n5 76
R47 a_56_297.n9 a_56_297.n8 76
R48 a_56_297.n2 a_56_297.n1 62.806
R49 a_56_297.n11 a_56_297.t1 31.52
R50 a_56_297.t0 a_56_297.n11 27.58
R51 a_56_297.n3 a_56_297.n2 13.145
R52 a_56_297.n8 a_56_297.n7 13.145
R53 a_56_297.n9 a_56_297.n6 12.991
R54 a_56_297.n10 a_56_297.n9 9.743
R55 a_56_297.n5 a_56_297.n4 1.46
R56 X.n2 X.n1 356.5
R57 X.n2 X.n0 292.5
R58 X.n5 X.n4 140.36
R59 X.n5 X.n3 49.316
R60 X.n6 X.n2 39.691
R61 X.n1 X.t1 29.55
R62 X.n1 X.t2 27.58
R63 X.n0 X.t3 27.58
R64 X.n0 X.t0 27.58
R65 X.n4 X.t5 25.846
R66 X.n4 X.t4 25.846
R67 X.n3 X.t6 25.846
R68 X.n3 X.t7 25.846
R69 X X.n5 6.956
R70 X X.n6 3.864
R71 X.n6 X 1.947
R72 VPWR.n3 VPWR.n2 459.425
R73 VPWR.n7 VPWR.n6 306.463
R74 VPWR.n1 VPWR.n0 306.255
R75 VPWR.n12 VPWR.n11 292.5
R76 VPWR.n2 VPWR.t3 103.19
R77 VPWR.n11 VPWR.t2 40.385
R78 VPWR.n6 VPWR.t5 35.46
R79 VPWR.n6 VPWR.t0 34.475
R80 VPWR.n2 VPWR.t7 33.518
R81 VPWR.n11 VPWR.t1 33.49
R82 VPWR.n0 VPWR.t4 26.595
R83 VPWR.n0 VPWR.t6 26.595
R84 VPWR.n14 VPWR.n13 4.65
R85 VPWR.n5 VPWR.n4 4.65
R86 VPWR.n8 VPWR.n7 4.65
R87 VPWR.n10 VPWR.n9 4.65
R88 VPWR.n3 VPWR.n1 4.618
R89 VPWR.n13 VPWR.n12 4.467
R90 VPWR.n5 VPWR.n3 0.4
R91 VPWR.n15 VPWR.n14 0.132
R92 VPWR VPWR.n15 0.129
R93 VPWR.n8 VPWR.n5 0.119
R94 VPWR.n10 VPWR.n8 0.119
R95 VPWR.n14 VPWR.n10 0.119
R96 VPB VPB.t2 319.626
R97 VPB.t2 VPB.t1 310.747
R98 VPB.t7 VPB.t3 301.869
R99 VPB.t0 VPB.t5 298.909
R100 VPB.t1 VPB.t0 266.355
R101 VPB.t5 VPB.t6 260.436
R102 VPB.t4 VPB.t7 254.517
R103 VPB.t6 VPB.t4 248.598
R104 B.n0 B.t1 237.326
R105 B.n0 B.t0 165.026
R106 B B.n0 79.274
R107  B 20.241
R108 a_152_47.t0 a_152_47.t1 69.23
R109 a_257_47.t0 a_257_47.t1 42.461
R110 C.n0 C.t0 241.534
R111 C.n0 C.t1 169.234
R112 C C.n0 79.895
C0 VGND VPWR 0.10fF
C1 X VGND 0.21fF
C2 X A_N 0.13fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__and4_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__and4_1 X C A B D VGND VPWR VNB VPB
X0 a_27_47.t4 C.t0 VPWR.t4 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1 a_197_47.t0 B.t0 a_109_47.t1 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 X.t1 a_27_47.t5 VPWR.t2 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 a_303_47.t1 C.t1 a_197_47.t1 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 a_27_47.t3 A.t0 VPWR.t3 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 VPWR.t1 D.t0 a_27_47.t1 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 VGND.t1 D.t1 a_303_47.t0 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7 VPWR.t0 B.t1 a_27_47.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 X.t0 a_27_47.t6 VGND.t0 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 a_109_47.t0 A.t1 a_27_47.t2 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
R0 C.n0 C.t0 334.721
R1 C.n0 C.t1 206.188
R2 C C.n0 78.346
R3 VPWR.n6 VPWR.t3 370.34
R4 VPWR.n2 VPWR.n1 307.239
R5 VPWR.n3 VPWR.n0 167.901
R6 VPWR.n0 VPWR.t1 117.449
R7 VPWR.n1 VPWR.t4 86.773
R8 VPWR.n1 VPWR.t0 86.773
R9 VPWR.n0 VPWR.t2 42.355
R10 VPWR.n5 VPWR.n4 4.65
R11 VPWR.n7 VPWR.n6 4.65
R12 VPWR.n3 VPWR.n2 3.75
R13 VPWR.n5 VPWR.n3 0.159
R14 VPWR.n7 VPWR.n5 0.119
R15 VPWR VPWR.n7 0.022
R16 a_27_47.n2 a_27_47.n1 329.364
R17 a_27_47.n4 a_27_47.n3 325.012
R18 a_27_47.n0 a_27_47.t5 230.791
R19 a_27_47.n3 a_27_47.t2 222.541
R20 a_27_47.n0 a_27_47.t6 158.491
R21 a_27_47.n2 a_27_47.n0 133.724
R22 a_27_47.t0 a_27_47.n4 82.083
R23 a_27_47.n4 a_27_47.t3 82.083
R24 a_27_47.n1 a_27_47.t1 65.666
R25 a_27_47.n1 a_27_47.t4 65.666
R26 a_27_47.n3 a_27_47.n2 64.752
R27 VPB.t1 VPB.t2 491.277
R28 VPB.t0 VPB.t4 307.788
R29 VPB.t3 VPB.t0 295.95
R30 VPB.t4 VPB.t1 254.517
R31 VPB VPB.t3 192.367
R32 B.n0 B.t1 334.721
R33 B.n0 B.t0 206.188
R34 B B.n0 90.445
R35 a_109_47.t0 a_109_47.t1 82.857
R36 a_197_47.t0 a_197_47.t1 108.571
R37 VNB VNB.t2 6470.59
R38 VNB.t0 VNB.t1 4274.85
R39 VNB.t3 VNB.t4 3429.41
R40 VNB.t4 VNB.t0 3105.88
R41 VNB.t2 VNB.t3 2847.06
R42 X.n2 X.n1 297.582
R43 X.n5 X.n2 292.5
R44 X.n3 X.t0 83.131
R45 X.n2 X.t1 26.595
R46 X X.n4 14.769
R47 X X.n0 10.584
R48 X.n5 X 10.584
R49 X X.n3 6.902
R50 X X.n0 6.153
R51 X X.n5 6.153
R52 X.n3 X 5.55
R53 X.n1 X 3.938
R54 X.n1 X 3.011
R55 X.n4 X 1.969
R56 X.n4 X 1.505
R57 a_303_47.t0 a_303_47.t1 94.285
R58 A.n0 A.t0 323.341
R59 A.n0 A.t1 194.808
R60 A A.n0 76.928
R61 D.n0 D.t0 330.119
R62 D.n0 D.t1 201.586
R63 D D.n0 78.514
R64 VGND.n0 VGND.t1 108.504
R65 VGND VGND.n0 72.066
R66 VGND.n0 VGND.t0 38.769
C0 VGND D 0.12fF
C1 X VGND 0.14fF
C2 VPWR X 0.15fF
C3 C D 0.25fF
C4 B C 0.23fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__and4_2.ext - technology: sky130A

.subckt sky130_fd_sc_hd__and4_2 X C A B D VGND VPWR VNB VPB
X0 VGND.t2 a_27_47.t5 X.t3 VNB.t5 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 VGND.t0 D.t0 a_304_47.t0 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 X.t1 a_27_47.t6 VPWR.t4 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 a_198_47.t0 B.t0 a_109_47.t1 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 a_27_47.t3 C.t0 VPWR.t2 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 VPWR.t3 a_27_47.t7 X.t0 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 a_304_47.t1 C.t1 a_198_47.t1 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7 a_27_47.t0 A.t0 VPWR.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 VPWR.t1 D.t1 a_27_47.t2 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9 X.t2 a_27_47.t8 VGND.t1 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 VPWR.t5 B.t1 a_27_47.t4 VPB.t5 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11 a_109_47.t0 A.t1 a_27_47.t1 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
R0 a_27_47.n3 a_27_47.n2 329.364
R1 a_27_47.n5 a_27_47.n4 325.012
R2 a_27_47.n4 a_27_47.t1 222.735
R3 a_27_47.n0 a_27_47.t7 212.079
R4 a_27_47.n1 a_27_47.t6 212.079
R5 a_27_47.n3 a_27_47.n1 152.354
R6 a_27_47.n0 a_27_47.t5 139.779
R7 a_27_47.n1 a_27_47.t8 139.779
R8 a_27_47.t0 a_27_47.n5 84.428
R9 a_27_47.n5 a_27_47.t4 82.083
R10 a_27_47.n1 a_27_47.n0 70.109
R11 a_27_47.n2 a_27_47.t2 65.666
R12 a_27_47.n2 a_27_47.t3 65.666
R13 a_27_47.n4 a_27_47.n3 64.752
R14 X.n4 X.n3 292.5
R15 X.n3 X.n2 147.091
R16 X X.n0 94.219
R17 X.n1 X.n0 92.5
R18 X.n3 X.t0 38.415
R19 X.n0 X.t3 36
R20 X.n3 X.t1 26.595
R21 X.n0 X.t2 24.923
R22 X.n6 X 21.942
R23 X.n1 X 11.271
R24 X.n2 X 10.551
R25 X.n5 X.n4 6.304
R26 X.n4 X 4.776
R27 X X.n5 3.657
R28 X X.n6 2.925
R29 X.n2 X 2.402
R30 X.n5 X 1.91
R31 X X.n1 1.719
R32 X.n6 X 1.528
R33 VGND.n0 VGND.t0 121.48
R34 VGND.n1 VGND.t2 100.6
R35 VGND.n1 VGND.n0 80.058
R36 VGND.n0 VGND.t1 15.993
R37 VGND VGND.n1 0.683
R38 VNB VNB.t0 6438.23
R39 VNB.t2 VNB.t4 3960.57
R40 VNB.t1 VNB.t3 3429.41
R41 VNB.t3 VNB.t2 3105.88
R42 VNB.t0 VNB.t1 2879.41
R43 VNB.t4 VNB.t5 2320.88
R44 D.n0 D.t1 330.119
R45 D.n0 D.t0 201.586
R46 D D.n0 78.707
R47  D 16.738
R48 a_304_47.t0 a_304_47.t1 94.285
R49 VPWR.n12 VPWR.t0 370.56
R50 VPWR.n8 VPWR.n7 307.239
R51 VPWR.n2 VPWR.t3 200.693
R52 VPWR.n1 VPWR.n0 164.214
R53 VPWR.n0 VPWR.t1 104.644
R54 VPWR.n7 VPWR.t2 86.773
R55 VPWR.n7 VPWR.t5 86.773
R56 VPWR.n0 VPWR.t4 42.355
R57 VPWR.n4 VPWR.n3 4.65
R58 VPWR.n6 VPWR.n5 4.65
R59 VPWR.n9 VPWR.n8 4.65
R60 VPWR.n11 VPWR.n10 4.65
R61 VPWR.n13 VPWR.n12 4.65
R62 VPWR.n2 VPWR.n1 4.016
R63 VPWR.n4 VPWR.n2 0.222
R64 VPWR.n6 VPWR.n4 0.119
R65 VPWR.n9 VPWR.n6 0.119
R66 VPWR.n11 VPWR.n9 0.119
R67 VPWR.n13 VPWR.n11 0.119
R68 VPWR VPWR.n13 0.02
R69 VPB.t1 VPB.t4 452.803
R70 VPB.t5 VPB.t2 307.788
R71 VPB.t0 VPB.t5 298.909
R72 VPB.t4 VPB.t3 284.112
R73 VPB.t2 VPB.t1 254.517
R74 VPB VPB.t0 189.408
R75 B.n0 B.t1 334.721
R76 B.n0 B.t0 206.188
R77 B B.n0 90.242
R78 a_109_47.t0 a_109_47.t1 84.285
R79 a_198_47.t0 a_198_47.t1 108.571
R80 C.n0 C.t0 334.721
R81 C.n0 C.t1 206.188
R82 C C.n0 78.346
R83 A.n0 A.t0 323.548
R84 A.n0 A.t1 195.015
R85 A.n1 A.n0 76
R86  A 21.229
R87 A.n1  17.795
R88 A A.n1 3.434
C0 C D 0.24fF
C1 VGND D 0.11fF
C2 B C 0.23fF
C3 X VGND 0.18fF
C4 VPWR X 0.27fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__and4_4.ext - technology: sky130A

.subckt sky130_fd_sc_hd__and4_4 X C A B D VGND VPWR VNB VPB
X0 VPWR.t6 a_27_47.t5 X.t0 VPB.t6 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 X.t7 a_27_47.t6 VPWR.t5 VPB.t5 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 a_188_47.t1 B.t0 a_109_47.t1 VNB.t6 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 VPWR.t4 a_27_47.t7 X.t6 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 VGND.t4 D.t0 a_285_47.t1 VNB.t7 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 VPWR.t7 D.t1 a_27_47.t4 VPB.t7 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 X.t5 a_27_47.t8 VPWR.t3 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 VGND.t3 a_27_47.t9 X.t4 VNB.t5 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 VPWR.t2 B.t1 a_27_47.t3 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 X.t3 a_27_47.t10 VGND.t2 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 X.t2 a_27_47.t11 VGND.t1 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 a_27_47.t2 C.t0 VPWR.t1 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 VGND.t0 a_27_47.t12 X.t1 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 a_27_47.t0 A.t0 VPWR.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14 a_285_47.t0 C.t1 a_188_47.t0 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X15 a_109_47.t0 A.t1 a_27_47.t1 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
R0 a_27_47.n11 a_27_47.t1 243.885
R1 a_27_47.n0 a_27_47.t5 212.079
R2 a_27_47.n2 a_27_47.t6 212.079
R3 a_27_47.n5 a_27_47.t7 212.079
R4 a_27_47.n6 a_27_47.t8 212.079
R5 a_27_47.n10 a_27_47.n9 177.361
R6 a_27_47.n12 a_27_47.n11 169.235
R7 a_27_47.n0 a_27_47.t12 139.779
R8 a_27_47.n2 a_27_47.t11 139.779
R9 a_27_47.n5 a_27_47.t9 139.779
R10 a_27_47.n6 a_27_47.t10 139.779
R11 a_27_47.n4 a_27_47.n1 94.921
R12 a_27_47.n10 a_27_47.n8 90.743
R13 a_27_47.n8 a_27_47.n7 76
R14 a_27_47.n4 a_27_47.n3 76
R15 a_27_47.n11 a_27_47.n10 59.857
R16 a_27_47.n9 a_27_47.t4 58.115
R17 a_27_47.n7 a_27_47.n6 48.2
R18 a_27_47.n1 a_27_47.n0 36.515
R19 a_27_47.n9 a_27_47.t2 26.595
R20 a_27_47.n12 a_27_47.t3 26.595
R21 a_27_47.t0 a_27_47.n12 26.595
R22 a_27_47.n3 a_27_47.n2 24.83
R23 a_27_47.n8 a_27_47.n4 18.921
R24 a_27_47.n7 a_27_47.n5 13.145
R25 X.n2 X.n1 224.473
R26 X.n5 X.n4 172.311
R27 X.n2 X.n0 168.571
R28 X.n5 X.n3 109.064
R29 X X.n5 27.648
R30 X.n1 X.t6 26.595
R31 X.n1 X.t5 26.595
R32 X.n0 X.t0 26.595
R33 X.n0 X.t7 26.595
R34 X.n4 X.t4 24.923
R35 X.n4 X.t3 24.923
R36 X.n3 X.t1 24.923
R37 X.n3 X.t2 24.923
R38 X X.n2 17.723
R39 VPWR.n2 VPWR.t6 194.747
R40 VPWR.n15 VPWR.t0 194.002
R41 VPWR.n1 VPWR.n0 169.933
R42 VPWR.n11 VPWR.n10 163.438
R43 VPWR.n6 VPWR.n5 163.438
R44 VPWR.n5 VPWR.t7 36.445
R45 VPWR.n10 VPWR.t1 30.535
R46 VPWR.n10 VPWR.t2 30.535
R47 VPWR.n5 VPWR.t3 28.565
R48 VPWR.n0 VPWR.t5 26.595
R49 VPWR.n0 VPWR.t4 26.595
R50 VPWR.n4 VPWR.n3 4.65
R51 VPWR.n7 VPWR.n6 4.65
R52 VPWR.n9 VPWR.n8 4.65
R53 VPWR.n12 VPWR.n11 4.65
R54 VPWR.n14 VPWR.n13 4.65
R55 VPWR.n16 VPWR.n15 4.65
R56 VPWR.n2 VPWR.n1 3.704
R57 VPWR.n4 VPWR.n2 0.269
R58 VPWR.n7 VPWR.n4 0.119
R59 VPWR.n9 VPWR.n7 0.119
R60 VPWR.n12 VPWR.n9 0.119
R61 VPWR.n14 VPWR.n12 0.119
R62 VPWR.n16 VPWR.n14 0.119
R63 VPWR VPWR.n16 0.02
R64 VPB.t1 VPB.t7 343.302
R65 VPB.t7 VPB.t3 284.112
R66 VPB.t2 VPB.t1 272.274
R67 VPB.t5 VPB.t6 248.598
R68 VPB.t4 VPB.t5 248.598
R69 VPB.t3 VPB.t4 248.598
R70 VPB.t0 VPB.t2 248.598
R71 VPB VPB.t0 189.408
R72 B.n0 B.t1 241.534
R73 B.n0 B.t0 169.234
R74  B.n0 77.983
R75  B 12.259
R76 a_109_47.t0 a_109_47.t1 45.23
R77 a_188_47.t0 a_188_47.t1 61.846
R78 VNB VNB.t0 6053.91
R79 VNB.t1 VNB.t7 2828.57
R80 VNB.t6 VNB.t1 2345.05
R81 VNB.t7 VNB.t4 2296.7
R82 VNB.t3 VNB.t2 2030.77
R83 VNB.t5 VNB.t3 2030.77
R84 VNB.t4 VNB.t5 2030.77
R85 VNB.t0 VNB.t6 1909.89
R86 D.n0 D.t1 241.534
R87 D.n0 D.t0 164.95
R88 D D.n0 101.645
R89 a_285_47.t0 a_285_47.t1 80.307
R90 VGND.n4 VGND.t0 192.14
R91 VGND.n1 VGND.n0 108.396
R92 VGND.n3 VGND.n2 107.433
R93 VGND.n0 VGND.t4 33.23
R94 VGND.n0 VGND.t2 26.769
R95 VGND.n2 VGND.t1 24.923
R96 VGND.n2 VGND.t3 24.923
R97 VGND.n6 VGND.n5 4.65
R98 VGND.n7 VGND.n1 4.097
R99 VGND.n4 VGND.n3 3.704
R100 VGND VGND.n7 0.482
R101 VGND.n6 VGND.n4 0.269
R102 VGND.n7 VGND.n6 0.135
R103 C.n0 C.t0 233.868
R104 C.n0 C.t1 161.568
R105  C.n0 78.47
R106  C 15.27
R107 A.n0 A.t0 230.361
R108 A.n0 A.t1 158.061
R109 A A.n0 79.434
R110  A 21.229
C0 C D 0.13fF
C1 B C 0.20fF
C2 X VGND 0.34fF
C3 VPWR X 0.53fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__and4b_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__and4b_1 VGND VPWR C A_N X D B VNB VPB
X0 a_297_47.t1 a_27_47.t2 a_193_413.t3 VNB.t5 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1 a_369_47.t0 B.t0 a_297_47.t0 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 VPWR.t1 D.t0 a_193_413.t1 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3 X.t0 a_193_413.t5 VGND.t0 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 VPWR.t5 A_N.t0 a_27_47.t1 VPB.t5 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 VGND.t1 D.t1 a_469_47.t0 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 X.t1 a_193_413.t6 VPWR.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 VPWR.t2 B.t1 a_193_413.t2 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 a_193_413.t0 C.t0 VPWR.t3 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9 a_193_413.t4 a_27_47.t3 VPWR.t4 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10 a_469_47.t1 C.t1 a_369_47.t1 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11 VGND.t2 A_N.t1 a_27_47.t0 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
R0 a_27_47.n1 a_27_47.t1 455.927
R1 a_27_47.n0 a_27_47.t3 334.721
R2 a_27_47.n0 a_27_47.t2 302.224
R3 a_27_47.t0 a_27_47.n1 201.168
R4 a_27_47.n1 a_27_47.n0 76
R5 a_193_413.n2 a_193_413.n1 311.7
R6 a_193_413.n4 a_193_413.n3 311.7
R7 a_193_413.n0 a_193_413.t6 241.534
R8 a_193_413.n2 a_193_413.t3 237.382
R9 a_193_413.n0 a_193_413.t5 169.234
R10 a_193_413.n3 a_193_413.n0 167.322
R11 a_193_413.n1 a_193_413.t4 126.642
R12 a_193_413.n3 a_193_413.n2 97.129
R13 a_193_413.n1 a_193_413.t2 93.809
R14 a_193_413.t0 a_193_413.n4 84.428
R15 a_193_413.n4 a_193_413.t1 63.321
R16 a_297_47.t0 a_297_47.t1 60
R17 VNB VNB.t3 6470.59
R18 VNB.t3 VNB.t5 6082.35
R19 VNB.t4 VNB.t1 3235.29
R20 VNB.t1 VNB.t2 2847.06
R21 VNB.t2 VNB.t0 2345.21
R22 VNB.t5 VNB.t4 2329.41
R23 B.n0 B.t1 295.43
R24 B.n0 B.t0 237.59
R25 B.n1 B.n0 76
R26 B B.n1 8
R27 B.n1 B 7.542
R28 a_369_47.t0 a_369_47.t1 100
R29 D.n0 D.t0 334.721
R30 D.n0 D.t1 206.188
R31 D.n1 D.n0 76
R32 D.n1 D 10.729
R33 D D.n1 2.07
R34 VPWR.n3 VPWR.n2 311.951
R35 VPWR.n11 VPWR.n10 307.239
R36 VPWR.n5 VPWR.n4 292.5
R37 VPWR.n1 VPWR.n0 292.5
R38 VPWR.n2 VPWR.t1 77.392
R39 VPWR.n0 VPWR.t3 63.321
R40 VPWR.n4 VPWR.t2 63.321
R41 VPWR.n10 VPWR.t4 63.321
R42 VPWR.n10 VPWR.t5 63.321
R43 VPWR.n2 VPWR.t0 41.041
R44 VPWR.n7 VPWR.n6 4.65
R45 VPWR.n9 VPWR.n8 4.65
R46 VPWR.n3 VPWR.n1 4.153
R47 VPWR.n12 VPWR.n11 3.932
R48 VPWR.n6 VPWR.n5 2.427
R49 VPWR.n7 VPWR.n3 0.221
R50 VPWR.n12 VPWR.n9 0.137
R51 VPWR VPWR.n12 0.123
R52 VPWR.n9 VPWR.n7 0.119
R53 VPB.t2 VPB.t3 449.844
R54 VPB.t4 VPB.t2 366.978
R55 VPB.t1 VPB.t0 281.152
R56 VPB.t3 VPB.t1 275.233
R57 VPB.t5 VPB.t4 248.598
R58 VPB VPB.t5 192.367
R59 VGND.n1 VGND.t2 149.228
R60 VGND.n1 VGND.n0 111.204
R61 VGND.n0 VGND.t0 48.285
R62 VGND.n0 VGND.t1 38.571
R63 VGND VGND.n1 0.143
R64 X.n1 X.t1 538.75
R65 X X.t1 442.957
R66 X.n0 X.t0 83.131
R67 X.n1 X.n0 68.483
R68 X X.n1 6.153
R69 X.n0 X 5.55
R70 A_N.n0 A_N.t0 323.341
R71 A_N.n0 A_N.t1 194.808
R72 A_N.n1 A_N.n0 76
R73 A_N.n1 A_N 9.994
R74 A_N A_N.n1 1.928
R75 a_469_47.t0 a_469_47.t1 82.857
R76 C.n0 C.t0 334.721
R77 C.n0 C.t1 206.188
R78 C.n1 C.n0 76
R79 C.n1 C 13.511
R80 C C.n1 2.607
C0 C B 0.20fF
C1 C D 0.25fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__and4b_2.ext - technology: sky130A

.subckt sky130_fd_sc_hd__and4b_2 VPWR VGND X A_N D C B VNB VPB
X0 VPWR.t6 a_193_413.t5 X.t2 VPB.t6 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_297_47.t0 a_27_413.t2 a_193_413.t0 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 a_369_47.t0 B.t0 a_297_47.t1 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3 X.t3 a_193_413.t6 VGND.t3 VNB.t6 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 VPWR.t3 D.t0 a_193_413.t3 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 VPWR.t0 A_N.t0 a_27_413.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 VGND.t1 D.t1 a_469_47.t1 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7 VGND.t2 a_193_413.t7 X.t0 VNB.t5 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 VPWR.t4 B.t1 a_193_413.t4 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9 a_193_413.t2 C.t0 VPWR.t2 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10 X.t1 a_193_413.t8 VPWR.t5 VPB.t5 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 a_193_413.t1 a_27_413.t3 VPWR.t1 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12 a_469_47.t0 C.t1 a_369_47.t1 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13 a_27_413.t1 A_N.t1 VGND.t0 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
R0 a_193_413.n3 a_193_413.n0 315.088
R1 a_193_413.n5 a_193_413.n4 312.314
R2 a_193_413.t0 a_193_413.n5 236.118
R3 a_193_413.n1 a_193_413.t5 212.079
R4 a_193_413.n2 a_193_413.t8 212.079
R5 a_193_413.n3 a_193_413.n2 170.506
R6 a_193_413.n4 a_193_413.t4 157.13
R7 a_193_413.n1 a_193_413.t7 139.779
R8 a_193_413.n2 a_193_413.t6 139.779
R9 a_193_413.n5 a_193_413.n3 84.705
R10 a_193_413.n0 a_193_413.t2 84.428
R11 a_193_413.n2 a_193_413.n1 66.457
R12 a_193_413.n0 a_193_413.t3 63.321
R13 a_193_413.n4 a_193_413.t1 63.321
R14 X.n4 X.n3 146.401
R15 X X.n0 93.033
R16 X.n3 X.t1 33.49
R17 X.n0 X.t3 31.384
R18 X.n3 X.t2 26.595
R19 X.n0 X.t0 24.923
R20 X X.n2 20.782
R21 X.n4 X 15.897
R22 X X.n1 11.894
R23 X X.n4 5.157
R24 X.n2 X 4.876
R25 X.n1 X 2.133
R26 X.n2 X 1.828
R27 X.n1 X 1.551
R28 VPWR.n1 VPWR.n0 307.239
R29 VPWR.n16 VPWR.n15 307.239
R30 VPWR.n10 VPWR.n9 292.5
R31 VPWR.n6 VPWR.n5 292.5
R32 VPWR.n2 VPWR.t6 194.496
R33 VPWR.n0 VPWR.t3 91.464
R34 VPWR.n5 VPWR.t2 63.321
R35 VPWR.n9 VPWR.t4 63.321
R36 VPWR.n15 VPWR.t1 63.321
R37 VPWR.n15 VPWR.t0 63.321
R38 VPWR.n0 VPWR.t5 27.955
R39 VPWR.n4 VPWR.n3 4.65
R40 VPWR.n8 VPWR.n7 4.65
R41 VPWR.n12 VPWR.n11 4.65
R42 VPWR.n14 VPWR.n13 4.65
R43 VPWR.n17 VPWR.n16 3.932
R44 VPWR.n2 VPWR.n1 3.787
R45 VPWR.n11 VPWR.n10 2.56
R46 VPWR.n4 VPWR.n2 0.256
R47 VPWR.n7 VPWR.n6 0.232
R48 VPWR.n17 VPWR.n14 0.137
R49 VPWR VPWR.n17 0.121
R50 VPWR.n8 VPWR.n4 0.119
R51 VPWR.n12 VPWR.n8 0.119
R52 VPWR.n14 VPWR.n12 0.119
R53 VPB.t4 VPB.t2 449.844
R54 VPB.t1 VPB.t4 366.978
R55 VPB.t3 VPB.t5 284.112
R56 VPB.t2 VPB.t3 275.233
R57 VPB.t5 VPB.t6 269.314
R58 VPB.t0 VPB.t1 248.598
R59 VPB VPB.t0 189.408
R60 a_27_413.t0 a_27_413.n1 457.278
R61 a_27_413.n0 a_27_413.t3 334.721
R62 a_27_413.n0 a_27_413.t2 305.801
R63 a_27_413.n1 a_27_413.t1 178.209
R64 a_27_413.n1 a_27_413.n0 76
R65 a_297_47.t0 a_297_47.t1 60
R66 VNB VNB.t0 6438.23
R67 VNB.t0 VNB.t2 6082.35
R68 VNB.t4 VNB.t1 3235.29
R69 VNB.t1 VNB.t3 2879.41
R70 VNB.t3 VNB.t6 2355.55
R71 VNB.t2 VNB.t4 2329.41
R72 VNB.t6 VNB.t5 2200
R73 B.n1 B.t0 255.46
R74 B.n0 B.t1 191.8
R75 B B.n0 83.854
R76 B.n2 B.n1 76
R77 B B.n2 11.927
R78 B.n2 B 7.854
R79 a_369_47.t0 a_369_47.t1 100
R80 VGND.n2 VGND.t2 194.076
R81 VGND.n13 VGND.t0 145.81
R82 VGND.n1 VGND.n0 107.239
R83 VGND.n0 VGND.t3 47.78
R84 VGND.n0 VGND.t1 38.571
R85 VGND.n14 VGND.n13 4.65
R86 VGND.n4 VGND.n3 4.65
R87 VGND.n6 VGND.n5 4.65
R88 VGND.n8 VGND.n7 4.65
R89 VGND.n10 VGND.n9 4.65
R90 VGND.n12 VGND.n11 4.65
R91 VGND.n2 VGND.n1 3.933
R92 VGND.n4 VGND.n2 0.233
R93 VGND.n6 VGND.n4 0.119
R94 VGND.n8 VGND.n6 0.119
R95 VGND.n10 VGND.n8 0.119
R96 VGND.n12 VGND.n10 0.119
R97 VGND.n14 VGND.n12 0.119
R98 VGND VGND.n14 0.02
R99 D.n0 D.t0 334.721
R100 D.n0 D.t1 206.188
R101 D.n1 D.n0 76
R102 D.n1 D 11.054
R103  D.n1 2.133
R104 A_N.n0 A_N.t0 323.548
R105 A_N.n0 A_N.t1 195.015
R106 A_N.n1 A_N.n0 76
R107 A_N.n1 A_N 18.24
R108 A_N A_N.n1 3.52
R109 a_469_47.t0 a_469_47.t1 84.285
R110 C.n0 C.t0 332.69
R111 C.n0 C.t1 204.157
R112 C.n1 C.n0 76
R113 C  13.815
R114 C.n1  11.58
R115  C.n1 2.234
C0 X VGND 0.18fF
C1 VPWR X 0.23fF
C2 C D 0.26fF
C3 B C 0.20fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__and4b_4.ext - technology: sky130A

.subckt sky130_fd_sc_hd__and4b_4 X D C B A_N VGND VPWR VNB VPB
X0 VPWR.t5 a_174_21.t5 X.t2 VPB.t5 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 X.t1 a_174_21.t6 VPWR.t4 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 a_815_47.t1 B.t0 a_701_47.t1 VNB.t6 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 VPWR.t3 a_174_21.t7 X.t0 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 VPWR.t1 C.t0 a_174_21.t1 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 a_174_21.t2 a_27_47.t2 a_815_47.t0 VNB.t5 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 X.t3 a_174_21.t8 VPWR.t2 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 VPWR.t7 A_N.t0 a_27_47.t0 VPB.t7 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 a_701_47.t0 C.t1 a_617_47.t0 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 a_174_21.t4 D.t0 VPWR.t8 VPB.t8 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 a_174_21.t0 B.t1 VPWR.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 VPWR.t6 a_27_47.t3 a_174_21.t3 VPB.t6 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 X.t7 a_174_21.t9 VGND.t5 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 X.t6 a_174_21.t10 VGND.t4 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14 a_617_47.t1 D.t1 VGND.t1 VNB.t8 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X15 VGND.t3 a_174_21.t11 X.t5 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X16 VGND.t2 a_174_21.t12 X.t4 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X17 VGND.t0 A_N.t1 a_27_47.t1 VNB.t7 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
R0 a_174_21.n11 a_174_21.n10 379.841
R1 a_174_21.n10 a_174_21.n0 292.5
R2 a_174_21.n9 a_174_21.t2 273.45
R3 a_174_21.n7 a_174_21.t5 212.079
R4 a_174_21.n1 a_174_21.t6 212.079
R5 a_174_21.n4 a_174_21.t7 212.079
R6 a_174_21.n3 a_174_21.t8 212.079
R7 a_174_21.n7 a_174_21.t12 139.779
R8 a_174_21.n1 a_174_21.t10 139.779
R9 a_174_21.n4 a_174_21.t11 139.779
R10 a_174_21.n3 a_174_21.t9 139.779
R11 a_174_21.n6 a_174_21.n5 101.6
R12 a_174_21.n8 a_174_21.n7 87.684
R13 a_174_21.n10 a_174_21.n9 79.435
R14 a_174_21.n6 a_174_21.n2 76
R15 a_174_21.n4 a_174_21.n3 61.345
R16 a_174_21.t0 a_174_21.n11 60.085
R17 a_174_21.n5 a_174_21.n4 35.054
R18 a_174_21.n0 a_174_21.t1 26.595
R19 a_174_21.n0 a_174_21.t4 26.595
R20 a_174_21.n11 a_174_21.t3 26.595
R21 a_174_21.n8 a_174_21.n6 25.6
R22 a_174_21.n2 a_174_21.n1 23.369
R23 a_174_21.n9 a_174_21.n8 13.552
R24 X.n2 X.n0 347.841
R25 X.n2 X.n1 292.5
R26 X.n5 X.n3 165.158
R27 X.n5 X.n4 113.702
R28 X.n0 X.t2 26.595
R29 X.n0 X.t1 26.595
R30 X.n1 X.t0 26.595
R31 X.n1 X.t3 26.595
R32 X.n3 X.t4 24.923
R33 X.n3 X.t6 24.923
R34 X.n4 X.t5 24.923
R35 X.n4 X.t7 24.923
R36 X X.n2 8.457
R37 X X.n5 1.371
R38 VPWR.n0 VPWR.t6 580.224
R39 VPWR.n2 VPWR.n1 307.239
R40 VPWR.n8 VPWR.n7 307.239
R41 VPWR.n13 VPWR.n12 307.239
R42 VPWR.n18 VPWR.n17 307.239
R43 VPWR.n7 VPWR.t8 102.44
R44 VPWR.n17 VPWR.t7 63.321
R45 VPWR.n1 VPWR.t0 56.145
R46 VPWR.n17 VPWR.t2 55.113
R47 VPWR.n1 VPWR.t1 26.595
R48 VPWR.n7 VPWR.t5 26.595
R49 VPWR.n12 VPWR.t4 26.595
R50 VPWR.n12 VPWR.t3 26.595
R51 VPWR.n4 VPWR.n3 4.65
R52 VPWR.n6 VPWR.n5 4.65
R53 VPWR.n9 VPWR.n8 4.65
R54 VPWR.n11 VPWR.n10 4.65
R55 VPWR.n14 VPWR.n13 4.65
R56 VPWR.n16 VPWR.n15 4.65
R57 VPWR.n19 VPWR.n18 3.932
R58 VPWR.n3 VPWR.n2 1.882
R59 VPWR.n4 VPWR.n0 0.214
R60 VPWR.n19 VPWR.n16 0.137
R61 VPWR VPWR.n19 0.121
R62 VPWR.n6 VPWR.n4 0.119
R63 VPWR.n9 VPWR.n6 0.119
R64 VPWR.n11 VPWR.n9 0.119
R65 VPWR.n14 VPWR.n11 0.119
R66 VPWR.n16 VPWR.n14 0.119
R67 VPB.t5 VPB.t8 476.479
R68 VPB.t0 VPB.t6 349.221
R69 VPB.t1 VPB.t0 337.383
R70 VPB.t7 VPB.t2 281.152
R71 VPB.t8 VPB.t1 248.598
R72 VPB.t4 VPB.t5 248.598
R73 VPB.t3 VPB.t4 248.598
R74 VPB.t2 VPB.t3 248.598
R75 VPB VPB.t7 189.408
R76 B.n0 B.t1 241.534
R77 B.n0 B.t0 169.234
R78 B B.n0 78.133
R79 a_701_47.t0 a_701_47.t1 77.538
R80 a_815_47.t0 a_815_47.t1 81.23
R81 VNB VNB.t7 6438.23
R82 VNB.t1 VNB.t8 3892.31
R83 VNB.t6 VNB.t5 2852.75
R84 VNB.t0 VNB.t6 2756.04
R85 VNB.t7 VNB.t4 2255.35
R86 VNB.t8 VNB.t0 2030.77
R87 VNB.t3 VNB.t1 2030.77
R88 VNB.t2 VNB.t3 2030.77
R89 VNB.t4 VNB.t2 2030.77
R90 C.n0 C.t0 241.534
R91 C.n0 C.t1 169.234
R92 C C.n0 79.352
R93 a_27_47.n1 a_27_47.n0 469.411
R94 a_27_47.t0 a_27_47.n1 370.59
R95 a_27_47.n1 a_27_47.t1 240.658
R96 a_27_47.n0 a_27_47.t3 230.361
R97 a_27_47.n0 a_27_47.t2 158.061
R98 A_N.n0 A_N.t0 334.721
R99 A_N.n0 A_N.t1 206.188
R100 A_N.n1 A_N.n0 76
R101 A_N.n1 A_N 10.422
R102 A_N A_N.n1 2.011
R103 a_617_47.t0 a_617_47.t1 49.846
R104 D.n0 D.t0 241.534
R105 D.n0 D.t1 169.234
R106 D D.n0 79.2
R107 VGND.n3 VGND.n0 109.922
R108 VGND.n2 VGND.n1 107.433
R109 VGND.n7 VGND.n6 107.239
R110 VGND.n0 VGND.t1 89.538
R111 VGND.n6 VGND.t0 54.285
R112 VGND.n0 VGND.t2 31.384
R113 VGND.n6 VGND.t5 25.934
R114 VGND.n1 VGND.t4 24.923
R115 VGND.n1 VGND.t3 24.923
R116 VGND.n5 VGND.n4 4.65
R117 VGND.n8 VGND.n7 4.017
R118 VGND.n3 VGND.n2 3.878
R119 VGND.n5 VGND.n3 0.244
R120 VGND.n8 VGND.n5 0.135
R121 VGND VGND.n8 0.123
C0 VPB VPWR 0.10fF
C1 X VGND 0.25fF
C2 VPWR VGND 0.11fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__and4bb_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__and4bb_1 VGND VPWR A_N D X C B_N VNB VPB
X0 VPWR.t5 D.t0 a_343_93.t4 VPB.t5 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1 a_223_47.t0 B_N.t0 VGND.t0 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 a_515_93.t1 a_223_47.t2 a_429_93.t1 VNB.t5 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3 a_223_47.t1 B_N.t1 VPWR.t6 VPB.t6 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 VPWR.t4 A_N.t0 a_27_47.t1 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 VGND.t2 A_N.t1 a_27_47.t0 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 X.t1 a_343_93.t5 VPWR.t3 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 a_429_93.t0 a_27_47.t2 a_343_93.t1 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 VGND.t3 D.t1 a_615_93.t1 VNB.t6 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9 a_343_93.t0 C.t0 VPWR.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10 a_343_93.t2 a_27_47.t3 VPWR.t1 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11 a_615_93.t0 C.t1 a_515_93.t0 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12 X.t0 a_343_93.t6 VGND.t1 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 VPWR.t2 a_223_47.t3 a_343_93.t3 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
R0 D.n0 D.t0 334.721
R1 D.n0 D.t1 132.281
R2 D.n1 D.n0 76
R3 D.n1 D 16.158
R4 D D.n1 2.76
R5 a_343_93.n2 a_343_93.n1 308.688
R6 a_343_93.n4 a_343_93.n3 308.688
R7 a_343_93.n2 a_343_93.t1 224.845
R8 a_343_93.n0 a_343_93.t5 224.803
R9 a_343_93.n3 a_343_93.n0 189.694
R10 a_343_93.n0 a_343_93.t6 152.503
R11 a_343_93.n4 a_343_93.t4 93.809
R12 a_343_93.t0 a_343_93.n4 79.738
R13 a_343_93.n3 a_343_93.n2 71.905
R14 a_343_93.n1 a_343_93.t2 68.011
R15 a_343_93.n1 a_343_93.t3 63.321
R16 VPWR.n8 VPWR.t1 384.631
R17 VPWR.n1 VPWR.n0 310.819
R18 VPWR.n3 VPWR.n2 307.239
R19 VPWR.n14 VPWR.n13 307.239
R20 VPWR.n0 VPWR.t5 152.44
R21 VPWR.n2 VPWR.t0 89.119
R22 VPWR.n2 VPWR.t2 75.047
R23 VPWR.n13 VPWR.t6 68.011
R24 VPWR.n13 VPWR.t4 63.321
R25 VPWR.n0 VPWR.t3 27.955
R26 VPWR.n5 VPWR.n4 4.65
R27 VPWR.n7 VPWR.n6 4.65
R28 VPWR.n10 VPWR.n9 4.65
R29 VPWR.n12 VPWR.n11 4.65
R30 VPWR.n9 VPWR.n8 4.141
R31 VPWR.n15 VPWR.n14 4.115
R32 VPWR.n4 VPWR.n3 3.011
R33 VPWR.n5 VPWR.n1 0.197
R34 VPWR.n15 VPWR.n12 0.133
R35 VPWR VPWR.n15 0.128
R36 VPWR.n7 VPWR.n5 0.119
R37 VPWR.n10 VPWR.n7 0.119
R38 VPWR.n12 VPWR.n10 0.119
R39 VPB.t6 VPB.t1 609.657
R40 VPB.t5 VPB.t3 361.059
R41 VPB.t0 VPB.t5 307.788
R42 VPB.t2 VPB.t0 295.95
R43 VPB VPB.t4 275.233
R44 VPB.t1 VPB.t2 254.517
R45 VPB.t4 VPB.t6 254.517
R46 B_N.n0 B_N.t1 376.398
R47 B_N.n0 B_N.t0 164.318
R48 B_N B_N.n0 110.599
R49 VGND.n2 VGND.n0 114.084
R50 VGND.n2 VGND.n1 110.512
R51 VGND.n0 VGND.t3 94.285
R52 VGND.n1 VGND.t0 41.428
R53 VGND.n1 VGND.t2 38.571
R54 VGND.n0 VGND.t1 24
R55 VGND VGND.n2 0.157
R56 a_223_47.n1 a_223_47.t1 554.563
R57 a_223_47.n0 a_223_47.t3 334.721
R58 a_223_47.n1 a_223_47.n0 208.818
R59 a_223_47.t0 a_223_47.n1 151.071
R60 a_223_47.n0 a_223_47.t2 132.281
R61 VNB VNB.t4 7376.47
R62 VNB.t1 VNB.t2 6697.78
R63 VNB.t0 VNB.t6 3364.71
R64 VNB.t5 VNB.t0 3235.29
R65 VNB.t6 VNB.t3 3186.59
R66 VNB.t2 VNB.t5 2782.35
R67 VNB.t4 VNB.t1 2782.35
R68 a_429_93.t0 a_429_93.t1 80
R69 a_515_93.t0 a_515_93.t1 100
R70 A_N.n0 A_N.t1 392.464
R71 A_N.n0 A_N.t0 148.251
R72 A_N A_N.n0 77.645
R73 a_27_47.n1 a_27_47.t1 480.811
R74 a_27_47.t0 a_27_47.n1 231.899
R75 a_27_47.n1 a_27_47.n0 229.633
R76 a_27_47.n0 a_27_47.t2 188.113
R77 a_27_47.n0 a_27_47.t3 166.691
R78 X.n0 X.t1 172.965
R79 X X.t0 134.464
R80 X.n0 X 12.564
R81 X X.n0 4.065
R82 a_615_93.t0 a_615_93.t1 105.714
R83 C.n0 C.t0 334.721
R84 C.n0 C.t1 132.281
R85 C.n1 C.n0 76
R86 C.n1 C 17.484
R87 C C.n1 3.06
C0 C D 0.22fF
C1 A_N B_N 0.11fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__and4bb_2.ext - technology: sky130A

.subckt sky130_fd_sc_hd__and4bb_2 VGND VPWR A_N C B_N X D VNB VPB
X0 a_174_21.t0 C.t0 VPWR.t1 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1 a_174_21.t2 a_27_47.t2 VPWR.t4 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 a_476_47.t0 a_27_47.t3 a_174_21.t3 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3 VPWR.t5 a_174_21.t5 X.t3 VPB.t6 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 X.t2 a_174_21.t6 VPWR.t6 VPB.t5 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 a_548_47.t0 a_505_280.t2 a_476_47.t1 VNB.t6 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 VPWR.t3 A_N.t0 a_27_47.t0 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7 X.t1 a_174_21.t7 VGND.t3 VNB.t5 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 VPWR.t2 D.t0 a_174_21.t1 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9 VGND.t0 D.t1 a_639_47.t0 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10 VPWR.t7 a_505_280.t3 a_174_21.t4 VPB.t7 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11 a_505_280.t0 B_N.t0 VPWR.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12 VGND.t2 a_174_21.t8 X.t0 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 a_505_280.t1 B_N.t1 VGND.t4 VNB.t7 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14 a_639_47.t1 C.t1 a_548_47.t1 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15 VGND.t1 A_N.t1 a_27_47.t1 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
R0 C.n0 C.t0 405.415
R1 C.n0 C.t1 135.495
R2 C.n1 C.n0 76
R3 C.n1 C 8.452
R4 C C.n1 7.969
R5 VPWR.n3 VPWR.n2 310.803
R6 VPWR.n15 VPWR.n14 307.239
R7 VPWR.n1 VPWR.n0 306.805
R8 VPWR.n9 VPWR.n8 164.624
R9 VPWR.n2 VPWR.t2 143.059
R10 VPWR.n8 VPWR.t5 90.682
R11 VPWR.n0 VPWR.t1 68.011
R12 VPWR.n2 VPWR.t0 63.321
R13 VPWR.n0 VPWR.t7 63.321
R14 VPWR.n14 VPWR.t3 63.321
R15 VPWR.n14 VPWR.t6 55.113
R16 VPWR.n8 VPWR.t4 35.178
R17 VPWR.n10 VPWR.n9 4.951
R18 VPWR.n5 VPWR.n4 4.65
R19 VPWR.n7 VPWR.n6 4.65
R20 VPWR.n11 VPWR.n10 4.65
R21 VPWR.n13 VPWR.n12 4.65
R22 VPWR.n3 VPWR.n1 3.976
R23 VPWR.n16 VPWR.n15 3.932
R24 VPWR.n5 VPWR.n3 0.21
R25 VPWR.n16 VPWR.n13 0.137
R26 VPWR VPWR.n16 0.121
R27 VPWR.n7 VPWR.n5 0.119
R28 VPWR.n11 VPWR.n7 0.119
R29 VPWR.n13 VPWR.n11 0.119
R30 a_174_21.n5 a_174_21.n4 372.688
R31 a_174_21.n4 a_174_21.n0 308.688
R32 a_174_21.n2 a_174_21.t5 212.079
R33 a_174_21.n1 a_174_21.t6 212.079
R34 a_174_21.n3 a_174_21.n2 167.247
R35 a_174_21.n3 a_174_21.t3 147.259
R36 a_174_21.n2 a_174_21.t8 139.779
R37 a_174_21.n1 a_174_21.t7 139.779
R38 a_174_21.n4 a_174_21.n3 112.564
R39 a_174_21.n0 a_174_21.t2 86.773
R40 a_174_21.n0 a_174_21.t4 63.321
R41 a_174_21.n5 a_174_21.t1 63.321
R42 a_174_21.t0 a_174_21.n5 63.321
R43 a_174_21.n2 a_174_21.n1 61.345
R44 VPB.t6 VPB.t4 506.074
R45 VPB.t2 VPB.t0 349.221
R46 VPB.t3 VPB.t5 281.152
R47 VPB.t4 VPB.t7 278.193
R48 VPB.t7 VPB.t1 254.517
R49 VPB.t1 VPB.t2 248.598
R50 VPB.t5 VPB.t6 248.598
R51 VPB VPB.t3 189.408
R52 a_27_47.t0 a_27_47.n1 398.738
R53 a_27_47.n0 a_27_47.t2 326.76
R54 a_27_47.n1 a_27_47.t1 253.046
R55 a_27_47.n1 a_27_47.n0 219.47
R56 a_27_47.n0 a_27_47.t3 149.407
R57 a_476_47.t0 a_476_47.t1 60
R58 VNB VNB.t2 6438.23
R59 VNB.t4 VNB.t3 5321.88
R60 VNB.t0 VNB.t7 3817.65
R61 VNB.t6 VNB.t1 2944.12
R62 VNB.t1 VNB.t0 2717.65
R63 VNB.t3 VNB.t6 2329.41
R64 VNB.t2 VNB.t5 2255.35
R65 VNB.t5 VNB.t4 2030.77
R66 X X.n0 303.024
R67 X X.n1 112.126
R68 X.n0 X.t3 26.595
R69 X.n0 X.t2 26.595
R70 X.n1 X.t0 24.923
R71 X.n1 X.t1 24.923
R72 a_505_280.t0 a_505_280.n1 370.59
R73 a_505_280.n0 a_505_280.t2 336.328
R74 a_505_280.n1 a_505_280.t1 243.519
R75 a_505_280.n1 a_505_280.n0 209.646
R76 a_505_280.n0 a_505_280.t3 204.581
R77 a_548_47.t0 a_548_47.t1 87.142
R78 A_N.n0 A_N.t0 323.341
R79 A_N.n0 A_N.t1 194.808
R80 A_N.n1 A_N.n0 76
R81 A_N.n1 A_N 20.266
R82 A_N A_N.n1 3.911
R83 VGND.n1 VGND.t2 190.315
R84 VGND.n2 VGND.n0 118.086
R85 VGND.n6 VGND.n5 107.239
R86 VGND.n0 VGND.t0 87.142
R87 VGND.n5 VGND.t3 41.648
R88 VGND.n0 VGND.t4 38.571
R89 VGND.n5 VGND.t1 38.571
R90 VGND.n4 VGND.n3 4.65
R91 VGND.n2 VGND.n1 3.992
R92 VGND.n7 VGND.n6 3.932
R93 VGND.n4 VGND.n2 0.138
R94 VGND.n7 VGND.n4 0.137
R95 VGND VGND.n7 0.121
R96 D.n0 D.t0 309.015
R97 D.n0 D.t1 231.895
R98  D.n0 81.665
R99  D 14.268
R100 a_639_47.t0 a_639_47.t1 77.142
R101 B_N.n0 B_N.t0 408.628
R102 B_N.n0 B_N.t1 132.281
R103 B_N.n1 B_N.n0 76
R104  B_N.n1 6.4
R105 B_N.n1 B_N 6.034
C0 D B_N 0.14fF
C1 D C 0.21fF
C2 VGND VPWR 0.10fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__and4bb_4.ext - technology: sky130A

.subckt sky130_fd_sc_hd__and4bb_4 C A_N D X B_N VGND VPWR VNB VPB
X0 VPWR.t4 a_174_21.t5 X.t6 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_174_21.t2 a_832_21.t2 a_766_47.t1 VNB.t5 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 X.t5 a_174_21.t6 VPWR.t3 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 a_832_21.t0 A_N.t0 VGND.t0 VNB.t9 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 a_766_47.t0 a_27_47.t2 a_652_47.t0 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 VPWR.t2 a_174_21.t7 X.t4 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 X.t3 a_174_21.t8 VPWR.t1 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 VPWR.t8 B_N.t0 a_27_47.t0 VPB.t8 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 a_652_47.t1 C.t0 a_556_47.t0 VNB.t6 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 a_832_21.t1 A_N.t1 VPWR.t9 VPB.t9 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10 X.t2 a_174_21.t9 VGND.t4 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 X.t1 a_174_21.t10 VGND.t3 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 a_556_47.t1 D.t0 VGND.t5 VNB.t7 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 a_174_21.t4 D.t1 VPWR.t7 VPB.t7 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14 VPWR.t5 C.t1 a_174_21.t1 VPB.t5 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 VGND.t2 a_174_21.t11 X.t0 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X16 VGND.t1 a_174_21.t12 X.t7 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X17 VPWR.t6 a_832_21.t3 a_174_21.t3 VPB.t6 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X18 a_174_21.t0 a_27_47.t3 VPWR.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X19 VGND.t6 B_N.t1 a_27_47.t1 VNB.t8 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
R0 a_174_21.n11 a_174_21.n10 368.547
R1 a_174_21.n10 a_174_21.n0 292.5
R2 a_174_21.n9 a_174_21.t2 259.797
R3 a_174_21.n7 a_174_21.t5 196.012
R4 a_174_21.n1 a_174_21.t6 196.012
R5 a_174_21.n4 a_174_21.t7 196.012
R6 a_174_21.n3 a_174_21.t8 196.012
R7 a_174_21.n7 a_174_21.t12 149.419
R8 a_174_21.n1 a_174_21.t10 149.419
R9 a_174_21.n4 a_174_21.t11 149.419
R10 a_174_21.n3 a_174_21.t9 149.419
R11 a_174_21.n6 a_174_21.n5 101.6
R12 a_174_21.n8 a_174_21.n7 82.885
R13 a_174_21.n6 a_174_21.n2 76
R14 a_174_21.n10 a_174_21.n9 64.752
R15 a_174_21.n4 a_174_21.n3 57.84
R16 a_174_21.n0 a_174_21.t4 38.415
R17 a_174_21.n11 a_174_21.t3 34.475
R18 a_174_21.t0 a_174_21.n11 30.535
R19 a_174_21.n5 a_174_21.n4 28.92
R20 a_174_21.n0 a_174_21.t1 26.595
R21 a_174_21.n8 a_174_21.n6 25.6
R22 a_174_21.n2 a_174_21.n1 17.902
R23 a_174_21.n9 a_174_21.n8 12.047
R24 X.n2 X.n0 349.347
R25 X.n2 X.n1 292.5
R26 X.n5 X.n3 166.664
R27 X.n5 X.n4 113.702
R28 X.n0 X.t6 26.595
R29 X.n0 X.t5 26.595
R30 X.n1 X.t4 26.595
R31 X.n1 X.t3 26.595
R32 X.n3 X.t7 24.923
R33 X.n3 X.t1 24.923
R34 X.n4 X.t0 24.923
R35 X.n4 X.t2 24.923
R36 X X.n2 8.457
R37 X X.n5 1.371
R38 VPWR.n13 VPWR.n12 307.239
R39 VPWR.n18 VPWR.n17 307.239
R40 VPWR.n23 VPWR.n22 307.239
R41 VPWR.n28 VPWR.n27 307.239
R42 VPWR.n7 VPWR.n6 292.5
R43 VPWR.n3 VPWR.n2 292.5
R44 VPWR.n1 VPWR.n0 292.5
R45 VPWR.n0 VPWR.t9 107.88
R46 VPWR.n6 VPWR.t6 65.479
R47 VPWR.n27 VPWR.t8 63.321
R48 VPWR.n27 VPWR.t1 55.113
R49 VPWR.n12 VPWR.t5 46.295
R50 VPWR.n17 VPWR.t7 42.355
R51 VPWR.n12 VPWR.t0 36.445
R52 VPWR.n17 VPWR.t4 26.595
R53 VPWR.n22 VPWR.t3 26.595
R54 VPWR.n22 VPWR.t2 26.595
R55 VPWR.n5 VPWR.n1 6.205
R56 VPWR.n5 VPWR.n4 4.65
R57 VPWR.n9 VPWR.n8 4.65
R58 VPWR.n11 VPWR.n10 4.65
R59 VPWR.n14 VPWR.n13 4.65
R60 VPWR.n16 VPWR.n15 4.65
R61 VPWR.n19 VPWR.n18 4.65
R62 VPWR.n21 VPWR.n20 4.65
R63 VPWR.n24 VPWR.n23 4.65
R64 VPWR.n26 VPWR.n25 4.65
R65 VPWR.n29 VPWR.n28 3.932
R66 VPWR.n8 VPWR.n7 3.607
R67 VPWR.n4 VPWR.n3 0.814
R68 VPWR.n29 VPWR.n26 0.137
R69 VPWR VPWR.n29 0.121
R70 VPWR.n9 VPWR.n5 0.119
R71 VPWR.n11 VPWR.n9 0.119
R72 VPWR.n14 VPWR.n11 0.119
R73 VPWR.n16 VPWR.n14 0.119
R74 VPWR.n19 VPWR.n16 0.119
R75 VPWR.n21 VPWR.n19 0.119
R76 VPWR.n24 VPWR.n21 0.119
R77 VPWR.n26 VPWR.n24 0.119
R78 VPB.t6 VPB.t9 754.672
R79 VPB.t5 VPB.t0 337.383
R80 VPB.t4 VPB.t7 295.95
R81 VPB.t0 VPB.t6 284.112
R82 VPB.t7 VPB.t5 284.112
R83 VPB.t8 VPB.t1 281.152
R84 VPB.t3 VPB.t4 248.598
R85 VPB.t2 VPB.t3 248.598
R86 VPB.t1 VPB.t2 248.598
R87 VPB VPB.t8 189.408
R88 a_832_21.n1 a_832_21.t1 480.432
R89 a_832_21.t0 a_832_21.n1 225.564
R90 a_832_21.n0 a_832_21.t3 212.079
R91 a_832_21.n1 a_832_21.n0 192.848
R92 a_832_21.n0 a_832_21.t2 139.779
R93 a_766_47.t0 a_766_47.t1 60.923
R94 VNB.t5 VNB.t9 7489.53
R95 VNB VNB.t8 6438.23
R96 VNB.t6 VNB.t0 2756.04
R97 VNB.t1 VNB.t7 2417.58
R98 VNB.t0 VNB.t5 2320.88
R99 VNB.t7 VNB.t6 2320.88
R100 VNB.t8 VNB.t4 2255.35
R101 VNB.t3 VNB.t1 2030.77
R102 VNB.t2 VNB.t3 2030.77
R103 VNB.t4 VNB.t2 2030.77
R104 A_N.n0 A_N.t1 334.721
R105 A_N.n0 A_N.t0 206.188
R106 A_N.n1 A_N.n0 76
R107 A_N.n1 A_N 10.133
R108 A_N A_N.n1 1.955
R109 VGND.n2 VGND.t0 195.425
R110 VGND.n6 VGND.n5 107.433
R111 VGND.n11 VGND.n10 107.239
R112 VGND.n1 VGND.n0 106.463
R113 VGND.n10 VGND.t6 54.285
R114 VGND.n0 VGND.t5 36
R115 VGND.n0 VGND.t1 28.615
R116 VGND.n10 VGND.t4 25.934
R117 VGND.n5 VGND.t3 24.923
R118 VGND.n5 VGND.t2 24.923
R119 VGND.n4 VGND.n3 4.65
R120 VGND.n7 VGND.n6 4.65
R121 VGND.n9 VGND.n8 4.65
R122 VGND.n2 VGND.n1 4.069
R123 VGND.n12 VGND.n11 4.017
R124 VGND.n4 VGND.n2 0.136
R125 VGND.n12 VGND.n9 0.135
R126 VGND VGND.n12 0.123
R127 VGND.n7 VGND.n4 0.119
R128 VGND.n9 VGND.n7 0.119
R129 a_27_47.n1 a_27_47.n0 470.54
R130 a_27_47.t0 a_27_47.n1 370.59
R131 a_27_47.n0 a_27_47.t3 241.534
R132 a_27_47.n1 a_27_47.t1 240.658
R133 a_27_47.n0 a_27_47.t2 169.234
R134 a_652_47.t0 a_652_47.t1 77.538
R135 B_N.n0 B_N.t0 334.721
R136 B_N.n0 B_N.t1 206.188
R137 B_N.n1 B_N.n0 76
R138 B_N.n1 B_N 10.422
R139 B_N B_N.n1 2.011
R140 C.n0 C.t1 234.17
R141 C.n0 C.t0 161.87
R142 C C.n0 78.386
R143 a_556_47.t0 a_556_47.t1 60.923
R144 D.n0 D.t1 241.534
R145 D.n0 D.t0 169.234
R146 D D.n0 81.624
C0 X VGND 0.26fF
C1 X B_N 0.10fF
C2 VPWR VGND 0.14fF
C3 VPWR VPB 0.12fF
C4 C D 0.11fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__buf_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__buf_1 VGND VPWR X A VNB VPB
X0 VPWR.t1 A.t0 a_27_47.t1 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X1 X.t1 a_27_47.t2 VGND.t0 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X2 X.t0 a_27_47.t3 VPWR.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X3 VGND.t1 A.t1 a_27_47.t0 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
R0 A.n0 A.t0 260.32
R1 A.n0 A.t1 175.167
R2 A A.n0 80.324
R3 a_27_47.t1 a_27_47.n1 259.364
R4 a_27_47.n0 a_27_47.t3 254.387
R5 a_27_47.n0 a_27_47.t2 211.007
R6 a_27_47.n1 a_27_47.t0 202.108
R7 a_27_47.n1 a_27_47.n0 76
R8 VPWR VPWR.n0 178.435
R9 VPWR.n0 VPWR.t0 36.158
R10 VPWR.n0 VPWR.t1 36.158
R11 VPB.t1 VPB.t0 260.436
R12 VPB VPB.t1 192.367
R13 VGND VGND.n0 119.156
R14 VGND.n0 VGND.t0 33.461
R15 VGND.n0 VGND.t1 33.461
R16 X.n1 X.t0 222.242
R17 X.n0 X.t1 123.653
R18 X X.n0 78.877
R19 X.n1 X 10.483
R20 X X.n1 5.504
R21 X.n0 X 5.169
R22 VNB VNB.t1 6215.08
R23 VNB.t1 VNB.t0 2482.05
C0 VPWR X 0.13fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__buf_2.ext - technology: sky130A

.subckt sky130_fd_sc_hd__buf_2 VPWR VGND X A VNB VPB
X0 VPWR.t1 a_27_47.t2 X.t3 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 X.t2 a_27_47.t3 VPWR.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 VPWR.t2 A.t0 a_27_47.t0 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X3 X.t1 a_27_47.t4 VGND.t2 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 VGND.t1 a_27_47.t5 X.t0 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 VGND.t0 A.t1 a_27_47.t1 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
R0 a_27_47.t0 a_27_47.n2 301.066
R1 a_27_47.n0 a_27_47.t2 212.079
R2 a_27_47.n1 a_27_47.t3 212.079
R3 a_27_47.n2 a_27_47.t1 208.998
R4 a_27_47.n0 a_27_47.t5 139.779
R5 a_27_47.n1 a_27_47.t4 139.779
R6 a_27_47.n2 a_27_47.n1 84.033
R7 a_27_47.n1 a_27_47.n0 61.345
R8 X.n1 X.n0 143.643
R9 X.n3 X.n2 92.5
R10 X X.n3 81.316
R11 X.n0 X.t3 26.595
R12 X.n0 X.t2 26.595
R13 X.n2 X.t0 24.923
R14 X.n2 X.t1 24.923
R15 X X.n1 9.024
R16 X.n1 X 7.642
R17 X.n3 X 5.27
R18 VPWR.n1 VPWR.n0 168.558
R19 VPWR.n1 VPWR.t1 156.28
R20 VPWR.n0 VPWR.t2 55.406
R21 VPWR.n0 VPWR.t0 34.09
R22 VPWR VPWR.n1 10.029
R23 VPB.t2 VPB.t0 281.152
R24 VPB.t0 VPB.t1 248.598
R25 VPB VPB.t2 192.367
R26 A.n0 A.t0 276.463
R27 A.n0 A.t1 196.13
R28 A A.n0 80.324
R29 VGND.n1 VGND.t1 112.799
R30 VGND.n1 VGND.n0 110.032
R31 VGND.n0 VGND.t0 51.428
R32 VGND.n0 VGND.t2 28.791
R33 VGND VGND.n1 10.029
R34 VNB VNB.t0 6470.59
R35 VNB.t0 VNB.t2 2255.35
R36 VNB.t2 VNB.t1 2030.77
C0 VPWR X 0.26fF
C1 X VGND 0.16fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__buf_4.ext - technology: sky130A

.subckt sky130_fd_sc_hd__buf_4 VPWR VGND X A VNB VPB
X0 VPWR.t3 a_27_47.t2 X.t3 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 X.t2 a_27_47.t3 VPWR.t2 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 VPWR.t1 a_27_47.t4 X.t1 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 X.t0 a_27_47.t5 VPWR.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 X.t7 a_27_47.t6 VGND.t3 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 X.t6 a_27_47.t7 VGND.t2 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 VGND.t1 a_27_47.t8 X.t5 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 VGND.t0 a_27_47.t9 X.t4 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 VPWR.t4 A.t0 a_27_47.t0 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 VGND.t4 A.t1 a_27_47.t1 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
R0 a_27_47.n0 a_27_47.t2 221.719
R1 a_27_47.n1 a_27_47.t3 221.719
R2 a_27_47.n2 a_27_47.t4 221.719
R3 a_27_47.n3 a_27_47.t5 221.719
R4 a_27_47.n5 a_27_47.t1 178.41
R5 a_27_47.t0 a_27_47.n5 174.113
R6 a_27_47.n0 a_27_47.t9 149.419
R7 a_27_47.n1 a_27_47.t7 149.419
R8 a_27_47.n2 a_27_47.t8 149.419
R9 a_27_47.n3 a_27_47.t6 149.419
R10 a_27_47.n5 a_27_47.n4 94.823
R11 a_27_47.n1 a_27_47.n0 74.977
R12 a_27_47.n2 a_27_47.n1 74.977
R13 a_27_47.n4 a_27_47.n2 59.803
R14 a_27_47.n4 a_27_47.n3 15.174
R15 X.n3 X.n1 197.594
R16 X.n3 X.n2 167.415
R17 X.n4 X.n0 138.052
R18 X X.n5 106.451
R19 X.n1 X.t1 26.595
R20 X.n1 X.t0 26.595
R21 X.n2 X.t3 26.595
R22 X.n2 X.t2 26.595
R23 X.n0 X.t5 24.923
R24 X.n0 X.t7 24.923
R25 X.n5 X.t4 24.923
R26 X.n5 X.t6 24.923
R27 X.n4 X 7.369
R28 X X.n3 2.197
R29 X X.n4 1.422
R30 VPWR.n1 VPWR.n0 170.914
R31 VPWR.n3 VPWR.n2 164.214
R32 VPWR.n4 VPWR.t3 149.534
R33 VPWR.n0 VPWR.t0 26.595
R34 VPWR.n0 VPWR.t4 26.595
R35 VPWR.n2 VPWR.t2 26.595
R36 VPWR.n2 VPWR.t1 26.595
R37 VPWR VPWR.n7 9.575
R38 VPWR.n6 VPWR.n5 4.65
R39 VPWR.n4 VPWR.n3 3.9
R40 VPWR.n7 VPWR.n1 3.464
R41 VPWR.n7 VPWR.n6 0.72
R42 VPWR.n6 VPWR.n4 0.29
R43 VPB.t2 VPB.t3 248.598
R44 VPB.t1 VPB.t2 248.598
R45 VPB.t0 VPB.t1 248.598
R46 VPB.t4 VPB.t0 248.598
R47 VPB VPB.t4 189.408
R48 VGND.n1 VGND.n0 113.833
R49 VGND.n3 VGND.n2 108.015
R50 VGND.n4 VGND.t0 107.174
R51 VGND.n0 VGND.t3 24.923
R52 VGND.n0 VGND.t4 24.923
R53 VGND.n2 VGND.t2 24.923
R54 VGND.n2 VGND.t1 24.923
R55 VGND VGND.n7 9.372
R56 VGND.n6 VGND.n5 4.65
R57 VGND.n4 VGND.n3 3.9
R58 VGND.n7 VGND.n1 3.266
R59 VGND.n7 VGND.n6 0.821
R60 VGND.n6 VGND.n4 0.29
R61 VNB VNB.t4 6053.91
R62 VNB.t2 VNB.t0 2030.77
R63 VNB.t1 VNB.t2 2030.77
R64 VNB.t3 VNB.t1 2030.77
R65 VNB.t4 VNB.t3 2030.77
R66 A.n0 A.t0 235.762
R67 A.n0 A.t1 163.462
R68 A A.n0 84.266
C0 VPWR X 0.50fF
C1 X VGND 0.35fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__buf_6.ext - technology: sky130A

.subckt sky130_fd_sc_hd__buf_6 VPWR VGND X A VNB VPB
X0 VPWR.t5 a_161_47.t4 X.t11 VPB.t5 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_161_47.t0 A.t0 VGND.t7 VNB.t7 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 X.t10 a_161_47.t5 VPWR.t4 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 VPWR.t3 a_161_47.t6 X.t9 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 VGND.t6 A.t1 a_161_47.t1 VNB.t6 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 X.t8 a_161_47.t7 VPWR.t2 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 VGND.t5 a_161_47.t8 X.t5 VNB.t5 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 VGND.t4 a_161_47.t9 X.t4 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 VPWR.t1 a_161_47.t10 X.t7 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 X.t6 a_161_47.t11 VPWR.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 X.t3 a_161_47.t12 VGND.t3 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 X.t2 a_161_47.t13 VGND.t2 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 X.t1 a_161_47.t14 VGND.t1 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 VPWR.t6 A.t2 a_161_47.t2 VPB.t6 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14 VGND.t0 a_161_47.t15 X.t0 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X15 a_161_47.t3 A.t3 VPWR.t7 VPB.t7 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
R0 a_161_47.n1 a_161_47.t4 221.719
R1 a_161_47.n2 a_161_47.t5 221.719
R2 a_161_47.n3 a_161_47.t6 221.719
R3 a_161_47.n4 a_161_47.t7 221.719
R4 a_161_47.n5 a_161_47.t10 221.719
R5 a_161_47.n6 a_161_47.t11 221.719
R6 a_161_47.n9 a_161_47.n8 150.153
R7 a_161_47.n1 a_161_47.t15 149.419
R8 a_161_47.n2 a_161_47.t14 149.419
R9 a_161_47.n3 a_161_47.t9 149.419
R10 a_161_47.n4 a_161_47.t13 149.419
R11 a_161_47.n5 a_161_47.t8 149.419
R12 a_161_47.n6 a_161_47.t12 149.419
R13 a_161_47.n8 a_161_47.n7 92.564
R14 a_161_47.n8 a_161_47.n0 91.229
R15 a_161_47.n2 a_161_47.n1 74.977
R16 a_161_47.n3 a_161_47.n2 74.977
R17 a_161_47.n4 a_161_47.n3 74.977
R18 a_161_47.n5 a_161_47.n4 74.977
R19 a_161_47.n7 a_161_47.n5 58.911
R20 a_161_47.t2 a_161_47.n9 26.595
R21 a_161_47.n9 a_161_47.t3 26.595
R22 a_161_47.n0 a_161_47.t1 24.923
R23 a_161_47.n0 a_161_47.t0 24.923
R24 a_161_47.n7 a_161_47.n6 16.066
R25 X X.n0 197.594
R26 X.n6 X.n4 165.218
R27 X.n7 X.n2 165.218
R28 X X.n1 138.052
R29 X.n6 X.n5 105.676
R30 X.n7 X.n3 105.676
R31 X.n0 X.t7 26.595
R32 X.n0 X.t6 26.595
R33 X.n4 X.t11 26.595
R34 X.n4 X.t10 26.595
R35 X.n2 X.t9 26.595
R36 X.n2 X.t8 26.595
R37 X.n1 X.t5 24.923
R38 X.n1 X.t3 24.923
R39 X.n5 X.t0 24.923
R40 X.n5 X.t1 24.923
R41 X.n3 X.t4 24.923
R42 X.n3 X.t2 24.923
R43 X.n7 X.n6 12.218
R44 X X.n7 5.963
R45 VPWR.n10 VPWR.n9 170.914
R46 VPWR.n2 VPWR.n1 164.214
R47 VPWR.n7 VPWR.n6 164.214
R48 VPWR.n0 VPWR.t7 159.459
R49 VPWR.n3 VPWR.t5 149.804
R50 VPWR.n1 VPWR.t4 26.595
R51 VPWR.n1 VPWR.t3 26.595
R52 VPWR.n6 VPWR.t2 26.595
R53 VPWR.n6 VPWR.t1 26.595
R54 VPWR.n9 VPWR.t0 26.595
R55 VPWR.n9 VPWR.t6 26.595
R56 VPWR.n17 VPWR.n0 21.835
R57 VPWR.n11 VPWR.n10 7.152
R58 VPWR VPWR.n17 6.023
R59 VPWR.n17 VPWR.n16 4.769
R60 VPWR.n5 VPWR.n4 4.65
R61 VPWR.n8 VPWR.n7 4.65
R62 VPWR.n12 VPWR.n11 4.65
R63 VPWR.n14 VPWR.n13 4.65
R64 VPWR.n16 VPWR.n15 4.65
R65 VPWR.n3 VPWR.n2 3.704
R66 VPWR.n5 VPWR.n3 0.269
R67 VPWR.n8 VPWR.n5 0.119
R68 VPWR.n12 VPWR.n8 0.119
R69 VPWR.n14 VPWR.n12 0.119
R70 VPWR.n16 VPWR.n14 0.119
R71 VPB VPB.t7 343.302
R72 VPB.t4 VPB.t5 248.598
R73 VPB.t3 VPB.t4 248.598
R74 VPB.t2 VPB.t3 248.598
R75 VPB.t1 VPB.t2 248.598
R76 VPB.t0 VPB.t1 248.598
R77 VPB.t6 VPB.t0 248.598
R78 VPB.t7 VPB.t6 248.598
R79 A.n0 A.t2 221.719
R80 A.n2 A.t3 221.719
R81 A.n0 A.t1 149.419
R82 A.n2 A.t0 149.419
R83 A.n3 A.n2 109.025
R84 A.n1 A 82.933
R85 A.n2 A.n1 51.77
R86 A.n1 A.n0 23.207
R87 A.n3 A 18.4
R88 A A.n3 8.266
R89 VGND.n0 VGND.t7 190.063
R90 VGND.n12 VGND.n11 116.217
R91 VGND.n2 VGND.n1 108.015
R92 VGND.n7 VGND.n6 108.015
R93 VGND.n3 VGND.t0 107.444
R94 VGND.n1 VGND.t1 24.923
R95 VGND.n1 VGND.t4 24.923
R96 VGND.n6 VGND.t2 24.923
R97 VGND.n6 VGND.t5 24.923
R98 VGND.n11 VGND.t3 24.923
R99 VGND.n11 VGND.t6 24.923
R100 VGND.n17 VGND.n0 21.835
R101 VGND.n13 VGND.n12 15.811
R102 VGND VGND.n17 6.023
R103 VGND.n17 VGND.n16 4.769
R104 VGND.n5 VGND.n4 4.65
R105 VGND.n8 VGND.n7 4.65
R106 VGND.n10 VGND.n9 4.65
R107 VGND.n14 VGND.n13 4.65
R108 VGND.n16 VGND.n15 4.65
R109 VGND.n3 VGND.n2 3.704
R110 VGND.n5 VGND.n3 0.269
R111 VGND.n8 VGND.n5 0.119
R112 VGND.n10 VGND.n8 0.119
R113 VGND.n14 VGND.n10 0.119
R114 VGND.n16 VGND.n14 0.119
R115 VNB VNB.t7 8127.47
R116 VNB.t1 VNB.t0 2030.77
R117 VNB.t4 VNB.t1 2030.77
R118 VNB.t2 VNB.t4 2030.77
R119 VNB.t5 VNB.t2 2030.77
R120 VNB.t3 VNB.t5 2030.77
R121 VNB.t6 VNB.t3 2030.77
R122 VNB.t7 VNB.t6 2030.77
C0 VPWR X 0.76fF
C1 VGND X 0.56fF
C2 VGND VPWR 0.12fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__buf_8.ext - technology: sky130A

.subckt sky130_fd_sc_hd__buf_8 A X VGND VPWR VNB VPB
X0 X.t13 a_27_47.t6 VGND.t3 VNB.t10 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 X.t12 a_27_47.t7 VGND.t10 VNB.t9 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 X.t11 a_27_47.t8 VGND.t9 VNB.t8 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 VPWR.t10 a_27_47.t9 X.t5 VPB.t10 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 X.t4 a_27_47.t10 VPWR.t9 VPB.t9 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 VGND.t8 a_27_47.t11 X.t10 VNB.t7 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 VPWR.t0 A.t0 a_27_47.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 VPWR.t8 a_27_47.t12 X.t3 VPB.t8 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 a_27_47.t1 A.t1 VPWR.t1 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 X.t2 a_27_47.t13 VPWR.t7 VPB.t7 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 a_27_47.t2 A.t2 VGND.t0 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 X.t9 a_27_47.t14 VGND.t7 VNB.t6 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 VPWR.t6 a_27_47.t15 X.t1 VPB.t6 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13 X.t0 a_27_47.t16 VPWR.t5 VPB.t5 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14 VGND.t1 A.t3 a_27_47.t3 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X15 VGND.t6 a_27_47.t17 X.t8 VNB.t5 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X16 VPWR.t4 a_27_47.t18 X.t15 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17 VGND.t5 a_27_47.t19 X.t7 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X18 VGND.t4 a_27_47.t20 X.t6 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X19 X.t14 a_27_47.t21 VPWR.t3 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X20 VPWR.t2 A.t4 a_27_47.t4 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X21 VGND.t2 A.t5 a_27_47.t5 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
R0 a_27_47.n0 a_27_47.t12 221.719
R1 a_27_47.n1 a_27_47.t13 221.719
R2 a_27_47.n2 a_27_47.t15 221.719
R3 a_27_47.n6 a_27_47.t16 221.719
R4 a_27_47.n9 a_27_47.t18 221.719
R5 a_27_47.n12 a_27_47.t21 221.719
R6 a_27_47.n15 a_27_47.t9 221.719
R7 a_27_47.n18 a_27_47.t10 221.719
R8 a_27_47.n22 a_27_47.t5 193.846
R9 a_27_47.n24 a_27_47.t4 173.405
R10 a_27_47.n0 a_27_47.t11 149.419
R11 a_27_47.n1 a_27_47.t8 149.419
R12 a_27_47.n2 a_27_47.t20 149.419
R13 a_27_47.n6 a_27_47.t7 149.419
R14 a_27_47.n9 a_27_47.t19 149.419
R15 a_27_47.n12 a_27_47.t6 149.419
R16 a_27_47.n15 a_27_47.t17 149.419
R17 a_27_47.n18 a_27_47.t14 149.419
R18 a_27_47.n25 a_27_47.n24 108.41
R19 a_27_47.n22 a_27_47.n21 105.676
R20 a_27_47.n5 a_27_47.n3 101.6
R21 a_27_47.n5 a_27_47.n4 76
R22 a_27_47.n8 a_27_47.n7 76
R23 a_27_47.n11 a_27_47.n10 76
R24 a_27_47.n14 a_27_47.n13 76
R25 a_27_47.n17 a_27_47.n16 76
R26 a_27_47.n20 a_27_47.n19 76
R27 a_27_47.n1 a_27_47.n0 74.977
R28 a_27_47.n3 a_27_47.n1 66.051
R29 a_27_47.n23 a_27_47.n22 48.962
R30 a_27_47.n24 a_27_47.n23 38.732
R31 a_27_47.n7 a_27_47.n6 37.488
R32 a_27_47.t0 a_27_47.n25 26.595
R33 a_27_47.n25 a_27_47.t1 26.595
R34 a_27_47.n8 a_27_47.n5 25.6
R35 a_27_47.n11 a_27_47.n8 25.6
R36 a_27_47.n14 a_27_47.n11 25.6
R37 a_27_47.n17 a_27_47.n14 25.6
R38 a_27_47.n20 a_27_47.n17 25.6
R39 a_27_47.n21 a_27_47.t3 24.923
R40 a_27_47.n21 a_27_47.t2 24.923
R41 a_27_47.n10 a_27_47.n9 23.207
R42 a_27_47.n19 a_27_47.n18 19.637
R43 a_27_47.n23 a_27_47.n20 18.447
R44 a_27_47.n3 a_27_47.n2 8.925
R45 a_27_47.n13 a_27_47.n12 8.925
R46 a_27_47.n16 a_27_47.n15 5.355
R47 VGND.n1 VGND.n0 108.015
R48 VGND.n6 VGND.n5 108.015
R49 VGND.n10 VGND.n9 108.015
R50 VGND.n16 VGND.n15 108.015
R51 VGND.n21 VGND.n20 108.015
R52 VGND.n2 VGND.t8 106.996
R53 VGND.n0 VGND.t9 24.923
R54 VGND.n0 VGND.t4 24.923
R55 VGND.n5 VGND.t10 24.923
R56 VGND.n5 VGND.t5 24.923
R57 VGND.n9 VGND.t3 24.923
R58 VGND.n9 VGND.t6 24.923
R59 VGND.n15 VGND.t7 24.923
R60 VGND.n15 VGND.t1 24.923
R61 VGND.n20 VGND.t0 24.923
R62 VGND.n20 VGND.t2 24.923
R63 VGND.n4 VGND.n3 4.65
R64 VGND.n8 VGND.n7 4.65
R65 VGND.n12 VGND.n11 4.65
R66 VGND.n14 VGND.n13 4.65
R67 VGND.n17 VGND.n16 4.65
R68 VGND.n19 VGND.n18 4.65
R69 VGND.n22 VGND.n21 3.932
R70 VGND.n2 VGND.n1 3.488
R71 VGND.n7 VGND.n6 3.388
R72 VGND.n11 VGND.n10 0.376
R73 VGND.n4 VGND.n2 0.263
R74 VGND.n22 VGND.n19 0.137
R75 VGND VGND.n22 0.121
R76 VGND.n8 VGND.n4 0.119
R77 VGND.n12 VGND.n8 0.119
R78 VGND.n14 VGND.n12 0.119
R79 VGND.n17 VGND.n14 0.119
R80 VGND.n19 VGND.n17 0.119
R81 X.n8 X.n7 228.465
R82 X.n11 X.n10 169.484
R83 X.n3 X.n2 168.923
R84 X.n9 X.n5 165.218
R85 X.n8 X.n6 165.218
R86 X X.n13 107.181
R87 X.n3 X.n1 105.676
R88 X.n4 X.n0 105.676
R89 X.n4 X.n3 63.247
R90 X.n9 X.n8 63.247
R91 X.n12 X.n4 50.447
R92 X.n11 X.n9 50.447
R93 X.n5 X.t1 26.595
R94 X.n5 X.t0 26.595
R95 X.n6 X.t15 26.595
R96 X.n6 X.t14 26.595
R97 X.n7 X.t5 26.595
R98 X.n7 X.t4 26.595
R99 X.n10 X.t3 26.595
R100 X.n10 X.t2 26.595
R101 X.n2 X.t8 24.923
R102 X.n2 X.t9 24.923
R103 X.n1 X.t7 24.923
R104 X.n1 X.t13 24.923
R105 X.n0 X.t6 24.923
R106 X.n0 X.t12 24.923
R107 X.n13 X.t10 24.923
R108 X.n13 X.t11 24.923
R109 X.n12 X 14.305
R110 X X.n11 4.266
R111 X X.n12 2.76
R112 VNB VNB.t2 6053.91
R113 VNB.t8 VNB.t7 2030.77
R114 VNB.t3 VNB.t8 2030.77
R115 VNB.t9 VNB.t3 2030.77
R116 VNB.t4 VNB.t9 2030.77
R117 VNB.t10 VNB.t4 2030.77
R118 VNB.t5 VNB.t10 2030.77
R119 VNB.t6 VNB.t5 2030.77
R120 VNB.t1 VNB.t6 2030.77
R121 VNB.t0 VNB.t1 2030.77
R122 VNB.t2 VNB.t0 2030.77
R123 VPWR.n22 VPWR.n21 174.594
R124 VPWR.n16 VPWR.n15 174.594
R125 VPWR.n1 VPWR.n0 164.214
R126 VPWR.n6 VPWR.n5 164.214
R127 VPWR.n10 VPWR.n9 164.214
R128 VPWR.n2 VPWR.t8 149.356
R129 VPWR.n0 VPWR.t7 26.595
R130 VPWR.n0 VPWR.t6 26.595
R131 VPWR.n5 VPWR.t5 26.595
R132 VPWR.n5 VPWR.t4 26.595
R133 VPWR.n9 VPWR.t3 26.595
R134 VPWR.n9 VPWR.t10 26.595
R135 VPWR.n21 VPWR.t1 26.595
R136 VPWR.n21 VPWR.t2 26.595
R137 VPWR.n15 VPWR.t9 26.595
R138 VPWR.n15 VPWR.t0 26.595
R139 VPWR.n17 VPWR.n16 6.776
R140 VPWR.n24 VPWR.n23 4.65
R141 VPWR.n4 VPWR.n3 4.65
R142 VPWR.n8 VPWR.n7 4.65
R143 VPWR.n12 VPWR.n11 4.65
R144 VPWR.n14 VPWR.n13 4.65
R145 VPWR.n18 VPWR.n17 4.65
R146 VPWR.n20 VPWR.n19 4.65
R147 VPWR.n2 VPWR.n1 3.488
R148 VPWR.n7 VPWR.n6 3.388
R149 VPWR.n23 VPWR.n22 0.752
R150 VPWR.n11 VPWR.n10 0.376
R151 VPWR.n4 VPWR.n2 0.263
R152 VPWR.n8 VPWR.n4 0.119
R153 VPWR.n12 VPWR.n8 0.119
R154 VPWR.n14 VPWR.n12 0.119
R155 VPWR.n18 VPWR.n14 0.119
R156 VPWR.n20 VPWR.n18 0.119
R157 VPWR.n24 VPWR.n20 0.119
R158 VPWR.n25 VPWR.n24 0.119
R159 VPWR VPWR.n25 0.02
R160 VPB.t7 VPB.t8 248.598
R161 VPB.t6 VPB.t7 248.598
R162 VPB.t5 VPB.t6 248.598
R163 VPB.t4 VPB.t5 248.598
R164 VPB.t3 VPB.t4 248.598
R165 VPB.t10 VPB.t3 248.598
R166 VPB.t9 VPB.t10 248.598
R167 VPB.t0 VPB.t9 248.598
R168 VPB.t1 VPB.t0 248.598
R169 VPB.t2 VPB.t1 248.598
R170 VPB VPB.t2 189.408
R171 A.n6 A.t4 235.762
R172 A.n0 A.t0 221.719
R173 A.n2 A.t1 221.719
R174 A.n6 A.t5 163.462
R175 A.n0 A.t3 149.419
R176 A.n2 A.t2 149.419
R177 A.n5 A.n4 76
R178 A.n7 A.n6 76
R179 A.n1 A.n0 58.018
R180 A.n5 A.n2 43.737
R181 A.n4 A.n3 21.76
R182 A.n7 A 19.52
R183 A.n6 A.n5 17.851
R184 A.n2 A.n1 16.959
R185 A A.n7 9.92
R186 A.n3 A 5.44
R187 A.n4 A 2.24
C0 VPB VPWR 0.12fF
C1 VGND X 0.80fF
C2 VGND VPWR 0.15fF
C3 VPWR X 1.02fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__buf_12.ext - technology: sky130A

.subckt sky130_fd_sc_hd__buf_12 A X VGND VPWR VNB VPB
X0 VGND.t11 a_109_47.t8 X.t10 VNB.t11 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 X.t0 a_109_47.t9 VPWR.t11 VPB.t11 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 VGND.t10 a_109_47.t10 X.t9 VNB.t10 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 VGND.t9 a_109_47.t11 X.t8 VNB.t9 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 VGND.t8 a_109_47.t12 X.t7 VNB.t8 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 X.t23 a_109_47.t13 VPWR.t10 VPB.t10 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 VPWR.t12 A.t0 a_109_47.t0 VPB.t12 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 X.t6 a_109_47.t14 VGND.t7 VNB.t7 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 X.t5 a_109_47.t15 VGND.t6 VNB.t6 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 X.t4 a_109_47.t16 VGND.t5 VNB.t5 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 a_109_47.t1 A.t1 VPWR.t13 VPB.t13 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 VPWR.t9 a_109_47.t17 X.t22 VPB.t9 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 X.t21 a_109_47.t18 VPWR.t8 VPB.t8 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13 VPWR.t14 A.t2 a_109_47.t2 VPB.t14 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14 VPWR.t7 a_109_47.t19 X.t20 VPB.t7 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 VGND.t12 A.t3 a_109_47.t3 VNB.t12 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X16 VGND.t13 A.t4 a_109_47.t4 VNB.t13 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X17 VGND.t4 a_109_47.t20 X.t3 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X18 X.t19 a_109_47.t21 VPWR.t6 VPB.t6 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X19 VPWR.t5 a_109_47.t22 X.t18 VPB.t5 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X20 a_109_47.t5 A.t5 VGND.t14 VNB.t14 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X21 X.t2 a_109_47.t23 VGND.t3 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X22 X.t17 a_109_47.t24 VPWR.t4 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X23 VPWR.t3 a_109_47.t25 X.t16 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X24 X.t1 a_109_47.t26 VGND.t2 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X25 X.t12 a_109_47.t27 VGND.t1 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X26 VPWR.t2 a_109_47.t28 X.t15 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X27 X.t14 a_109_47.t29 VPWR.t1 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X28 a_109_47.t6 A.t6 VPWR.t15 VPB.t15 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X29 VPWR.t0 a_109_47.t30 X.t13 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X30 a_109_47.t7 A.t7 VGND.t15 VNB.t15 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X31 VGND.t0 a_109_47.t31 X.t11 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
R0 a_109_47.n1 a_109_47.t25 221.719
R1 a_109_47.n2 a_109_47.t29 221.719
R2 a_109_47.n3 a_109_47.t30 221.719
R3 a_109_47.n4 a_109_47.t9 221.719
R4 a_109_47.n5 a_109_47.t17 221.719
R5 a_109_47.n6 a_109_47.t18 221.719
R6 a_109_47.n7 a_109_47.t19 221.719
R7 a_109_47.n11 a_109_47.t21 221.719
R8 a_109_47.n14 a_109_47.t22 221.719
R9 a_109_47.n17 a_109_47.t24 221.719
R10 a_109_47.n20 a_109_47.t28 221.719
R11 a_109_47.n23 a_109_47.t13 221.719
R12 a_109_47.n28 a_109_47.n27 168.923
R13 a_109_47.n1 a_109_47.t20 149.419
R14 a_109_47.n2 a_109_47.t15 149.419
R15 a_109_47.n3 a_109_47.t11 149.419
R16 a_109_47.n4 a_109_47.t14 149.419
R17 a_109_47.n5 a_109_47.t31 149.419
R18 a_109_47.n6 a_109_47.t16 149.419
R19 a_109_47.n7 a_109_47.t12 149.419
R20 a_109_47.n11 a_109_47.t27 149.419
R21 a_109_47.n14 a_109_47.t10 149.419
R22 a_109_47.n17 a_109_47.t26 149.419
R23 a_109_47.n20 a_109_47.t8 149.419
R24 a_109_47.n23 a_109_47.t23 149.419
R25 a_109_47.n30 a_109_47.n0 146.81
R26 a_109_47.n31 a_109_47.n30 108.41
R27 a_109_47.n28 a_109_47.n26 105.676
R28 a_109_47.n10 a_109_47.n8 101.6
R29 a_109_47.n10 a_109_47.n9 76
R30 a_109_47.n13 a_109_47.n12 76
R31 a_109_47.n16 a_109_47.n15 76
R32 a_109_47.n19 a_109_47.n18 76
R33 a_109_47.n22 a_109_47.n21 76
R34 a_109_47.n25 a_109_47.n24 76
R35 a_109_47.n2 a_109_47.n1 74.977
R36 a_109_47.n3 a_109_47.n2 74.977
R37 a_109_47.n4 a_109_47.n3 74.977
R38 a_109_47.n5 a_109_47.n4 74.977
R39 a_109_47.n6 a_109_47.n5 74.977
R40 a_109_47.n8 a_109_47.n6 66.051
R41 a_109_47.n29 a_109_47.n28 48.962
R42 a_109_47.n30 a_109_47.n29 38.732
R43 a_109_47.n12 a_109_47.n11 37.488
R44 a_109_47.n0 a_109_47.t2 26.595
R45 a_109_47.n0 a_109_47.t6 26.595
R46 a_109_47.t0 a_109_47.n31 26.595
R47 a_109_47.n31 a_109_47.t1 26.595
R48 a_109_47.n13 a_109_47.n10 25.6
R49 a_109_47.n16 a_109_47.n13 25.6
R50 a_109_47.n19 a_109_47.n16 25.6
R51 a_109_47.n22 a_109_47.n19 25.6
R52 a_109_47.n25 a_109_47.n22 25.6
R53 a_109_47.n27 a_109_47.t3 24.923
R54 a_109_47.n27 a_109_47.t7 24.923
R55 a_109_47.n26 a_109_47.t4 24.923
R56 a_109_47.n26 a_109_47.t5 24.923
R57 a_109_47.n15 a_109_47.n14 23.207
R58 a_109_47.n24 a_109_47.n23 19.637
R59 a_109_47.n29 a_109_47.n25 18.447
R60 a_109_47.n8 a_109_47.n7 8.925
R61 a_109_47.n18 a_109_47.n17 8.925
R62 a_109_47.n21 a_109_47.n20 5.355
R63 X.n3 X.n2 228.465
R64 X.n8 X.n7 168.923
R65 X.n4 X.n0 165.218
R66 X.n3 X.n1 165.218
R67 X.n16 X.n14 165.218
R68 X.n17 X.n12 165.218
R69 X.n18 X.n10 165.218
R70 X.n8 X.n6 105.676
R71 X.n9 X.n5 105.676
R72 X.n16 X.n15 105.676
R73 X.n17 X.n13 105.676
R74 X.n18 X.n11 105.676
R75 X.n4 X.n3 63.247
R76 X.n9 X.n8 63.247
R77 X X.n4 50.447
R78 X X.n9 50.447
R79 X.n0 X.t20 26.595
R80 X.n0 X.t19 26.595
R81 X.n1 X.t18 26.595
R82 X.n1 X.t17 26.595
R83 X.n2 X.t15 26.595
R84 X.n2 X.t23 26.595
R85 X.n14 X.t16 26.595
R86 X.n14 X.t14 26.595
R87 X.n12 X.t13 26.595
R88 X.n12 X.t0 26.595
R89 X.n10 X.t22 26.595
R90 X.n10 X.t21 26.595
R91 X.n7 X.t10 24.923
R92 X.n7 X.t2 24.923
R93 X.n6 X.t9 24.923
R94 X.n6 X.t1 24.923
R95 X.n5 X.t7 24.923
R96 X.n5 X.t12 24.923
R97 X.n15 X.t3 24.923
R98 X.n15 X.t5 24.923
R99 X.n13 X.t8 24.923
R100 X.n13 X.t6 24.923
R101 X.n11 X.t11 24.923
R102 X.n11 X.t4 24.923
R103 X.n17 X.n16 12.218
R104 X.n18 X.n17 12.218
R105 X X.n18 2.472
R106 VGND.n35 VGND.t15 181.861
R107 VGND.n1 VGND.n0 108.015
R108 VGND.n6 VGND.n5 108.015
R109 VGND.n11 VGND.n10 108.015
R110 VGND.n16 VGND.n15 108.015
R111 VGND.n20 VGND.n19 108.015
R112 VGND.n26 VGND.n25 108.015
R113 VGND.n31 VGND.n30 108.015
R114 VGND.n2 VGND.t4 94.664
R115 VGND.n0 VGND.t6 24.923
R116 VGND.n0 VGND.t9 24.923
R117 VGND.n5 VGND.t7 24.923
R118 VGND.n5 VGND.t0 24.923
R119 VGND.n10 VGND.t5 24.923
R120 VGND.n10 VGND.t8 24.923
R121 VGND.n15 VGND.t1 24.923
R122 VGND.n15 VGND.t10 24.923
R123 VGND.n19 VGND.t2 24.923
R124 VGND.n19 VGND.t11 24.923
R125 VGND.n25 VGND.t3 24.923
R126 VGND.n25 VGND.t13 24.923
R127 VGND.n30 VGND.t14 24.923
R128 VGND.n30 VGND.t12 24.923
R129 VGND VGND.n35 4.738
R130 VGND.n4 VGND.n3 4.65
R131 VGND.n7 VGND.n6 4.65
R132 VGND.n9 VGND.n8 4.65
R133 VGND.n12 VGND.n11 4.65
R134 VGND.n14 VGND.n13 4.65
R135 VGND.n18 VGND.n17 4.65
R136 VGND.n22 VGND.n21 4.65
R137 VGND.n24 VGND.n23 4.65
R138 VGND.n27 VGND.n26 4.65
R139 VGND.n29 VGND.n28 4.65
R140 VGND.n32 VGND.n31 4.65
R141 VGND.n34 VGND.n33 4.65
R142 VGND.n2 VGND.n1 3.89
R143 VGND.n21 VGND.n20 3.388
R144 VGND.n17 VGND.n16 0.376
R145 VGND.n4 VGND.n2 0.277
R146 VGND.n7 VGND.n4 0.119
R147 VGND.n9 VGND.n7 0.119
R148 VGND.n12 VGND.n9 0.119
R149 VGND.n14 VGND.n12 0.119
R150 VGND.n18 VGND.n14 0.119
R151 VGND.n22 VGND.n18 0.119
R152 VGND.n24 VGND.n22 0.119
R153 VGND.n27 VGND.n24 0.119
R154 VGND.n29 VGND.n27 0.119
R155 VGND.n32 VGND.n29 0.119
R156 VGND.n34 VGND.n32 0.119
R157 VGND VGND.n34 0.031
R158 VNB VNB.n0 4917.65
R159 VNB.t6 VNB.t4 2030.77
R160 VNB.t9 VNB.t6 2030.77
R161 VNB.t7 VNB.t9 2030.77
R162 VNB.t0 VNB.t7 2030.77
R163 VNB.t5 VNB.t0 2030.77
R164 VNB.t8 VNB.t5 2030.77
R165 VNB.t1 VNB.t8 2030.77
R166 VNB.t10 VNB.t1 2030.77
R167 VNB.t2 VNB.t10 2030.77
R168 VNB.t11 VNB.t2 2030.77
R169 VNB.t3 VNB.t11 2030.77
R170 VNB.t13 VNB.t3 2030.77
R171 VNB.t14 VNB.t13 2030.77
R172 VNB.t12 VNB.t14 2030.77
R173 VNB.n0 VNB.t12 1136.26
R174 VNB.n0 VNB.t15 894.505
R175 VPWR.n37 VPWR.t15 201.189
R176 VPWR.n32 VPWR.n31 174.594
R177 VPWR.n26 VPWR.n25 174.594
R178 VPWR.n20 VPWR.n19 164.214
R179 VPWR.n16 VPWR.n15 164.214
R180 VPWR.n11 VPWR.n10 164.214
R181 VPWR.n6 VPWR.n5 164.214
R182 VPWR.n1 VPWR.n0 164.214
R183 VPWR.n2 VPWR.t3 149.44
R184 VPWR.n31 VPWR.t13 26.595
R185 VPWR.n31 VPWR.t14 26.595
R186 VPWR.n25 VPWR.t10 26.595
R187 VPWR.n25 VPWR.t12 26.595
R188 VPWR.n19 VPWR.t4 26.595
R189 VPWR.n19 VPWR.t2 26.595
R190 VPWR.n15 VPWR.t6 26.595
R191 VPWR.n15 VPWR.t5 26.595
R192 VPWR.n10 VPWR.t8 26.595
R193 VPWR.n10 VPWR.t7 26.595
R194 VPWR.n5 VPWR.t11 26.595
R195 VPWR.n5 VPWR.t9 26.595
R196 VPWR.n0 VPWR.t1 26.595
R197 VPWR.n0 VPWR.t0 26.595
R198 VPWR.n27 VPWR.n26 9.788
R199 VPWR VPWR.n37 6.996
R200 VPWR.n4 VPWR.n3 4.65
R201 VPWR.n7 VPWR.n6 4.65
R202 VPWR.n9 VPWR.n8 4.65
R203 VPWR.n12 VPWR.n11 4.65
R204 VPWR.n14 VPWR.n13 4.65
R205 VPWR.n18 VPWR.n17 4.65
R206 VPWR.n22 VPWR.n21 4.65
R207 VPWR.n24 VPWR.n23 4.65
R208 VPWR.n28 VPWR.n27 4.65
R209 VPWR.n30 VPWR.n29 4.65
R210 VPWR.n34 VPWR.n33 4.65
R211 VPWR.n36 VPWR.n35 4.65
R212 VPWR.n2 VPWR.n1 3.89
R213 VPWR.n33 VPWR.n32 3.764
R214 VPWR.n21 VPWR.n20 3.388
R215 VPWR.n17 VPWR.n16 0.376
R216 VPWR.n4 VPWR.n2 0.277
R217 VPWR.n7 VPWR.n4 0.119
R218 VPWR.n9 VPWR.n7 0.119
R219 VPWR.n12 VPWR.n9 0.119
R220 VPWR.n14 VPWR.n12 0.119
R221 VPWR.n18 VPWR.n14 0.119
R222 VPWR.n22 VPWR.n18 0.119
R223 VPWR.n24 VPWR.n22 0.119
R224 VPWR.n28 VPWR.n24 0.119
R225 VPWR.n30 VPWR.n28 0.119
R226 VPWR.n34 VPWR.n30 0.119
R227 VPWR.n36 VPWR.n34 0.119
R228 VPWR VPWR.n36 0.031
R229 VPB.t1 VPB.t3 248.598
R230 VPB.t0 VPB.t1 248.598
R231 VPB.t11 VPB.t0 248.598
R232 VPB.t9 VPB.t11 248.598
R233 VPB.t8 VPB.t9 248.598
R234 VPB.t7 VPB.t8 248.598
R235 VPB.t6 VPB.t7 248.598
R236 VPB.t5 VPB.t6 248.598
R237 VPB.t4 VPB.t5 248.598
R238 VPB.t2 VPB.t4 248.598
R239 VPB.t10 VPB.t2 248.598
R240 VPB.t12 VPB.t10 248.598
R241 VPB.t13 VPB.t12 248.598
R242 VPB.t14 VPB.t13 248.598
R243 VPB VPB.t14 189.408
R244 VPB VPB.t15 59.19
R245 A.n9 A.t6 235.552
R246 A.n2 A.t0 221.719
R247 A.n4 A.t1 221.719
R248 A.n0 A.t2 221.719
R249 A.n9 A.t7 163.252
R250 A.n2 A.t4 149.419
R251 A.n4 A.t5 149.419
R252 A.n0 A.t3 149.419
R253 A.n6 A.n5 76
R254 A.n8 A.n7 76
R255 A.n10 A.n9 76
R256 A.n3 A.n2 58.018
R257 A.n5 A.n4 43.737
R258 A.n9 A.n8 32.133
R259 A.n5 A.n0 31.24
R260 A.n8 A.n0 29.455
R261 A.n6 A.n1 21.76
R262 A.n7 A 19.52
R263 A.n4 A.n3 16.959
R264 A.n10 A 11.84
R265 A.n7 A 9.92
R266 A A.n10 9.92
R267 A.n1 A 5.44
R268 A A.n6 2.24
C0 VPWR VGND 0.19fF
C1 VPWR X 1.56fF
C2 VPWR VPB 0.15fF
C3 X VGND 1.23fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__buf_16.ext - technology: sky130A

.subckt sky130_fd_sc_hd__buf_16 A X VGND VPWR VNB VPB
X0 VGND.t21 A.t0 a_109_47.t11 VNB.t21 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 X.t15 a_109_47.t12 VPWR.t15 VPB.t15 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 VGND.t3 a_109_47.t13 X.t31 VNB.t15 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 VGND.t2 a_109_47.t14 X.t30 VNB.t14 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 X.t14 a_109_47.t15 VPWR.t14 VPB.t14 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 VGND.t1 a_109_47.t16 X.t29 VNB.t13 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 VPWR.t13 a_109_47.t17 X.t13 VPB.t13 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 a_109_47.t6 A.t1 VPWR.t21 VPB.t21 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 X.t12 a_109_47.t18 VPWR.t12 VPB.t12 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 VPWR.t20 A.t2 a_109_47.t5 VPB.t20 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 X.t28 a_109_47.t19 VGND.t0 VNB.t12 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 X.t27 a_109_47.t20 VGND.t15 VNB.t11 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 X.t26 a_109_47.t21 VGND.t14 VNB.t10 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 X.t25 a_109_47.t22 VGND.t13 VNB.t9 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14 a_109_47.t4 A.t3 VPWR.t19 VPB.t19 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 VPWR.t11 a_109_47.t23 X.t11 VPB.t11 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16 X.t24 a_109_47.t24 VGND.t12 VNB.t8 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X17 X.t10 a_109_47.t25 VPWR.t10 VPB.t10 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X18 VPWR.t18 A.t4 a_109_47.t3 VPB.t18 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X19 VPWR.t9 a_109_47.t26 X.t9 VPB.t9 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X20 VGND.t20 A.t5 a_109_47.t10 VNB.t20 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X21 VGND.t19 A.t6 a_109_47.t9 VNB.t19 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X22 VGND.t11 a_109_47.t27 X.t23 VNB.t7 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X23 X.t8 a_109_47.t28 VPWR.t8 VPB.t8 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X24 VGND.t10 a_109_47.t29 X.t22 VNB.t6 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X25 VPWR.t7 a_109_47.t30 X.t7 VPB.t7 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X26 VGND.t9 a_109_47.t31 X.t21 VNB.t5 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X27 VPWR.t6 a_109_47.t32 X.t6 VPB.t6 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X28 X.t5 a_109_47.t33 VPWR.t5 VPB.t5 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X29 VGND.t8 a_109_47.t34 X.t20 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X30 a_109_47.t2 A.t7 VGND.t18 VNB.t18 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X31 a_109_47.t1 A.t8 VGND.t17 VNB.t17 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X32 X.t4 a_109_47.t35 VPWR.t4 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X33 VPWR.t3 a_109_47.t36 X.t3 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X34 X.t19 a_109_47.t37 VGND.t7 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X35 X.t18 a_109_47.t38 VGND.t6 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X36 VPWR.t17 A.t9 a_109_47.t8 VPB.t17 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X37 X.t2 a_109_47.t39 VPWR.t2 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X38 X.t17 a_109_47.t40 VGND.t5 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X39 a_109_47.t7 A.t10 VPWR.t16 VPB.t16 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X40 VPWR.t1 a_109_47.t41 X.t1 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X41 VPWR.t0 a_109_47.t42 X.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X42 a_109_47.t0 A.t11 VGND.t16 VNB.t16 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X43 VGND.t4 a_109_47.t43 X.t16 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
R0 A.n0 A.t9 221.719
R1 A.n2 A.t1 221.719
R2 A.n5 A.t2 221.719
R3 A.n13 A.t3 221.719
R4 A.n10 A.t4 221.719
R5 A.n8 A.t10 221.719
R6 A.n0 A.t0 149.419
R7 A.n2 A.t8 149.419
R8 A.n5 A.t6 149.419
R9 A.n13 A.t7 149.419
R10 A.n10 A.t5 149.419
R11 A.n8 A.t11 149.419
R12 A.n12 A.n9 97.76
R13 A.n1 A 95.84
R14 A.n4 A.n3 76
R15 A.n7 A.n6 76
R16 A.n15 A.n14 76
R17 A.n12 A.n11 76
R18 A.n1 A.n0 48.2
R19 A.n3 A.n2 33.918
R20 A.n2 A.n1 26.777
R21 A.n9 A.n8 23.207
R22 A.n7 A.n4 21.76
R23 A.n15 A.n12 21.76
R24 A.n6 A.n5 19.637
R25 A A.n15 16
R26 A.n11 A.n10 8.925
R27 A A.n7 5.76
R28 A.n14 A.n13 5.355
R29 A.n4 A 1.92
R30 a_109_47.n5 a_109_47.t42 221.719
R31 a_109_47.n6 a_109_47.t15 221.719
R32 a_109_47.n8 a_109_47.t17 221.719
R33 a_109_47.n13 a_109_47.t18 221.719
R34 a_109_47.n16 a_109_47.t30 221.719
R35 a_109_47.n19 a_109_47.t33 221.719
R36 a_109_47.n22 a_109_47.t36 221.719
R37 a_109_47.n27 a_109_47.t39 221.719
R38 a_109_47.n30 a_109_47.t41 221.719
R39 a_109_47.n33 a_109_47.t12 221.719
R40 a_109_47.n36 a_109_47.t23 221.719
R41 a_109_47.n41 a_109_47.t25 221.719
R42 a_109_47.n44 a_109_47.t26 221.719
R43 a_109_47.n47 a_109_47.t28 221.719
R44 a_109_47.n50 a_109_47.t32 221.719
R45 a_109_47.n53 a_109_47.t35 221.719
R46 a_109_47.n5 a_109_47.t34 149.419
R47 a_109_47.n6 a_109_47.t40 149.419
R48 a_109_47.n8 a_109_47.t31 149.419
R49 a_109_47.n13 a_109_47.t24 149.419
R50 a_109_47.n16 a_109_47.t29 149.419
R51 a_109_47.n19 a_109_47.t22 149.419
R52 a_109_47.n22 a_109_47.t27 149.419
R53 a_109_47.n27 a_109_47.t20 149.419
R54 a_109_47.n30 a_109_47.t14 149.419
R55 a_109_47.n33 a_109_47.t19 149.419
R56 a_109_47.n36 a_109_47.t43 149.419
R57 a_109_47.n41 a_109_47.t21 149.419
R58 a_109_47.n44 a_109_47.t16 149.419
R59 a_109_47.n47 a_109_47.t38 149.419
R60 a_109_47.n50 a_109_47.t13 149.419
R61 a_109_47.n53 a_109_47.t37 149.419
R62 a_109_47.n61 a_109_47.n60 146.811
R63 a_109_47.n58 a_109_47.n57 108.41
R64 a_109_47.n60 a_109_47.n59 108.41
R65 a_109_47.n2 a_109_47.n0 90.831
R66 a_109_47.n55 a_109_47.n54 76
R67 a_109_47.n10 a_109_47.n9 76
R68 a_109_47.n12 a_109_47.n11 76
R69 a_109_47.n15 a_109_47.n14 76
R70 a_109_47.n18 a_109_47.n17 76
R71 a_109_47.n21 a_109_47.n20 76
R72 a_109_47.n24 a_109_47.n23 76
R73 a_109_47.n26 a_109_47.n25 76
R74 a_109_47.n29 a_109_47.n28 76
R75 a_109_47.n32 a_109_47.n31 76
R76 a_109_47.n35 a_109_47.n34 76
R77 a_109_47.n38 a_109_47.n37 76
R78 a_109_47.n40 a_109_47.n39 76
R79 a_109_47.n43 a_109_47.n42 76
R80 a_109_47.n46 a_109_47.n45 76
R81 a_109_47.n49 a_109_47.n48 76
R82 a_109_47.n52 a_109_47.n51 76
R83 a_109_47.n10 a_109_47.n7 53.45
R84 a_109_47.n2 a_109_47.n1 52.431
R85 a_109_47.n4 a_109_47.n3 52.431
R86 a_109_47.n4 a_109_47.n2 38.4
R87 a_109_47.n60 a_109_47.n58 38.4
R88 a_109_47.n7 a_109_47.n5 37.805
R89 a_109_47.n42 a_109_47.n41 37.488
R90 a_109_47.n28 a_109_47.n27 33.918
R91 a_109_47.n56 a_109_47.n4 31.074
R92 a_109_47.n58 a_109_47.n56 31.074
R93 a_109_47.n14 a_109_47.n13 30.348
R94 a_109_47.n57 a_109_47.t8 26.595
R95 a_109_47.n57 a_109_47.t6 26.595
R96 a_109_47.n59 a_109_47.t5 26.595
R97 a_109_47.n59 a_109_47.t4 26.595
R98 a_109_47.t3 a_109_47.n61 26.595
R99 a_109_47.n61 a_109_47.t7 26.595
R100 a_109_47.n0 a_109_47.t10 24.923
R101 a_109_47.n0 a_109_47.t0 24.923
R102 a_109_47.n1 a_109_47.t9 24.923
R103 a_109_47.n1 a_109_47.t2 24.923
R104 a_109_47.n3 a_109_47.t11 24.923
R105 a_109_47.n3 a_109_47.t1 24.923
R106 a_109_47.n45 a_109_47.n44 23.207
R107 a_109_47.n12 a_109_47.n10 21.76
R108 a_109_47.n15 a_109_47.n12 21.76
R109 a_109_47.n18 a_109_47.n15 21.76
R110 a_109_47.n21 a_109_47.n18 21.76
R111 a_109_47.n24 a_109_47.n21 21.76
R112 a_109_47.n26 a_109_47.n24 21.76
R113 a_109_47.n29 a_109_47.n26 21.76
R114 a_109_47.n32 a_109_47.n29 21.76
R115 a_109_47.n35 a_109_47.n32 21.76
R116 a_109_47.n38 a_109_47.n35 21.76
R117 a_109_47.n40 a_109_47.n38 21.76
R118 a_109_47.n43 a_109_47.n40 21.76
R119 a_109_47.n46 a_109_47.n43 21.76
R120 a_109_47.n49 a_109_47.n46 21.76
R121 a_109_47.n52 a_109_47.n49 21.76
R122 a_109_47.n55 a_109_47.n52 21.76
R123 a_109_47.n7 a_109_47.n6 21.46
R124 a_109_47.n56 a_109_47.n55 20.8
R125 a_109_47.n31 a_109_47.n30 19.637
R126 a_109_47.n54 a_109_47.n53 19.637
R127 a_109_47.n9 a_109_47.n8 16.066
R128 a_109_47.n17 a_109_47.n16 16.066
R129 a_109_47.n23 a_109_47.n22 12.496
R130 a_109_47.n37 a_109_47.n36 8.925
R131 a_109_47.n48 a_109_47.n47 8.925
R132 a_109_47.n34 a_109_47.n33 5.355
R133 a_109_47.n51 a_109_47.n50 5.355
R134 a_109_47.n20 a_109_47.n19 1.785
R135 VGND.n0 VGND.t8 197.155
R136 VGND.n2 VGND.n1 116.217
R137 VGND.n8 VGND.n7 116.217
R138 VGND.n12 VGND.n11 116.217
R139 VGND.n18 VGND.n17 116.217
R140 VGND.n24 VGND.n23 116.217
R141 VGND.n30 VGND.n29 116.217
R142 VGND.n36 VGND.n35 116.217
R143 VGND.n40 VGND.n39 116.217
R144 VGND.n46 VGND.n45 116.217
R145 VGND.n52 VGND.n51 116.217
R146 VGND.n57 VGND.t16 114.773
R147 VGND.n1 VGND.t5 24.923
R148 VGND.n1 VGND.t9 24.923
R149 VGND.n7 VGND.t12 24.923
R150 VGND.n7 VGND.t10 24.923
R151 VGND.n11 VGND.t13 24.923
R152 VGND.n11 VGND.t11 24.923
R153 VGND.n17 VGND.t15 24.923
R154 VGND.n17 VGND.t2 24.923
R155 VGND.n23 VGND.t0 24.923
R156 VGND.n23 VGND.t4 24.923
R157 VGND.n29 VGND.t14 24.923
R158 VGND.n29 VGND.t1 24.923
R159 VGND.n35 VGND.t6 24.923
R160 VGND.n35 VGND.t3 24.923
R161 VGND.n39 VGND.t7 24.923
R162 VGND.n39 VGND.t21 24.923
R163 VGND.n45 VGND.t17 24.923
R164 VGND.n45 VGND.t19 24.923
R165 VGND.n51 VGND.t18 24.923
R166 VGND.n51 VGND.t20 24.923
R167 VGND.n9 VGND.n8 17.317
R168 VGND.n41 VGND.n40 15.811
R169 VGND.n37 VGND.n36 12.8
R170 VGND.n3 VGND.n2 11.294
R171 VGND.n13 VGND.n12 11.294
R172 VGND.n47 VGND.n46 9.788
R173 VGND.n58 VGND.n57 6.908
R174 VGND.n31 VGND.n30 6.776
R175 VGND.n19 VGND.n18 5.27
R176 VGND.n4 VGND.n3 4.65
R177 VGND.n6 VGND.n5 4.65
R178 VGND.n10 VGND.n9 4.65
R179 VGND.n14 VGND.n13 4.65
R180 VGND.n16 VGND.n15 4.65
R181 VGND.n20 VGND.n19 4.65
R182 VGND.n22 VGND.n21 4.65
R183 VGND.n26 VGND.n25 4.65
R184 VGND.n28 VGND.n27 4.65
R185 VGND.n32 VGND.n31 4.65
R186 VGND.n34 VGND.n33 4.65
R187 VGND.n38 VGND.n37 4.65
R188 VGND.n42 VGND.n41 4.65
R189 VGND.n44 VGND.n43 4.65
R190 VGND.n48 VGND.n47 4.65
R191 VGND.n50 VGND.n49 4.65
R192 VGND.n54 VGND.n53 4.65
R193 VGND.n56 VGND.n55 4.65
R194 VGND.n53 VGND.n52 3.764
R195 VGND.n25 VGND.n24 0.752
R196 VGND.n4 VGND.n0 0.517
R197 VGND.n6 VGND.n4 0.119
R198 VGND.n10 VGND.n6 0.119
R199 VGND.n14 VGND.n10 0.119
R200 VGND.n16 VGND.n14 0.119
R201 VGND.n20 VGND.n16 0.119
R202 VGND.n22 VGND.n20 0.119
R203 VGND.n26 VGND.n22 0.119
R204 VGND.n28 VGND.n26 0.119
R205 VGND.n32 VGND.n28 0.119
R206 VGND.n34 VGND.n32 0.119
R207 VGND.n38 VGND.n34 0.119
R208 VGND.n42 VGND.n38 0.119
R209 VGND.n44 VGND.n42 0.119
R210 VGND.n48 VGND.n44 0.119
R211 VGND.n50 VGND.n48 0.119
R212 VGND.n54 VGND.n50 0.119
R213 VGND.n56 VGND.n54 0.119
R214 VGND.n58 VGND.n56 0.119
R215 VGND VGND.n58 0.02
R216 VNB VNB.t16 6053.91
R217 VNB.t1 VNB.t4 2030.77
R218 VNB.t5 VNB.t1 2030.77
R219 VNB.t8 VNB.t5 2030.77
R220 VNB.t6 VNB.t8 2030.77
R221 VNB.t9 VNB.t6 2030.77
R222 VNB.t7 VNB.t9 2030.77
R223 VNB.t11 VNB.t7 2030.77
R224 VNB.t14 VNB.t11 2030.77
R225 VNB.t12 VNB.t14 2030.77
R226 VNB.t0 VNB.t12 2030.77
R227 VNB.t10 VNB.t0 2030.77
R228 VNB.t13 VNB.t10 2030.77
R229 VNB.t2 VNB.t13 2030.77
R230 VNB.t15 VNB.t2 2030.77
R231 VNB.t3 VNB.t15 2030.77
R232 VNB.t21 VNB.t3 2030.77
R233 VNB.t17 VNB.t21 2030.77
R234 VNB.t19 VNB.t17 2030.77
R235 VNB.t18 VNB.t19 2030.77
R236 VNB.t20 VNB.t18 2030.77
R237 VNB.t16 VNB.t20 2030.77
R238 VPWR.n0 VPWR.t0 208.281
R239 VPWR.n52 VPWR.n51 174.594
R240 VPWR.n46 VPWR.n45 174.594
R241 VPWR.n40 VPWR.n39 174.594
R242 VPWR.n36 VPWR.n35 174.594
R243 VPWR.n30 VPWR.n29 174.594
R244 VPWR.n24 VPWR.n23 174.594
R245 VPWR.n18 VPWR.n17 174.594
R246 VPWR.n12 VPWR.n11 174.594
R247 VPWR.n8 VPWR.n7 174.594
R248 VPWR.n2 VPWR.n1 174.594
R249 VPWR.n57 VPWR.t16 159.459
R250 VPWR.n51 VPWR.t19 26.595
R251 VPWR.n51 VPWR.t18 26.595
R252 VPWR.n45 VPWR.t21 26.595
R253 VPWR.n45 VPWR.t20 26.595
R254 VPWR.n39 VPWR.t4 26.595
R255 VPWR.n39 VPWR.t17 26.595
R256 VPWR.n35 VPWR.t8 26.595
R257 VPWR.n35 VPWR.t6 26.595
R258 VPWR.n29 VPWR.t10 26.595
R259 VPWR.n29 VPWR.t9 26.595
R260 VPWR.n23 VPWR.t15 26.595
R261 VPWR.n23 VPWR.t11 26.595
R262 VPWR.n17 VPWR.t2 26.595
R263 VPWR.n17 VPWR.t1 26.595
R264 VPWR.n11 VPWR.t5 26.595
R265 VPWR.n11 VPWR.t3 26.595
R266 VPWR.n7 VPWR.t12 26.595
R267 VPWR.n7 VPWR.t7 26.595
R268 VPWR.n1 VPWR.t14 26.595
R269 VPWR.n1 VPWR.t13 26.595
R270 VPWR.n9 VPWR.n8 17.317
R271 VPWR.n41 VPWR.n40 15.811
R272 VPWR.n37 VPWR.n36 12.8
R273 VPWR.n3 VPWR.n2 11.294
R274 VPWR.n13 VPWR.n12 11.294
R275 VPWR.n47 VPWR.n46 9.788
R276 VPWR.n58 VPWR.n57 6.908
R277 VPWR.n31 VPWR.n30 6.776
R278 VPWR.n19 VPWR.n18 5.27
R279 VPWR.n4 VPWR.n3 4.65
R280 VPWR.n6 VPWR.n5 4.65
R281 VPWR.n10 VPWR.n9 4.65
R282 VPWR.n14 VPWR.n13 4.65
R283 VPWR.n16 VPWR.n15 4.65
R284 VPWR.n20 VPWR.n19 4.65
R285 VPWR.n22 VPWR.n21 4.65
R286 VPWR.n26 VPWR.n25 4.65
R287 VPWR.n28 VPWR.n27 4.65
R288 VPWR.n32 VPWR.n31 4.65
R289 VPWR.n34 VPWR.n33 4.65
R290 VPWR.n38 VPWR.n37 4.65
R291 VPWR.n42 VPWR.n41 4.65
R292 VPWR.n44 VPWR.n43 4.65
R293 VPWR.n48 VPWR.n47 4.65
R294 VPWR.n50 VPWR.n49 4.65
R295 VPWR.n54 VPWR.n53 4.65
R296 VPWR.n56 VPWR.n55 4.65
R297 VPWR.n53 VPWR.n52 3.764
R298 VPWR.n25 VPWR.n24 0.752
R299 VPWR.n4 VPWR.n0 0.517
R300 VPWR.n6 VPWR.n4 0.119
R301 VPWR.n10 VPWR.n6 0.119
R302 VPWR.n14 VPWR.n10 0.119
R303 VPWR.n16 VPWR.n14 0.119
R304 VPWR.n20 VPWR.n16 0.119
R305 VPWR.n22 VPWR.n20 0.119
R306 VPWR.n26 VPWR.n22 0.119
R307 VPWR.n28 VPWR.n26 0.119
R308 VPWR.n32 VPWR.n28 0.119
R309 VPWR.n34 VPWR.n32 0.119
R310 VPWR.n38 VPWR.n34 0.119
R311 VPWR.n42 VPWR.n38 0.119
R312 VPWR.n44 VPWR.n42 0.119
R313 VPWR.n48 VPWR.n44 0.119
R314 VPWR.n50 VPWR.n48 0.119
R315 VPWR.n54 VPWR.n50 0.119
R316 VPWR.n56 VPWR.n54 0.119
R317 VPWR.n58 VPWR.n56 0.119
R318 VPWR VPWR.n58 0.02
R319 X.n2 X.n0 146.81
R320 X.n2 X.n1 108.41
R321 X.n4 X.n3 108.41
R322 X.n6 X.n5 108.41
R323 X.n8 X.n7 108.41
R324 X.n10 X.n9 108.41
R325 X.n12 X.n11 108.41
R326 X.n14 X.n13 108.41
R327 X.n17 X.n15 90.831
R328 X.n17 X.n16 52.431
R329 X.n19 X.n18 52.431
R330 X.n21 X.n20 52.431
R331 X.n23 X.n22 52.431
R332 X.n25 X.n24 52.431
R333 X.n27 X.n26 52.431
R334 X.n29 X.n28 52.431
R335 X X.n29 40.47
R336 X.n19 X.n17 38.4
R337 X.n21 X.n19 38.4
R338 X.n23 X.n21 38.4
R339 X.n25 X.n23 38.4
R340 X.n27 X.n25 38.4
R341 X.n29 X.n27 38.4
R342 X.n4 X.n2 38.4
R343 X.n6 X.n4 38.4
R344 X.n8 X.n6 38.4
R345 X.n10 X.n8 38.4
R346 X.n12 X.n10 38.4
R347 X.n14 X.n12 38.4
R348 X X.n14 33.733
R349 X.n0 X.t6 26.595
R350 X.n0 X.t4 26.595
R351 X.n1 X.t9 26.595
R352 X.n1 X.t8 26.595
R353 X.n3 X.t11 26.595
R354 X.n3 X.t10 26.595
R355 X.n5 X.t1 26.595
R356 X.n5 X.t15 26.595
R357 X.n7 X.t3 26.595
R358 X.n7 X.t2 26.595
R359 X.n9 X.t7 26.595
R360 X.n9 X.t5 26.595
R361 X.n11 X.t13 26.595
R362 X.n11 X.t12 26.595
R363 X.n13 X.t0 26.595
R364 X.n13 X.t14 26.595
R365 X.n15 X.t31 24.923
R366 X.n15 X.t19 24.923
R367 X.n16 X.t29 24.923
R368 X.n16 X.t18 24.923
R369 X.n18 X.t16 24.923
R370 X.n18 X.t26 24.923
R371 X.n20 X.t30 24.923
R372 X.n20 X.t28 24.923
R373 X.n22 X.t23 24.923
R374 X.n22 X.t27 24.923
R375 X.n24 X.t22 24.923
R376 X.n24 X.t25 24.923
R377 X.n26 X.t21 24.923
R378 X.n26 X.t24 24.923
R379 X.n28 X.t20 24.923
R380 X.n28 X.t17 24.923
R381 VPB.t14 VPB.t0 248.598
R382 VPB.t13 VPB.t14 248.598
R383 VPB.t12 VPB.t13 248.598
R384 VPB.t7 VPB.t12 248.598
R385 VPB.t5 VPB.t7 248.598
R386 VPB.t3 VPB.t5 248.598
R387 VPB.t2 VPB.t3 248.598
R388 VPB.t1 VPB.t2 248.598
R389 VPB.t15 VPB.t1 248.598
R390 VPB.t11 VPB.t15 248.598
R391 VPB.t10 VPB.t11 248.598
R392 VPB.t9 VPB.t10 248.598
R393 VPB.t8 VPB.t9 248.598
R394 VPB.t6 VPB.t8 248.598
R395 VPB.t4 VPB.t6 248.598
R396 VPB.t17 VPB.t4 248.598
R397 VPB.t21 VPB.t17 248.598
R398 VPB.t20 VPB.t21 248.598
R399 VPB.t19 VPB.t20 248.598
R400 VPB.t18 VPB.t19 248.598
R401 VPB.t16 VPB.t18 248.598
R402 VPB VPB.t16 189.408
C0 VPB VPWR 0.20fF
C1 VPWR VGND 0.23fF
C2 VPWR X 2.21fF
C3 X VGND 1.82fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__bufbuf_8.ext - technology: sky130A

.subckt sky130_fd_sc_hd__bufbuf_8 A X VGND VPWR VNB VPB
X0 a_318_47.t2 a_206_47.t2 VPWR.t9 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 VPWR.t0 a_318_47.t6 X.t10 VPB.t12 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 VPWR.t8 a_206_47.t3 a_318_47.t1 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 X.t2 a_318_47.t7 VGND.t12 VNB.t12 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 X.t9 a_318_47.t8 VPWR.t1 VPB.t11 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 VPWR.t2 a_318_47.t9 X.t8 VPB.t10 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 X.t7 a_318_47.t10 VPWR.t3 VPB.t9 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 VGND.t2 a_206_47.t4 a_318_47.t5 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 VPWR.t4 a_318_47.t11 X.t6 VPB.t8 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 X.t5 a_318_47.t12 VPWR.t5 VPB.t7 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 a_318_47.t4 a_206_47.t5 VGND.t1 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 X.t1 a_318_47.t13 VGND.t11 VNB.t11 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 a_206_47.t0 a_27_47.t2 VGND.t3 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 X.t0 a_318_47.t14 VGND.t10 VNB.t10 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14 a_206_47.t1 a_27_47.t3 VPWR.t10 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 VPWR.t11 a_318_47.t15 X.t4 VPB.t6 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16 VGND.t0 a_206_47.t6 a_318_47.t3 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X17 VGND.t9 a_318_47.t16 X.t15 VNB.t9 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X18 VGND.t8 a_318_47.t17 X.t14 VNB.t8 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X19 VGND.t7 a_318_47.t18 X.t13 VNB.t7 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X20 X.t3 a_318_47.t19 VPWR.t12 VPB.t5 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X21 VGND.t6 a_318_47.t20 X.t12 VNB.t6 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X22 VPWR.t7 a_206_47.t7 a_318_47.t0 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X23 VPWR.t6 A.t0 a_27_47.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X24 VGND.t4 A.t1 a_27_47.t1 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X25 X.t11 a_318_47.t21 VGND.t5 VNB.t5 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
R0 a_206_47.n0 a_206_47.t7 221.719
R1 a_206_47.n2 a_206_47.t2 221.719
R2 a_206_47.n3 a_206_47.t3 221.719
R3 a_206_47.t1 a_206_47.n6 153.428
R4 a_206_47.n0 a_206_47.t6 149.419
R5 a_206_47.n2 a_206_47.t5 149.419
R6 a_206_47.n3 a_206_47.t4 149.419
R7 a_206_47.n6 a_206_47.t0 110.027
R8 a_206_47.n5 a_206_47.n1 97.76
R9 a_206_47.n5 a_206_47.n4 76
R10 a_206_47.n6 a_206_47.n5 53.76
R11 a_206_47.n1 a_206_47.n0 51.77
R12 a_206_47.n4 a_206_47.n2 37.488
R13 a_206_47.n4 a_206_47.n3 37.488
R14 VPWR.n32 VPWR.n31 344.076
R15 VPWR.n0 VPWR.t0 210.284
R16 VPWR.n24 VPWR.n23 174.594
R17 VPWR.n18 VPWR.n17 174.594
R18 VPWR.n12 VPWR.n11 174.594
R19 VPWR.n6 VPWR.n5 174.594
R20 VPWR.n2 VPWR.n1 174.594
R21 VPWR.n31 VPWR.t10 50.601
R22 VPWR.n31 VPWR.t6 41.554
R23 VPWR.n23 VPWR.t9 26.595
R24 VPWR.n23 VPWR.t8 26.595
R25 VPWR.n17 VPWR.t12 26.595
R26 VPWR.n17 VPWR.t7 26.595
R27 VPWR.n11 VPWR.t5 26.595
R28 VPWR.n11 VPWR.t11 26.595
R29 VPWR.n5 VPWR.t3 26.595
R30 VPWR.n5 VPWR.t4 26.595
R31 VPWR.n1 VPWR.t1 26.595
R32 VPWR.n1 VPWR.t2 26.595
R33 VPWR.n3 VPWR.n2 15.435
R34 VPWR.n7 VPWR.n6 13.176
R35 VPWR.n13 VPWR.n12 7.152
R36 VPWR.n25 VPWR.n24 4.894
R37 VPWR.n34 VPWR.n33 4.65
R38 VPWR.n4 VPWR.n3 4.65
R39 VPWR.n8 VPWR.n7 4.65
R40 VPWR.n10 VPWR.n9 4.65
R41 VPWR.n14 VPWR.n13 4.65
R42 VPWR.n16 VPWR.n15 4.65
R43 VPWR.n20 VPWR.n19 4.65
R44 VPWR.n22 VPWR.n21 4.65
R45 VPWR.n26 VPWR.n25 4.65
R46 VPWR.n28 VPWR.n27 4.65
R47 VPWR.n30 VPWR.n29 4.65
R48 VPWR.n19 VPWR.n18 1.129
R49 VPWR.n33 VPWR.n32 0.752
R50 VPWR.n4 VPWR.n0 0.47
R51 VPWR.n8 VPWR.n4 0.119
R52 VPWR.n10 VPWR.n8 0.119
R53 VPWR.n14 VPWR.n10 0.119
R54 VPWR.n16 VPWR.n14 0.119
R55 VPWR.n20 VPWR.n16 0.119
R56 VPWR.n22 VPWR.n20 0.119
R57 VPWR.n26 VPWR.n22 0.119
R58 VPWR.n28 VPWR.n26 0.119
R59 VPWR.n30 VPWR.n28 0.119
R60 VPWR.n34 VPWR.n30 0.119
R61 VPWR.n35 VPWR.n34 0.119
R62 VPWR VPWR.n35 0.02
R63 a_318_47.n2 a_318_47.t6 221.719
R64 a_318_47.n3 a_318_47.t8 221.719
R65 a_318_47.n4 a_318_47.t9 221.719
R66 a_318_47.n6 a_318_47.t10 221.719
R67 a_318_47.n9 a_318_47.t11 221.719
R68 a_318_47.n12 a_318_47.t12 221.719
R69 a_318_47.n15 a_318_47.t15 221.719
R70 a_318_47.n18 a_318_47.t19 221.719
R71 a_318_47.n22 a_318_47.t1 173.405
R72 a_318_47.n2 a_318_47.t18 149.419
R73 a_318_47.n3 a_318_47.t21 149.419
R74 a_318_47.n4 a_318_47.t16 149.419
R75 a_318_47.n6 a_318_47.t7 149.419
R76 a_318_47.n9 a_318_47.t20 149.419
R77 a_318_47.n12 a_318_47.t14 149.419
R78 a_318_47.n15 a_318_47.t17 149.419
R79 a_318_47.n18 a_318_47.t13 149.419
R80 a_318_47.n1 a_318_47.t5 130.27
R81 a_318_47.n23 a_318_47.n22 108.41
R82 a_318_47.n8 a_318_47.n5 97.76
R83 a_318_47.n20 a_318_47.n19 76
R84 a_318_47.n8 a_318_47.n7 76
R85 a_318_47.n11 a_318_47.n10 76
R86 a_318_47.n14 a_318_47.n13 76
R87 a_318_47.n17 a_318_47.n16 76
R88 a_318_47.n3 a_318_47.n2 74.977
R89 a_318_47.n4 a_318_47.n3 74.977
R90 a_318_47.n1 a_318_47.n0 52.431
R91 a_318_47.n5 a_318_47.n4 48.2
R92 a_318_47.n7 a_318_47.n6 33.918
R93 a_318_47.n21 a_318_47.n1 32
R94 a_318_47.n22 a_318_47.n21 32
R95 a_318_47.n23 a_318_47.t0 26.595
R96 a_318_47.t2 a_318_47.n23 26.595
R97 a_318_47.n0 a_318_47.t3 24.923
R98 a_318_47.n0 a_318_47.t4 24.923
R99 a_318_47.n19 a_318_47.n18 23.207
R100 a_318_47.n11 a_318_47.n8 21.76
R101 a_318_47.n14 a_318_47.n11 21.76
R102 a_318_47.n17 a_318_47.n14 21.76
R103 a_318_47.n20 a_318_47.n17 21.76
R104 a_318_47.n21 a_318_47.n20 21.76
R105 a_318_47.n10 a_318_47.n9 19.637
R106 a_318_47.n16 a_318_47.n15 8.925
R107 a_318_47.n13 a_318_47.n12 5.355
R108 VPB.t4 VPB.t2 574.143
R109 VPB.t0 VPB.t4 287.071
R110 VPB.t11 VPB.t12 248.598
R111 VPB.t10 VPB.t11 248.598
R112 VPB.t9 VPB.t10 248.598
R113 VPB.t8 VPB.t9 248.598
R114 VPB.t7 VPB.t8 248.598
R115 VPB.t6 VPB.t7 248.598
R116 VPB.t5 VPB.t6 248.598
R117 VPB.t1 VPB.t5 248.598
R118 VPB.t3 VPB.t1 248.598
R119 VPB.t2 VPB.t3 248.598
R120 VPB VPB.t0 189.408
R121 X.n2 X.n0 146.81
R122 X.n2 X.n1 108.41
R123 X.n4 X.n3 108.41
R124 X.n6 X.n5 108.41
R125 X.n9 X.n7 90.831
R126 X.n9 X.n8 52.431
R127 X.n11 X.n10 52.431
R128 X.n13 X.n12 52.431
R129 X.n11 X.n9 38.4
R130 X.n13 X.n11 38.4
R131 X.n4 X.n2 38.4
R132 X.n6 X.n4 38.4
R133 X X.n13 36.329
R134 X X.n6 29.592
R135 X.n0 X.t4 26.595
R136 X.n0 X.t3 26.595
R137 X.n1 X.t6 26.595
R138 X.n1 X.t5 26.595
R139 X.n3 X.t8 26.595
R140 X.n3 X.t7 26.595
R141 X.n5 X.t10 26.595
R142 X.n5 X.t9 26.595
R143 X.n7 X.t14 24.923
R144 X.n7 X.t1 24.923
R145 X.n8 X.t12 24.923
R146 X.n8 X.t0 24.923
R147 X.n10 X.t15 24.923
R148 X.n10 X.t2 24.923
R149 X.n12 X.t13 24.923
R150 X.n12 X.t11 24.923
R151 VGND.n0 VGND.t7 199.159
R152 VGND.n2 VGND.n1 116.217
R153 VGND.n6 VGND.n5 116.217
R154 VGND.n12 VGND.n11 116.217
R155 VGND.n18 VGND.n17 116.217
R156 VGND.n24 VGND.n23 116.217
R157 VGND.n32 VGND.n31 116.217
R158 VGND.n31 VGND.t3 44
R159 VGND.n31 VGND.t4 38.571
R160 VGND.n1 VGND.t5 24.923
R161 VGND.n1 VGND.t9 24.923
R162 VGND.n5 VGND.t12 24.923
R163 VGND.n5 VGND.t6 24.923
R164 VGND.n11 VGND.t10 24.923
R165 VGND.n11 VGND.t8 24.923
R166 VGND.n17 VGND.t11 24.923
R167 VGND.n17 VGND.t0 24.923
R168 VGND.n23 VGND.t1 24.923
R169 VGND.n23 VGND.t2 24.923
R170 VGND.n3 VGND.n2 15.435
R171 VGND.n7 VGND.n6 13.176
R172 VGND.n13 VGND.n12 7.152
R173 VGND.n25 VGND.n24 4.894
R174 VGND.n4 VGND.n3 4.65
R175 VGND.n8 VGND.n7 4.65
R176 VGND.n10 VGND.n9 4.65
R177 VGND.n14 VGND.n13 4.65
R178 VGND.n16 VGND.n15 4.65
R179 VGND.n20 VGND.n19 4.65
R180 VGND.n22 VGND.n21 4.65
R181 VGND.n26 VGND.n25 4.65
R182 VGND.n28 VGND.n27 4.65
R183 VGND.n30 VGND.n29 4.65
R184 VGND.n34 VGND.n33 4.65
R185 VGND.n19 VGND.n18 1.129
R186 VGND.n33 VGND.n32 0.752
R187 VGND.n4 VGND.n0 0.47
R188 VGND.n8 VGND.n4 0.119
R189 VGND.n10 VGND.n8 0.119
R190 VGND.n14 VGND.n10 0.119
R191 VGND.n16 VGND.n14 0.119
R192 VGND.n20 VGND.n16 0.119
R193 VGND.n22 VGND.n20 0.119
R194 VGND.n26 VGND.n22 0.119
R195 VGND.n28 VGND.n26 0.119
R196 VGND.n30 VGND.n28 0.119
R197 VGND.n34 VGND.n30 0.119
R198 VGND.n35 VGND.n34 0.119
R199 VGND VGND.n35 0.02
R200 VNB VNB.t4 6438.23
R201 VNB.t3 VNB.t2 4690.11
R202 VNB.t4 VNB.t3 2303.7
R203 VNB.t5 VNB.t7 2030.77
R204 VNB.t9 VNB.t5 2030.77
R205 VNB.t12 VNB.t9 2030.77
R206 VNB.t6 VNB.t12 2030.77
R207 VNB.t10 VNB.t6 2030.77
R208 VNB.t8 VNB.t10 2030.77
R209 VNB.t11 VNB.t8 2030.77
R210 VNB.t0 VNB.t11 2030.77
R211 VNB.t1 VNB.t0 2030.77
R212 VNB.t2 VNB.t1 2030.77
R213 a_27_47.t0 a_27_47.n1 252.095
R214 a_27_47.n0 a_27_47.t3 239.984
R215 a_27_47.n1 a_27_47.t1 176.662
R216 a_27_47.n0 a_27_47.t2 167.684
R217 a_27_47.n1 a_27_47.n0 76
R218 A.n0 A.t1 195.015
R219 A.n0 A.t0 172.521
R220 A A.n0 84
C0 VPWR VPB 0.15fF
C1 X VGND 0.89fF
C2 VPWR VGND 0.15fF
C3 VPWR X 1.08fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__bufbuf_16.ext - technology: sky130A

.subckt sky130_fd_sc_hd__bufbuf_16 A X VGND VPWR VNB VPB
X0 X.t15 a_549_47.t12 VPWR.t14 VPB.t20 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 X.t28 a_549_47.t13 VGND.t17 VNB.t17 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 VPWR.t24 a_215_47.t6 a_549_47.t5 VPB.t24 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 VGND.t18 a_109_47.t2 a_215_47.t0 VNB.t18 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 X.t14 a_549_47.t14 VPWR.t13 VPB.t19 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 VGND.t19 a_109_47.t3 a_215_47.t1 VNB.t19 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 VGND.t21 a_215_47.t7 a_549_47.t6 VNB.t21 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 a_549_47.t7 a_215_47.t8 VPWR.t25 VPB.t25 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 VPWR.t12 a_549_47.t15 X.t13 VPB.t18 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 VGND.t22 a_215_47.t9 a_549_47.t8 VNB.t22 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 VGND.t16 a_549_47.t16 X.t27 VNB.t16 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 VGND.t15 a_549_47.t17 X.t26 VNB.t15 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 X.t12 a_549_47.t18 VPWR.t11 VPB.t17 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13 X.t25 a_549_47.t19 VGND.t14 VNB.t14 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14 a_549_47.t9 a_215_47.t10 VGND.t23 VNB.t23 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X15 VPWR.t10 a_549_47.t20 X.t11 VPB.t16 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16 X.t24 a_549_47.t21 VGND.t13 VNB.t13 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X17 VPWR.t9 a_549_47.t22 X.t10 VPB.t15 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X18 X.t9 a_549_47.t23 VPWR.t8 VPB.t14 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X19 a_549_47.t10 a_215_47.t11 VGND.t24 VNB.t24 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X20 a_549_47.t11 a_215_47.t12 VGND.t25 VNB.t25 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X21 X.t23 a_549_47.t24 VGND.t12 VNB.t12 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X22 X.t8 a_549_47.t25 VPWR.t7 VPB.t13 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X23 VPWR.t0 a_215_47.t13 a_549_47.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X24 VPWR.t6 a_549_47.t26 X.t7 VPB.t12 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X25 VGND.t11 a_549_47.t27 X.t22 VNB.t11 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X26 VPWR.t5 a_549_47.t28 X.t6 VPB.t11 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X27 a_549_47.t1 a_215_47.t14 VPWR.t1 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X28 X.t5 a_549_47.t29 VPWR.t20 VPB.t10 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X29 VGND.t10 a_549_47.t30 X.t21 VNB.t10 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X30 VGND.t9 a_549_47.t31 X.t20 VNB.t9 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X31 X.t4 a_549_47.t32 VPWR.t19 VPB.t9 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X32 VGND.t0 a_215_47.t15 a_549_47.t2 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X33 VGND.t8 a_549_47.t33 X.t19 VNB.t8 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X34 VGND.t7 a_549_47.t34 X.t18 VNB.t7 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X35 VPWR.t21 a_109_47.t4 a_215_47.t2 VPB.t21 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X36 VGND.t6 a_549_47.t35 X.t17 VNB.t6 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X37 a_215_47.t3 a_109_47.t5 VPWR.t22 VPB.t22 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X38 VPWR.t18 a_549_47.t36 X.t3 VPB.t8 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X39 X.t16 a_549_47.t37 VGND.t5 VNB.t5 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X40 a_215_47.t4 a_109_47.t6 VGND.t20 VNB.t20 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X41 VPWR.t23 a_109_47.t7 a_215_47.t5 VPB.t23 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X42 X.t2 a_549_47.t38 VPWR.t17 VPB.t7 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X43 VPWR.t2 a_215_47.t16 a_549_47.t3 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X44 X.t31 a_549_47.t39 VGND.t4 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X45 X.t30 a_549_47.t40 VGND.t3 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X46 a_109_47.t0 A.t0 VPWR.t4 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X47 VPWR.t16 a_549_47.t41 X.t1 VPB.t6 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X48 a_549_47.t4 a_215_47.t17 VPWR.t3 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X49 VPWR.t15 a_549_47.t42 X.t0 VPB.t5 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X50 a_109_47.t1 A.t1 VGND.t1 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X51 X.t29 a_549_47.t43 VGND.t2 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
R0 a_549_47.n5 a_549_47.t26 221.719
R1 a_549_47.n6 a_549_47.t29 221.719
R2 a_549_47.n8 a_549_47.t41 221.719
R3 a_549_47.n13 a_549_47.t12 221.719
R4 a_549_47.n16 a_549_47.t22 221.719
R5 a_549_47.n19 a_549_47.t25 221.719
R6 a_549_47.n22 a_549_47.t28 221.719
R7 a_549_47.n27 a_549_47.t32 221.719
R8 a_549_47.n30 a_549_47.t42 221.719
R9 a_549_47.n33 a_549_47.t14 221.719
R10 a_549_47.n36 a_549_47.t15 221.719
R11 a_549_47.n41 a_549_47.t18 221.719
R12 a_549_47.n44 a_549_47.t20 221.719
R13 a_549_47.n47 a_549_47.t23 221.719
R14 a_549_47.n50 a_549_47.t36 221.719
R15 a_549_47.n53 a_549_47.t38 221.719
R16 a_549_47.n5 a_549_47.t31 149.419
R17 a_549_47.n6 a_549_47.t37 149.419
R18 a_549_47.n8 a_549_47.t27 149.419
R19 a_549_47.n13 a_549_47.t19 149.419
R20 a_549_47.n16 a_549_47.t17 149.419
R21 a_549_47.n19 a_549_47.t13 149.419
R22 a_549_47.n22 a_549_47.t16 149.419
R23 a_549_47.n27 a_549_47.t43 149.419
R24 a_549_47.n30 a_549_47.t35 149.419
R25 a_549_47.n33 a_549_47.t40 149.419
R26 a_549_47.n36 a_549_47.t34 149.419
R27 a_549_47.n41 a_549_47.t39 149.419
R28 a_549_47.n44 a_549_47.t33 149.419
R29 a_549_47.n47 a_549_47.t24 149.419
R30 a_549_47.n50 a_549_47.t30 149.419
R31 a_549_47.n53 a_549_47.t21 149.419
R32 a_549_47.n61 a_549_47.n60 146.811
R33 a_549_47.n58 a_549_47.n57 108.41
R34 a_549_47.n60 a_549_47.n59 108.41
R35 a_549_47.n10 a_549_47.n7 97.76
R36 a_549_47.n2 a_549_47.n0 90.831
R37 a_549_47.n55 a_549_47.n54 76
R38 a_549_47.n10 a_549_47.n9 76
R39 a_549_47.n12 a_549_47.n11 76
R40 a_549_47.n15 a_549_47.n14 76
R41 a_549_47.n18 a_549_47.n17 76
R42 a_549_47.n21 a_549_47.n20 76
R43 a_549_47.n24 a_549_47.n23 76
R44 a_549_47.n26 a_549_47.n25 76
R45 a_549_47.n29 a_549_47.n28 76
R46 a_549_47.n32 a_549_47.n31 76
R47 a_549_47.n35 a_549_47.n34 76
R48 a_549_47.n38 a_549_47.n37 76
R49 a_549_47.n40 a_549_47.n39 76
R50 a_549_47.n43 a_549_47.n42 76
R51 a_549_47.n46 a_549_47.n45 76
R52 a_549_47.n49 a_549_47.n48 76
R53 a_549_47.n52 a_549_47.n51 76
R54 a_549_47.n7 a_549_47.n5 73.192
R55 a_549_47.n2 a_549_47.n1 52.431
R56 a_549_47.n4 a_549_47.n3 52.431
R57 a_549_47.n4 a_549_47.n2 38.4
R58 a_549_47.n60 a_549_47.n58 38.4
R59 a_549_47.n42 a_549_47.n41 37.488
R60 a_549_47.n28 a_549_47.n27 33.918
R61 a_549_47.n56 a_549_47.n4 31.074
R62 a_549_47.n58 a_549_47.n56 31.074
R63 a_549_47.n14 a_549_47.n13 30.348
R64 a_549_47.n57 a_549_47.t3 26.595
R65 a_549_47.n57 a_549_47.t4 26.595
R66 a_549_47.n59 a_549_47.t5 26.595
R67 a_549_47.n59 a_549_47.t7 26.595
R68 a_549_47.t0 a_549_47.n61 26.595
R69 a_549_47.n61 a_549_47.t1 26.595
R70 a_549_47.n0 a_549_47.t6 24.923
R71 a_549_47.n0 a_549_47.t9 24.923
R72 a_549_47.n1 a_549_47.t8 24.923
R73 a_549_47.n1 a_549_47.t10 24.923
R74 a_549_47.n3 a_549_47.t2 24.923
R75 a_549_47.n3 a_549_47.t11 24.923
R76 a_549_47.n45 a_549_47.n44 23.207
R77 a_549_47.n12 a_549_47.n10 21.76
R78 a_549_47.n15 a_549_47.n12 21.76
R79 a_549_47.n18 a_549_47.n15 21.76
R80 a_549_47.n21 a_549_47.n18 21.76
R81 a_549_47.n24 a_549_47.n21 21.76
R82 a_549_47.n26 a_549_47.n24 21.76
R83 a_549_47.n29 a_549_47.n26 21.76
R84 a_549_47.n32 a_549_47.n29 21.76
R85 a_549_47.n35 a_549_47.n32 21.76
R86 a_549_47.n38 a_549_47.n35 21.76
R87 a_549_47.n40 a_549_47.n38 21.76
R88 a_549_47.n43 a_549_47.n40 21.76
R89 a_549_47.n46 a_549_47.n43 21.76
R90 a_549_47.n49 a_549_47.n46 21.76
R91 a_549_47.n52 a_549_47.n49 21.76
R92 a_549_47.n55 a_549_47.n52 21.76
R93 a_549_47.n56 a_549_47.n55 20.8
R94 a_549_47.n31 a_549_47.n30 19.637
R95 a_549_47.n54 a_549_47.n53 19.637
R96 a_549_47.n9 a_549_47.n8 16.066
R97 a_549_47.n17 a_549_47.n16 16.066
R98 a_549_47.n23 a_549_47.n22 12.496
R99 a_549_47.n37 a_549_47.n36 8.925
R100 a_549_47.n48 a_549_47.n47 8.925
R101 a_549_47.n34 a_549_47.n33 5.355
R102 a_549_47.n51 a_549_47.n50 5.355
R103 a_549_47.n7 a_549_47.n6 1.785
R104 a_549_47.n20 a_549_47.n19 1.785
R105 VPWR.n0 VPWR.t6 206.354
R106 VPWR.n64 VPWR.n63 174.594
R107 VPWR.n58 VPWR.n57 174.594
R108 VPWR.n52 VPWR.n51 174.594
R109 VPWR.n48 VPWR.n47 174.594
R110 VPWR.n42 VPWR.n41 174.594
R111 VPWR.n36 VPWR.n35 174.594
R112 VPWR.n30 VPWR.n29 174.594
R113 VPWR.n24 VPWR.n23 174.594
R114 VPWR.n18 VPWR.n17 174.594
R115 VPWR.n14 VPWR.n13 174.594
R116 VPWR.n8 VPWR.n7 174.594
R117 VPWR.n2 VPWR.n1 174.594
R118 VPWR.n71 VPWR.t4 159.459
R119 VPWR.n63 VPWR.t22 26.595
R120 VPWR.n63 VPWR.t23 26.595
R121 VPWR.n57 VPWR.t1 26.595
R122 VPWR.n57 VPWR.t21 26.595
R123 VPWR.n51 VPWR.t25 26.595
R124 VPWR.n51 VPWR.t0 26.595
R125 VPWR.n47 VPWR.t3 26.595
R126 VPWR.n47 VPWR.t24 26.595
R127 VPWR.n41 VPWR.t17 26.595
R128 VPWR.n41 VPWR.t2 26.595
R129 VPWR.n35 VPWR.t8 26.595
R130 VPWR.n35 VPWR.t18 26.595
R131 VPWR.n29 VPWR.t11 26.595
R132 VPWR.n29 VPWR.t10 26.595
R133 VPWR.n23 VPWR.t13 26.595
R134 VPWR.n23 VPWR.t12 26.595
R135 VPWR.n17 VPWR.t19 26.595
R136 VPWR.n17 VPWR.t15 26.595
R137 VPWR.n13 VPWR.t7 26.595
R138 VPWR.n13 VPWR.t5 26.595
R139 VPWR.n7 VPWR.t14 26.595
R140 VPWR.n7 VPWR.t9 26.595
R141 VPWR.n1 VPWR.t20 26.595
R142 VPWR.n1 VPWR.t16 26.595
R143 VPWR.n49 VPWR.n48 17.317
R144 VPWR.n15 VPWR.n14 15.811
R145 VPWR.n19 VPWR.n18 12.8
R146 VPWR.n43 VPWR.n42 11.294
R147 VPWR.n53 VPWR.n52 11.294
R148 VPWR.n9 VPWR.n8 9.788
R149 VPWR.n72 VPWR.n71 6.908
R150 VPWR.n25 VPWR.n24 6.776
R151 VPWR.n37 VPWR.n36 5.27
R152 VPWR.n59 VPWR.n58 5.27
R153 VPWR.n4 VPWR.n3 4.65
R154 VPWR.n6 VPWR.n5 4.65
R155 VPWR.n10 VPWR.n9 4.65
R156 VPWR.n12 VPWR.n11 4.65
R157 VPWR.n16 VPWR.n15 4.65
R158 VPWR.n20 VPWR.n19 4.65
R159 VPWR.n22 VPWR.n21 4.65
R160 VPWR.n26 VPWR.n25 4.65
R161 VPWR.n28 VPWR.n27 4.65
R162 VPWR.n32 VPWR.n31 4.65
R163 VPWR.n34 VPWR.n33 4.65
R164 VPWR.n38 VPWR.n37 4.65
R165 VPWR.n40 VPWR.n39 4.65
R166 VPWR.n44 VPWR.n43 4.65
R167 VPWR.n46 VPWR.n45 4.65
R168 VPWR.n50 VPWR.n49 4.65
R169 VPWR.n54 VPWR.n53 4.65
R170 VPWR.n56 VPWR.n55 4.65
R171 VPWR.n60 VPWR.n59 4.65
R172 VPWR.n62 VPWR.n61 4.65
R173 VPWR.n66 VPWR.n65 4.65
R174 VPWR.n68 VPWR.n67 4.65
R175 VPWR.n70 VPWR.n69 4.65
R176 VPWR.n3 VPWR.n2 3.764
R177 VPWR.n4 VPWR.n0 0.861
R178 VPWR.n31 VPWR.n30 0.752
R179 VPWR.n65 VPWR.n64 0.752
R180 VPWR.n6 VPWR.n4 0.119
R181 VPWR.n10 VPWR.n6 0.119
R182 VPWR.n12 VPWR.n10 0.119
R183 VPWR.n16 VPWR.n12 0.119
R184 VPWR.n20 VPWR.n16 0.119
R185 VPWR.n22 VPWR.n20 0.119
R186 VPWR.n26 VPWR.n22 0.119
R187 VPWR.n28 VPWR.n26 0.119
R188 VPWR.n32 VPWR.n28 0.119
R189 VPWR.n34 VPWR.n32 0.119
R190 VPWR.n38 VPWR.n34 0.119
R191 VPWR.n40 VPWR.n38 0.119
R192 VPWR.n44 VPWR.n40 0.119
R193 VPWR.n46 VPWR.n44 0.119
R194 VPWR.n50 VPWR.n46 0.119
R195 VPWR.n54 VPWR.n50 0.119
R196 VPWR.n56 VPWR.n54 0.119
R197 VPWR.n60 VPWR.n56 0.119
R198 VPWR.n62 VPWR.n60 0.119
R199 VPWR.n66 VPWR.n62 0.119
R200 VPWR.n68 VPWR.n66 0.119
R201 VPWR.n70 VPWR.n68 0.119
R202 VPWR.n72 VPWR.n70 0.119
R203 VPWR VPWR.n72 0.02
R204 X.n2 X.n0 146.81
R205 X.n2 X.n1 108.41
R206 X.n4 X.n3 108.41
R207 X.n6 X.n5 108.41
R208 X.n8 X.n7 108.41
R209 X.n10 X.n9 108.41
R210 X.n12 X.n11 108.41
R211 X.n14 X.n13 108.41
R212 X.n17 X.n15 90.831
R213 X.n17 X.n16 52.431
R214 X.n19 X.n18 52.431
R215 X.n21 X.n20 52.431
R216 X.n23 X.n22 52.431
R217 X.n25 X.n24 52.431
R218 X.n27 X.n26 52.431
R219 X.n29 X.n28 52.431
R220 X.n19 X.n17 38.4
R221 X.n21 X.n19 38.4
R222 X.n23 X.n21 38.4
R223 X.n25 X.n23 38.4
R224 X.n27 X.n25 38.4
R225 X.n29 X.n27 38.4
R226 X.n4 X.n2 38.4
R227 X.n6 X.n4 38.4
R228 X.n8 X.n6 38.4
R229 X.n10 X.n8 38.4
R230 X.n12 X.n10 38.4
R231 X.n14 X.n12 38.4
R232 X X.n29 27.481
R233 X.n0 X.t3 26.595
R234 X.n0 X.t2 26.595
R235 X.n1 X.t11 26.595
R236 X.n1 X.t9 26.595
R237 X.n3 X.t13 26.595
R238 X.n3 X.t12 26.595
R239 X.n5 X.t0 26.595
R240 X.n5 X.t14 26.595
R241 X.n7 X.t6 26.595
R242 X.n7 X.t4 26.595
R243 X.n9 X.t10 26.595
R244 X.n9 X.t8 26.595
R245 X.n11 X.t1 26.595
R246 X.n11 X.t15 26.595
R247 X.n13 X.t7 26.595
R248 X.n13 X.t5 26.595
R249 X.n15 X.t21 24.923
R250 X.n15 X.t24 24.923
R251 X.n16 X.t19 24.923
R252 X.n16 X.t23 24.923
R253 X.n18 X.t18 24.923
R254 X.n18 X.t31 24.923
R255 X.n20 X.t17 24.923
R256 X.n20 X.t30 24.923
R257 X.n22 X.t27 24.923
R258 X.n22 X.t29 24.923
R259 X.n24 X.t26 24.923
R260 X.n24 X.t28 24.923
R261 X.n26 X.t22 24.923
R262 X.n26 X.t25 24.923
R263 X.n28 X.t20 24.923
R264 X.n28 X.t16 24.923
R265 X X.n14 17.442
R266 VPB.t4 VPB.t23 556.386
R267 VPB.t10 VPB.t12 248.598
R268 VPB.t6 VPB.t10 248.598
R269 VPB.t20 VPB.t6 248.598
R270 VPB.t15 VPB.t20 248.598
R271 VPB.t13 VPB.t15 248.598
R272 VPB.t11 VPB.t13 248.598
R273 VPB.t9 VPB.t11 248.598
R274 VPB.t5 VPB.t9 248.598
R275 VPB.t19 VPB.t5 248.598
R276 VPB.t18 VPB.t19 248.598
R277 VPB.t17 VPB.t18 248.598
R278 VPB.t16 VPB.t17 248.598
R279 VPB.t14 VPB.t16 248.598
R280 VPB.t8 VPB.t14 248.598
R281 VPB.t7 VPB.t8 248.598
R282 VPB.t2 VPB.t7 248.598
R283 VPB.t3 VPB.t2 248.598
R284 VPB.t24 VPB.t3 248.598
R285 VPB.t25 VPB.t24 248.598
R286 VPB.t0 VPB.t25 248.598
R287 VPB.t1 VPB.t0 248.598
R288 VPB.t21 VPB.t1 248.598
R289 VPB.t22 VPB.t21 248.598
R290 VPB.t23 VPB.t22 248.598
R291 VPB VPB.t4 189.408
R292 VGND.n0 VGND.t9 195.229
R293 VGND.n2 VGND.n1 116.217
R294 VGND.n8 VGND.n7 116.217
R295 VGND.n14 VGND.n13 116.217
R296 VGND.n18 VGND.n17 116.217
R297 VGND.n24 VGND.n23 116.217
R298 VGND.n30 VGND.n29 116.217
R299 VGND.n36 VGND.n35 116.217
R300 VGND.n42 VGND.n41 116.217
R301 VGND.n48 VGND.n47 116.217
R302 VGND.n52 VGND.n51 116.217
R303 VGND.n58 VGND.n57 116.217
R304 VGND.n64 VGND.n63 116.217
R305 VGND.n71 VGND.t1 114.773
R306 VGND.n1 VGND.t5 24.923
R307 VGND.n1 VGND.t11 24.923
R308 VGND.n7 VGND.t14 24.923
R309 VGND.n7 VGND.t15 24.923
R310 VGND.n13 VGND.t17 24.923
R311 VGND.n13 VGND.t16 24.923
R312 VGND.n17 VGND.t2 24.923
R313 VGND.n17 VGND.t6 24.923
R314 VGND.n23 VGND.t3 24.923
R315 VGND.n23 VGND.t7 24.923
R316 VGND.n29 VGND.t4 24.923
R317 VGND.n29 VGND.t8 24.923
R318 VGND.n35 VGND.t12 24.923
R319 VGND.n35 VGND.t10 24.923
R320 VGND.n41 VGND.t13 24.923
R321 VGND.n41 VGND.t0 24.923
R322 VGND.n47 VGND.t25 24.923
R323 VGND.n47 VGND.t22 24.923
R324 VGND.n51 VGND.t24 24.923
R325 VGND.n51 VGND.t21 24.923
R326 VGND.n57 VGND.t23 24.923
R327 VGND.n57 VGND.t19 24.923
R328 VGND.n63 VGND.t20 24.923
R329 VGND.n63 VGND.t18 24.923
R330 VGND.n49 VGND.n48 17.317
R331 VGND.n15 VGND.n14 15.811
R332 VGND.n19 VGND.n18 12.8
R333 VGND.n43 VGND.n42 11.294
R334 VGND.n53 VGND.n52 11.294
R335 VGND.n9 VGND.n8 9.788
R336 VGND.n72 VGND.n71 6.908
R337 VGND.n25 VGND.n24 6.776
R338 VGND.n37 VGND.n36 5.27
R339 VGND.n59 VGND.n58 5.27
R340 VGND.n4 VGND.n3 4.65
R341 VGND.n6 VGND.n5 4.65
R342 VGND.n10 VGND.n9 4.65
R343 VGND.n12 VGND.n11 4.65
R344 VGND.n16 VGND.n15 4.65
R345 VGND.n20 VGND.n19 4.65
R346 VGND.n22 VGND.n21 4.65
R347 VGND.n26 VGND.n25 4.65
R348 VGND.n28 VGND.n27 4.65
R349 VGND.n32 VGND.n31 4.65
R350 VGND.n34 VGND.n33 4.65
R351 VGND.n38 VGND.n37 4.65
R352 VGND.n40 VGND.n39 4.65
R353 VGND.n44 VGND.n43 4.65
R354 VGND.n46 VGND.n45 4.65
R355 VGND.n50 VGND.n49 4.65
R356 VGND.n54 VGND.n53 4.65
R357 VGND.n56 VGND.n55 4.65
R358 VGND.n60 VGND.n59 4.65
R359 VGND.n62 VGND.n61 4.65
R360 VGND.n66 VGND.n65 4.65
R361 VGND.n68 VGND.n67 4.65
R362 VGND.n70 VGND.n69 4.65
R363 VGND.n3 VGND.n2 3.764
R364 VGND.n4 VGND.n0 0.861
R365 VGND.n31 VGND.n30 0.752
R366 VGND.n65 VGND.n64 0.752
R367 VGND.n6 VGND.n4 0.119
R368 VGND.n10 VGND.n6 0.119
R369 VGND.n12 VGND.n10 0.119
R370 VGND.n16 VGND.n12 0.119
R371 VGND.n20 VGND.n16 0.119
R372 VGND.n22 VGND.n20 0.119
R373 VGND.n26 VGND.n22 0.119
R374 VGND.n28 VGND.n26 0.119
R375 VGND.n32 VGND.n28 0.119
R376 VGND.n34 VGND.n32 0.119
R377 VGND.n38 VGND.n34 0.119
R378 VGND.n40 VGND.n38 0.119
R379 VGND.n44 VGND.n40 0.119
R380 VGND.n46 VGND.n44 0.119
R381 VGND.n50 VGND.n46 0.119
R382 VGND.n54 VGND.n50 0.119
R383 VGND.n56 VGND.n54 0.119
R384 VGND.n60 VGND.n56 0.119
R385 VGND.n62 VGND.n60 0.119
R386 VGND.n66 VGND.n62 0.119
R387 VGND.n68 VGND.n66 0.119
R388 VGND.n70 VGND.n68 0.119
R389 VGND.n72 VGND.n70 0.119
R390 VGND VGND.n72 0.02
R391 VNB VNB.t1 6053.91
R392 VNB.t1 VNB.t18 4545.05
R393 VNB.t5 VNB.t9 2030.77
R394 VNB.t11 VNB.t5 2030.77
R395 VNB.t14 VNB.t11 2030.77
R396 VNB.t15 VNB.t14 2030.77
R397 VNB.t17 VNB.t15 2030.77
R398 VNB.t16 VNB.t17 2030.77
R399 VNB.t2 VNB.t16 2030.77
R400 VNB.t6 VNB.t2 2030.77
R401 VNB.t3 VNB.t6 2030.77
R402 VNB.t7 VNB.t3 2030.77
R403 VNB.t4 VNB.t7 2030.77
R404 VNB.t8 VNB.t4 2030.77
R405 VNB.t12 VNB.t8 2030.77
R406 VNB.t10 VNB.t12 2030.77
R407 VNB.t13 VNB.t10 2030.77
R408 VNB.t0 VNB.t13 2030.77
R409 VNB.t25 VNB.t0 2030.77
R410 VNB.t22 VNB.t25 2030.77
R411 VNB.t24 VNB.t22 2030.77
R412 VNB.t21 VNB.t24 2030.77
R413 VNB.t23 VNB.t21 2030.77
R414 VNB.t19 VNB.t23 2030.77
R415 VNB.t20 VNB.t19 2030.77
R416 VNB.t18 VNB.t20 2030.77
R417 a_215_47.n2 a_215_47.t16 221.719
R418 a_215_47.n4 a_215_47.t17 221.719
R419 a_215_47.n7 a_215_47.t6 221.719
R420 a_215_47.n10 a_215_47.t8 221.719
R421 a_215_47.n13 a_215_47.t13 221.719
R422 a_215_47.n16 a_215_47.t14 221.719
R423 a_215_47.n20 a_215_47.t5 173.405
R424 a_215_47.n2 a_215_47.t15 149.419
R425 a_215_47.n4 a_215_47.t12 149.419
R426 a_215_47.n7 a_215_47.t9 149.419
R427 a_215_47.n10 a_215_47.t11 149.419
R428 a_215_47.n13 a_215_47.t7 149.419
R429 a_215_47.n16 a_215_47.t10 149.419
R430 a_215_47.n1 a_215_47.t0 130.27
R431 a_215_47.n21 a_215_47.n20 108.41
R432 a_215_47.n6 a_215_47.n3 97.76
R433 a_215_47.n18 a_215_47.n17 76
R434 a_215_47.n6 a_215_47.n5 76
R435 a_215_47.n9 a_215_47.n8 76
R436 a_215_47.n12 a_215_47.n11 76
R437 a_215_47.n15 a_215_47.n14 76
R438 a_215_47.n1 a_215_47.n0 52.431
R439 a_215_47.n3 a_215_47.n2 48.2
R440 a_215_47.n5 a_215_47.n4 33.918
R441 a_215_47.n19 a_215_47.n1 32
R442 a_215_47.n20 a_215_47.n19 32
R443 a_215_47.t2 a_215_47.n21 26.595
R444 a_215_47.n21 a_215_47.t3 26.595
R445 a_215_47.n0 a_215_47.t1 24.923
R446 a_215_47.n0 a_215_47.t4 24.923
R447 a_215_47.n17 a_215_47.n16 23.207
R448 a_215_47.n9 a_215_47.n6 21.76
R449 a_215_47.n12 a_215_47.n9 21.76
R450 a_215_47.n15 a_215_47.n12 21.76
R451 a_215_47.n18 a_215_47.n15 21.76
R452 a_215_47.n19 a_215_47.n18 21.76
R453 a_215_47.n8 a_215_47.n7 19.637
R454 a_215_47.n14 a_215_47.n13 8.925
R455 a_215_47.n11 a_215_47.n10 5.355
R456 a_109_47.n0 a_109_47.t4 221.719
R457 a_109_47.n2 a_109_47.t5 221.719
R458 a_109_47.n3 a_109_47.t7 221.719
R459 a_109_47.t0 a_109_47.n6 153.009
R460 a_109_47.n0 a_109_47.t3 149.419
R461 a_109_47.n2 a_109_47.t6 149.419
R462 a_109_47.n3 a_109_47.t2 149.419
R463 a_109_47.n6 a_109_47.t1 109.873
R464 a_109_47.n5 a_109_47.n1 97.76
R465 a_109_47.n5 a_109_47.n4 76
R466 a_109_47.n1 a_109_47.n0 51.77
R467 a_109_47.n6 a_109_47.n5 49.6
R468 a_109_47.n4 a_109_47.n2 37.488
R469 a_109_47.n4 a_109_47.n3 37.488
R470 A.n0 A.t0 230.361
R471 A.n0 A.t1 158.061
R472 A A.n0 84
C0 VGND VPWR 0.27fF
C1 X VGND 1.76fF
C2 X VPWR 2.13fF
C3 VPB VPWR 0.24fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__bufinv_8.ext - technology: sky130A

.subckt sky130_fd_sc_hd__bufinv_8 A Y VGND VPWR VNB VPB
X0 VPWR.t11 a_215_47.t6 Y.t15 VPB.t11 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 VGND.t2 a_109_47.t2 a_215_47.t4 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 VGND.t1 a_109_47.t3 a_215_47.t5 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 VGND.t11 a_215_47.t7 Y.t5 VNB.t11 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 Y.t14 a_215_47.t8 VPWR.t10 VPB.t10 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 VGND.t10 a_215_47.t9 Y.t4 VNB.t10 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 Y.t11 a_215_47.t10 VGND.t9 VNB.t9 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 Y.t10 a_215_47.t11 VGND.t8 VNB.t8 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 Y.t9 a_215_47.t12 VGND.t7 VNB.t7 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 Y.t8 a_215_47.t13 VGND.t6 VNB.t6 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 VPWR.t9 a_215_47.t14 Y.t13 VPB.t9 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 Y.t12 a_215_47.t15 VPWR.t8 VPB.t8 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 VGND.t5 a_215_47.t16 Y.t7 VNB.t5 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 VGND.t4 a_215_47.t17 Y.t6 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14 VPWR.t0 a_109_47.t4 a_215_47.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 a_215_47.t1 a_109_47.t5 VPWR.t1 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16 VPWR.t7 a_215_47.t18 Y.t3 VPB.t7 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17 a_215_47.t2 a_109_47.t6 VGND.t0 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X18 VPWR.t2 a_109_47.t7 a_215_47.t3 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X19 Y.t2 a_215_47.t19 VPWR.t6 VPB.t6 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X20 VPWR.t5 a_215_47.t20 Y.t1 VPB.t5 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X21 a_109_47.t0 A.t0 VPWR.t3 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X22 Y.t0 a_215_47.t21 VPWR.t4 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X23 a_109_47.t1 A.t1 VGND.t3 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
R0 a_215_47.n2 a_215_47.t18 221.719
R1 a_215_47.n4 a_215_47.t19 221.719
R2 a_215_47.n7 a_215_47.t20 221.719
R3 a_215_47.n12 a_215_47.t21 221.719
R4 a_215_47.n15 a_215_47.t6 221.719
R5 a_215_47.n18 a_215_47.t8 221.719
R6 a_215_47.n21 a_215_47.t14 221.719
R7 a_215_47.n24 a_215_47.t15 221.719
R8 a_215_47.n28 a_215_47.t3 173.405
R9 a_215_47.n2 a_215_47.t16 149.419
R10 a_215_47.n4 a_215_47.t11 149.419
R11 a_215_47.n7 a_215_47.t17 149.419
R12 a_215_47.n12 a_215_47.t13 149.419
R13 a_215_47.n15 a_215_47.t9 149.419
R14 a_215_47.n18 a_215_47.t12 149.419
R15 a_215_47.n21 a_215_47.t7 149.419
R16 a_215_47.n24 a_215_47.t10 149.419
R17 a_215_47.n1 a_215_47.t4 130.27
R18 a_215_47.n29 a_215_47.n28 108.41
R19 a_215_47.n6 a_215_47.n3 97.76
R20 a_215_47.n26 a_215_47.n25 76
R21 a_215_47.n6 a_215_47.n5 76
R22 a_215_47.n9 a_215_47.n8 76
R23 a_215_47.n11 a_215_47.n10 76
R24 a_215_47.n14 a_215_47.n13 76
R25 a_215_47.n17 a_215_47.n16 76
R26 a_215_47.n20 a_215_47.n19 76
R27 a_215_47.n23 a_215_47.n22 76
R28 a_215_47.n1 a_215_47.n0 52.431
R29 a_215_47.n13 a_215_47.n12 33.918
R30 a_215_47.n27 a_215_47.n1 32
R31 a_215_47.n28 a_215_47.n27 32
R32 a_215_47.t0 a_215_47.n29 26.595
R33 a_215_47.n29 a_215_47.t1 26.595
R34 a_215_47.n0 a_215_47.t5 24.923
R35 a_215_47.n0 a_215_47.t2 24.923
R36 a_215_47.n25 a_215_47.n24 23.207
R37 a_215_47.n9 a_215_47.n6 21.76
R38 a_215_47.n11 a_215_47.n9 21.76
R39 a_215_47.n14 a_215_47.n11 21.76
R40 a_215_47.n17 a_215_47.n14 21.76
R41 a_215_47.n20 a_215_47.n17 21.76
R42 a_215_47.n23 a_215_47.n20 21.76
R43 a_215_47.n26 a_215_47.n23 21.76
R44 a_215_47.n27 a_215_47.n26 21.76
R45 a_215_47.n16 a_215_47.n15 19.637
R46 a_215_47.n3 a_215_47.n2 16.066
R47 a_215_47.n8 a_215_47.n7 12.496
R48 a_215_47.n22 a_215_47.n21 8.925
R49 a_215_47.n19 a_215_47.n18 5.355
R50 a_215_47.n5 a_215_47.n4 1.785
R51 Y.n2 Y.n0 146.81
R52 Y.n2 Y.n1 108.41
R53 Y.n4 Y.n3 108.41
R54 Y.n6 Y.n5 108.41
R55 Y.n9 Y.n7 90.831
R56 Y.n9 Y.n8 52.431
R57 Y.n11 Y.n10 52.431
R58 Y.n13 Y.n12 52.431
R59 Y Y.n13 39.969
R60 Y.n11 Y.n9 38.4
R61 Y.n13 Y.n11 38.4
R62 Y.n4 Y.n2 38.4
R63 Y.n6 Y.n4 38.4
R64 Y Y.n6 33.319
R65 Y.n0 Y.t13 26.595
R66 Y.n0 Y.t12 26.595
R67 Y.n1 Y.t15 26.595
R68 Y.n1 Y.t14 26.595
R69 Y.n3 Y.t1 26.595
R70 Y.n3 Y.t0 26.595
R71 Y.n5 Y.t3 26.595
R72 Y.n5 Y.t2 26.595
R73 Y.n7 Y.t5 24.923
R74 Y.n7 Y.t11 24.923
R75 Y.n8 Y.t4 24.923
R76 Y.n8 Y.t9 24.923
R77 Y.n10 Y.t6 24.923
R78 Y.n10 Y.t8 24.923
R79 Y.n12 Y.t7 24.923
R80 Y.n12 Y.t10 24.923
R81 VPWR.n0 VPWR.t7 208.281
R82 VPWR.n24 VPWR.n23 174.594
R83 VPWR.n18 VPWR.n17 174.594
R84 VPWR.n12 VPWR.n11 174.594
R85 VPWR.n8 VPWR.n7 174.594
R86 VPWR.n2 VPWR.n1 174.594
R87 VPWR.n31 VPWR.t3 159.459
R88 VPWR.n23 VPWR.t1 26.595
R89 VPWR.n23 VPWR.t2 26.595
R90 VPWR.n17 VPWR.t8 26.595
R91 VPWR.n17 VPWR.t0 26.595
R92 VPWR.n11 VPWR.t10 26.595
R93 VPWR.n11 VPWR.t9 26.595
R94 VPWR.n7 VPWR.t4 26.595
R95 VPWR.n7 VPWR.t11 26.595
R96 VPWR.n1 VPWR.t6 26.595
R97 VPWR.n1 VPWR.t5 26.595
R98 VPWR.n9 VPWR.n8 17.317
R99 VPWR.n3 VPWR.n2 11.294
R100 VPWR.n13 VPWR.n12 11.294
R101 VPWR.n32 VPWR.n31 6.908
R102 VPWR.n19 VPWR.n18 5.27
R103 VPWR.n4 VPWR.n3 4.65
R104 VPWR.n6 VPWR.n5 4.65
R105 VPWR.n10 VPWR.n9 4.65
R106 VPWR.n14 VPWR.n13 4.65
R107 VPWR.n16 VPWR.n15 4.65
R108 VPWR.n20 VPWR.n19 4.65
R109 VPWR.n22 VPWR.n21 4.65
R110 VPWR.n26 VPWR.n25 4.65
R111 VPWR.n28 VPWR.n27 4.65
R112 VPWR.n30 VPWR.n29 4.65
R113 VPWR.n25 VPWR.n24 0.752
R114 VPWR.n4 VPWR.n0 0.517
R115 VPWR.n6 VPWR.n4 0.119
R116 VPWR.n10 VPWR.n6 0.119
R117 VPWR.n14 VPWR.n10 0.119
R118 VPWR.n16 VPWR.n14 0.119
R119 VPWR.n20 VPWR.n16 0.119
R120 VPWR.n22 VPWR.n20 0.119
R121 VPWR.n26 VPWR.n22 0.119
R122 VPWR.n28 VPWR.n26 0.119
R123 VPWR.n30 VPWR.n28 0.119
R124 VPWR.n32 VPWR.n30 0.119
R125 VPWR VPWR.n32 0.02
R126 VPB.t3 VPB.t2 556.386
R127 VPB.t6 VPB.t7 248.598
R128 VPB.t5 VPB.t6 248.598
R129 VPB.t4 VPB.t5 248.598
R130 VPB.t11 VPB.t4 248.598
R131 VPB.t10 VPB.t11 248.598
R132 VPB.t9 VPB.t10 248.598
R133 VPB.t8 VPB.t9 248.598
R134 VPB.t0 VPB.t8 248.598
R135 VPB.t1 VPB.t0 248.598
R136 VPB.t2 VPB.t1 248.598
R137 VPB VPB.t3 189.408
R138 a_109_47.n0 a_109_47.t4 221.719
R139 a_109_47.n2 a_109_47.t5 221.719
R140 a_109_47.n3 a_109_47.t7 221.719
R141 a_109_47.t0 a_109_47.n6 154.753
R142 a_109_47.n0 a_109_47.t3 149.419
R143 a_109_47.n2 a_109_47.t6 149.419
R144 a_109_47.n3 a_109_47.t2 149.419
R145 a_109_47.n6 a_109_47.t1 107.967
R146 a_109_47.n5 a_109_47.n1 97.76
R147 a_109_47.n5 a_109_47.n4 76
R148 a_109_47.n6 a_109_47.n5 55.04
R149 a_109_47.n1 a_109_47.n0 51.77
R150 a_109_47.n4 a_109_47.n2 37.488
R151 a_109_47.n4 a_109_47.n3 37.488
R152 VGND.n0 VGND.t5 197.155
R153 VGND.n2 VGND.n1 116.217
R154 VGND.n8 VGND.n7 116.217
R155 VGND.n12 VGND.n11 116.217
R156 VGND.n18 VGND.n17 116.217
R157 VGND.n24 VGND.n23 116.217
R158 VGND.n31 VGND.t3 114.773
R159 VGND.n1 VGND.t8 24.923
R160 VGND.n1 VGND.t4 24.923
R161 VGND.n7 VGND.t6 24.923
R162 VGND.n7 VGND.t10 24.923
R163 VGND.n11 VGND.t7 24.923
R164 VGND.n11 VGND.t11 24.923
R165 VGND.n17 VGND.t9 24.923
R166 VGND.n17 VGND.t1 24.923
R167 VGND.n23 VGND.t0 24.923
R168 VGND.n23 VGND.t2 24.923
R169 VGND.n9 VGND.n8 17.317
R170 VGND.n3 VGND.n2 11.294
R171 VGND.n13 VGND.n12 11.294
R172 VGND.n32 VGND.n31 6.908
R173 VGND.n19 VGND.n18 5.27
R174 VGND.n4 VGND.n3 4.65
R175 VGND.n6 VGND.n5 4.65
R176 VGND.n10 VGND.n9 4.65
R177 VGND.n14 VGND.n13 4.65
R178 VGND.n16 VGND.n15 4.65
R179 VGND.n20 VGND.n19 4.65
R180 VGND.n22 VGND.n21 4.65
R181 VGND.n26 VGND.n25 4.65
R182 VGND.n28 VGND.n27 4.65
R183 VGND.n30 VGND.n29 4.65
R184 VGND.n25 VGND.n24 0.752
R185 VGND.n4 VGND.n0 0.517
R186 VGND.n6 VGND.n4 0.119
R187 VGND.n10 VGND.n6 0.119
R188 VGND.n14 VGND.n10 0.119
R189 VGND.n16 VGND.n14 0.119
R190 VGND.n20 VGND.n16 0.119
R191 VGND.n22 VGND.n20 0.119
R192 VGND.n26 VGND.n22 0.119
R193 VGND.n28 VGND.n26 0.119
R194 VGND.n30 VGND.n28 0.119
R195 VGND.n32 VGND.n30 0.119
R196 VGND VGND.n32 0.02
R197 VNB VNB.t3 6053.91
R198 VNB.t3 VNB.t2 4545.05
R199 VNB.t8 VNB.t5 2030.77
R200 VNB.t4 VNB.t8 2030.77
R201 VNB.t6 VNB.t4 2030.77
R202 VNB.t10 VNB.t6 2030.77
R203 VNB.t7 VNB.t10 2030.77
R204 VNB.t11 VNB.t7 2030.77
R205 VNB.t9 VNB.t11 2030.77
R206 VNB.t1 VNB.t9 2030.77
R207 VNB.t0 VNB.t1 2030.77
R208 VNB.t2 VNB.t0 2030.77
R209 A.n0 A.t0 230.154
R210 A.n0 A.t1 157.854
R211 A A.n0 84
C0 VGND Y 0.89fF
C1 VGND VPWR 0.14fF
C2 VPWR Y 1.08fF
C3 VPB VPWR 0.14fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__bufinv_16.ext - technology: sky130A

.subckt sky130_fd_sc_hd__bufinv_16 A Y VGND VPWR VNB VPB
X0 a_361_47.t5 a_27_47.t6 VGND.t15 VNB.t7 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 VPWR.t24 a_361_47.t12 Y.t24 VPB.t24 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 a_361_47.t4 a_27_47.t7 VGND.t14 VNB.t6 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 Y.t15 a_361_47.t13 VGND.t19 VNB.t23 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 VPWR.t23 a_361_47.t14 Y.t23 VPB.t23 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 Y.t14 a_361_47.t15 VGND.t1 VNB.t22 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 Y.t22 a_361_47.t16 VPWR.t22 VPB.t22 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 VPWR.t8 a_27_47.t8 a_361_47.t11 VPB.t8 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 VPWR.t21 a_361_47.t17 Y.t21 VPB.t21 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 VPWR.t20 a_361_47.t18 Y.t20 VPB.t20 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 VGND.t2 a_361_47.t19 Y.t13 VNB.t21 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 a_361_47.t10 a_27_47.t9 VPWR.t7 VPB.t7 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 VGND.t3 a_361_47.t20 Y.t12 VNB.t20 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 VGND.t4 a_361_47.t21 Y.t11 VNB.t19 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14 VGND.t16 a_361_47.t22 Y.t10 VNB.t18 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X15 VGND.t17 a_361_47.t23 Y.t9 VNB.t17 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X16 VPWR.t2 A.t0 a_27_47.t4 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17 Y.t19 a_361_47.t24 VPWR.t19 VPB.t19 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X18 VGND.t18 a_361_47.t25 Y.t8 VNB.t16 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X19 VPWR.t18 a_361_47.t26 Y.t18 VPB.t18 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X20 a_27_47.t0 A.t1 VPWR.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X21 Y.t31 a_361_47.t27 VPWR.t17 VPB.t17 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X22 a_27_47.t1 A.t2 VGND.t5 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X23 a_361_47.t3 a_27_47.t10 VGND.t13 VNB.t5 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X24 Y.t30 a_361_47.t28 VPWR.t16 VPB.t16 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X25 Y.t7 a_361_47.t29 VGND.t20 VNB.t15 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X26 VPWR.t6 a_27_47.t11 a_361_47.t9 VPB.t6 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X27 Y.t6 a_361_47.t30 VGND.t21 VNB.t14 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X28 Y.t29 a_361_47.t31 VPWR.t15 VPB.t15 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X29 Y.t5 a_361_47.t32 VGND.t22 VNB.t13 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X30 a_361_47.t8 a_27_47.t12 VPWR.t5 VPB.t5 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X31 VPWR.t14 a_361_47.t33 Y.t28 VPB.t14 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X32 Y.t4 a_361_47.t34 VGND.t23 VNB.t12 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X33 VGND.t6 A.t3 a_27_47.t2 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X34 VGND.t12 a_27_47.t13 a_361_47.t2 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X35 VPWR.t4 a_27_47.t14 a_361_47.t7 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X36 Y.t27 a_361_47.t35 VPWR.t13 VPB.t13 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X37 VGND.t11 a_27_47.t15 a_361_47.t1 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X38 VGND.t10 a_27_47.t16 a_361_47.t0 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X39 a_361_47.t6 a_27_47.t17 VPWR.t3 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X40 VPWR.t12 a_361_47.t36 Y.t26 VPB.t12 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X41 VPWR.t11 a_361_47.t37 Y.t25 VPB.t11 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X42 VGND.t7 a_361_47.t38 Y.t3 VNB.t11 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X43 VGND.t8 a_361_47.t39 Y.t2 VNB.t10 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X44 VPWR.t1 A.t4 a_27_47.t3 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X45 Y.t17 a_361_47.t40 VPWR.t10 VPB.t10 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X46 Y.t1 a_361_47.t41 VGND.t9 VNB.t9 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X47 Y.t16 a_361_47.t42 VPWR.t9 VPB.t9 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X48 VGND.t24 A.t5 a_27_47.t5 VNB.t24 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X49 Y.t0 a_361_47.t43 VGND.t0 VNB.t8 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
R0 a_27_47.n2 a_27_47.t11 221.719
R1 a_27_47.n4 a_27_47.t12 221.719
R2 a_27_47.n7 a_27_47.t14 221.719
R3 a_27_47.n10 a_27_47.t17 221.719
R4 a_27_47.n13 a_27_47.t8 221.719
R5 a_27_47.n16 a_27_47.t9 221.719
R6 a_27_47.n20 a_27_47.t3 173.405
R7 a_27_47.n2 a_27_47.t16 149.419
R8 a_27_47.n4 a_27_47.t7 149.419
R9 a_27_47.n7 a_27_47.t15 149.419
R10 a_27_47.n10 a_27_47.t6 149.419
R11 a_27_47.n13 a_27_47.t13 149.419
R12 a_27_47.n16 a_27_47.t10 149.419
R13 a_27_47.n1 a_27_47.t5 130.27
R14 a_27_47.n21 a_27_47.n20 108.41
R15 a_27_47.n6 a_27_47.n3 97.76
R16 a_27_47.n18 a_27_47.n17 76
R17 a_27_47.n6 a_27_47.n5 76
R18 a_27_47.n9 a_27_47.n8 76
R19 a_27_47.n12 a_27_47.n11 76
R20 a_27_47.n15 a_27_47.n14 76
R21 a_27_47.n1 a_27_47.n0 52.431
R22 a_27_47.n3 a_27_47.n2 48.2
R23 a_27_47.n5 a_27_47.n4 33.918
R24 a_27_47.n19 a_27_47.n1 32
R25 a_27_47.n20 a_27_47.n19 32
R26 a_27_47.n21 a_27_47.t4 26.595
R27 a_27_47.t0 a_27_47.n21 26.595
R28 a_27_47.n0 a_27_47.t2 24.923
R29 a_27_47.n0 a_27_47.t1 24.923
R30 a_27_47.n17 a_27_47.n16 23.207
R31 a_27_47.n9 a_27_47.n6 21.76
R32 a_27_47.n12 a_27_47.n9 21.76
R33 a_27_47.n15 a_27_47.n12 21.76
R34 a_27_47.n18 a_27_47.n15 21.76
R35 a_27_47.n19 a_27_47.n18 21.76
R36 a_27_47.n8 a_27_47.n7 19.637
R37 a_27_47.n14 a_27_47.n13 8.925
R38 a_27_47.n11 a_27_47.n10 5.355
R39 VGND.n0 VGND.t2 196.044
R40 VGND.n2 VGND.n1 116.217
R41 VGND.n8 VGND.n7 116.217
R42 VGND.n14 VGND.n13 116.217
R43 VGND.n18 VGND.n17 116.217
R44 VGND.n24 VGND.n23 116.217
R45 VGND.n30 VGND.n29 116.217
R46 VGND.n36 VGND.n35 116.217
R47 VGND.n42 VGND.n41 116.217
R48 VGND.n48 VGND.n47 116.217
R49 VGND.n52 VGND.n51 116.217
R50 VGND.n58 VGND.n57 116.217
R51 VGND.n64 VGND.n63 116.217
R52 VGND.n1 VGND.t9 24.923
R53 VGND.n1 VGND.t8 24.923
R54 VGND.n7 VGND.t23 24.923
R55 VGND.n7 VGND.t7 24.923
R56 VGND.n13 VGND.t22 24.923
R57 VGND.n13 VGND.t18 24.923
R58 VGND.n17 VGND.t21 24.923
R59 VGND.n17 VGND.t17 24.923
R60 VGND.n23 VGND.t20 24.923
R61 VGND.n23 VGND.t4 24.923
R62 VGND.n29 VGND.t19 24.923
R63 VGND.n29 VGND.t3 24.923
R64 VGND.n35 VGND.t0 24.923
R65 VGND.n35 VGND.t16 24.923
R66 VGND.n41 VGND.t1 24.923
R67 VGND.n41 VGND.t10 24.923
R68 VGND.n47 VGND.t14 24.923
R69 VGND.n47 VGND.t11 24.923
R70 VGND.n51 VGND.t15 24.923
R71 VGND.n51 VGND.t12 24.923
R72 VGND.n57 VGND.t13 24.923
R73 VGND.n57 VGND.t6 24.923
R74 VGND.n63 VGND.t5 24.923
R75 VGND.n63 VGND.t24 24.923
R76 VGND.n49 VGND.n48 15.811
R77 VGND.n15 VGND.n14 14.305
R78 VGND.n19 VGND.n18 14.305
R79 VGND.n53 VGND.n52 12.8
R80 VGND.n43 VGND.n42 9.788
R81 VGND.n9 VGND.n8 8.282
R82 VGND.n25 VGND.n24 8.282
R83 VGND.n59 VGND.n58 6.776
R84 VGND.n4 VGND.n3 4.65
R85 VGND.n6 VGND.n5 4.65
R86 VGND.n10 VGND.n9 4.65
R87 VGND.n12 VGND.n11 4.65
R88 VGND.n16 VGND.n15 4.65
R89 VGND.n20 VGND.n19 4.65
R90 VGND.n22 VGND.n21 4.65
R91 VGND.n26 VGND.n25 4.65
R92 VGND.n28 VGND.n27 4.65
R93 VGND.n32 VGND.n31 4.65
R94 VGND.n34 VGND.n33 4.65
R95 VGND.n38 VGND.n37 4.65
R96 VGND.n40 VGND.n39 4.65
R97 VGND.n44 VGND.n43 4.65
R98 VGND.n46 VGND.n45 4.65
R99 VGND.n50 VGND.n49 4.65
R100 VGND.n54 VGND.n53 4.65
R101 VGND.n56 VGND.n55 4.65
R102 VGND.n60 VGND.n59 4.65
R103 VGND.n62 VGND.n61 4.65
R104 VGND.n66 VGND.n65 4.65
R105 VGND.n37 VGND.n36 3.764
R106 VGND.n3 VGND.n2 2.258
R107 VGND.n31 VGND.n30 2.258
R108 VGND.n4 VGND.n0 1.02
R109 VGND.n65 VGND.n64 0.752
R110 VGND.n6 VGND.n4 0.119
R111 VGND.n10 VGND.n6 0.119
R112 VGND.n12 VGND.n10 0.119
R113 VGND.n16 VGND.n12 0.119
R114 VGND.n20 VGND.n16 0.119
R115 VGND.n22 VGND.n20 0.119
R116 VGND.n26 VGND.n22 0.119
R117 VGND.n28 VGND.n26 0.119
R118 VGND.n32 VGND.n28 0.119
R119 VGND.n34 VGND.n32 0.119
R120 VGND.n38 VGND.n34 0.119
R121 VGND.n40 VGND.n38 0.119
R122 VGND.n44 VGND.n40 0.119
R123 VGND.n46 VGND.n44 0.119
R124 VGND.n50 VGND.n46 0.119
R125 VGND.n54 VGND.n50 0.119
R126 VGND.n56 VGND.n54 0.119
R127 VGND.n60 VGND.n56 0.119
R128 VGND.n62 VGND.n60 0.119
R129 VGND.n66 VGND.n62 0.119
R130 VGND.n67 VGND.n66 0.119
R131 VGND VGND.n67 0.02
R132 a_361_47.n6 a_361_47.t17 221.719
R133 a_361_47.n7 a_361_47.t28 221.719
R134 a_361_47.n9 a_361_47.t37 221.719
R135 a_361_47.n14 a_361_47.t42 221.719
R136 a_361_47.n17 a_361_47.t14 221.719
R137 a_361_47.n20 a_361_47.t16 221.719
R138 a_361_47.n23 a_361_47.t18 221.719
R139 a_361_47.n28 a_361_47.t31 221.719
R140 a_361_47.n31 a_361_47.t33 221.719
R141 a_361_47.n34 a_361_47.t35 221.719
R142 a_361_47.n37 a_361_47.t36 221.719
R143 a_361_47.n42 a_361_47.t40 221.719
R144 a_361_47.n45 a_361_47.t12 221.719
R145 a_361_47.n48 a_361_47.t24 221.719
R146 a_361_47.n51 a_361_47.t26 221.719
R147 a_361_47.n54 a_361_47.t27 221.719
R148 a_361_47.n6 a_361_47.t19 149.419
R149 a_361_47.n7 a_361_47.t41 149.419
R150 a_361_47.n9 a_361_47.t39 149.419
R151 a_361_47.n14 a_361_47.t34 149.419
R152 a_361_47.n17 a_361_47.t38 149.419
R153 a_361_47.n20 a_361_47.t32 149.419
R154 a_361_47.n23 a_361_47.t25 149.419
R155 a_361_47.n28 a_361_47.t30 149.419
R156 a_361_47.n31 a_361_47.t23 149.419
R157 a_361_47.n34 a_361_47.t29 149.419
R158 a_361_47.n37 a_361_47.t21 149.419
R159 a_361_47.n42 a_361_47.t13 149.419
R160 a_361_47.n45 a_361_47.t20 149.419
R161 a_361_47.n48 a_361_47.t43 149.419
R162 a_361_47.n51 a_361_47.t22 149.419
R163 a_361_47.n54 a_361_47.t15 149.419
R164 a_361_47.n3 a_361_47.n1 146.81
R165 a_361_47.n3 a_361_47.n2 108.41
R166 a_361_47.n5 a_361_47.n4 108.41
R167 a_361_47.n11 a_361_47.n8 97.76
R168 a_361_47.n60 a_361_47.n0 90.831
R169 a_361_47.n56 a_361_47.n55 76
R170 a_361_47.n11 a_361_47.n10 76
R171 a_361_47.n13 a_361_47.n12 76
R172 a_361_47.n16 a_361_47.n15 76
R173 a_361_47.n19 a_361_47.n18 76
R174 a_361_47.n22 a_361_47.n21 76
R175 a_361_47.n25 a_361_47.n24 76
R176 a_361_47.n27 a_361_47.n26 76
R177 a_361_47.n30 a_361_47.n29 76
R178 a_361_47.n33 a_361_47.n32 76
R179 a_361_47.n36 a_361_47.n35 76
R180 a_361_47.n39 a_361_47.n38 76
R181 a_361_47.n41 a_361_47.n40 76
R182 a_361_47.n44 a_361_47.n43 76
R183 a_361_47.n47 a_361_47.n46 76
R184 a_361_47.n50 a_361_47.n49 76
R185 a_361_47.n53 a_361_47.n52 76
R186 a_361_47.n8 a_361_47.n6 73.192
R187 a_361_47.n59 a_361_47.n58 52.431
R188 a_361_47.n61 a_361_47.n60 52.431
R189 a_361_47.n5 a_361_47.n3 38.4
R190 a_361_47.n60 a_361_47.n59 38.4
R191 a_361_47.n43 a_361_47.n42 37.488
R192 a_361_47.n29 a_361_47.n28 33.918
R193 a_361_47.n57 a_361_47.n5 31.074
R194 a_361_47.n59 a_361_47.n57 31.074
R195 a_361_47.n15 a_361_47.n14 30.348
R196 a_361_47.n1 a_361_47.t11 26.595
R197 a_361_47.n1 a_361_47.t10 26.595
R198 a_361_47.n2 a_361_47.t7 26.595
R199 a_361_47.n2 a_361_47.t6 26.595
R200 a_361_47.n4 a_361_47.t9 26.595
R201 a_361_47.n4 a_361_47.t8 26.595
R202 a_361_47.n58 a_361_47.t0 24.923
R203 a_361_47.n58 a_361_47.t4 24.923
R204 a_361_47.n0 a_361_47.t2 24.923
R205 a_361_47.n0 a_361_47.t3 24.923
R206 a_361_47.n61 a_361_47.t1 24.923
R207 a_361_47.t5 a_361_47.n61 24.923
R208 a_361_47.n46 a_361_47.n45 23.207
R209 a_361_47.n13 a_361_47.n11 21.76
R210 a_361_47.n16 a_361_47.n13 21.76
R211 a_361_47.n19 a_361_47.n16 21.76
R212 a_361_47.n22 a_361_47.n19 21.76
R213 a_361_47.n25 a_361_47.n22 21.76
R214 a_361_47.n27 a_361_47.n25 21.76
R215 a_361_47.n30 a_361_47.n27 21.76
R216 a_361_47.n33 a_361_47.n30 21.76
R217 a_361_47.n36 a_361_47.n33 21.76
R218 a_361_47.n39 a_361_47.n36 21.76
R219 a_361_47.n41 a_361_47.n39 21.76
R220 a_361_47.n44 a_361_47.n41 21.76
R221 a_361_47.n47 a_361_47.n44 21.76
R222 a_361_47.n50 a_361_47.n47 21.76
R223 a_361_47.n53 a_361_47.n50 21.76
R224 a_361_47.n56 a_361_47.n53 21.76
R225 a_361_47.n57 a_361_47.n56 20.8
R226 a_361_47.n32 a_361_47.n31 19.637
R227 a_361_47.n55 a_361_47.n54 19.637
R228 a_361_47.n10 a_361_47.n9 16.066
R229 a_361_47.n18 a_361_47.n17 16.066
R230 a_361_47.n24 a_361_47.n23 12.496
R231 a_361_47.n38 a_361_47.n37 8.925
R232 a_361_47.n49 a_361_47.n48 8.925
R233 a_361_47.n35 a_361_47.n34 5.355
R234 a_361_47.n52 a_361_47.n51 5.355
R235 a_361_47.n8 a_361_47.n7 1.785
R236 a_361_47.n21 a_361_47.n20 1.785
R237 VNB VNB.t24 6053.91
R238 VNB.t9 VNB.t21 2030.77
R239 VNB.t10 VNB.t9 2030.77
R240 VNB.t12 VNB.t10 2030.77
R241 VNB.t11 VNB.t12 2030.77
R242 VNB.t13 VNB.t11 2030.77
R243 VNB.t16 VNB.t13 2030.77
R244 VNB.t14 VNB.t16 2030.77
R245 VNB.t17 VNB.t14 2030.77
R246 VNB.t15 VNB.t17 2030.77
R247 VNB.t19 VNB.t15 2030.77
R248 VNB.t23 VNB.t19 2030.77
R249 VNB.t20 VNB.t23 2030.77
R250 VNB.t8 VNB.t20 2030.77
R251 VNB.t18 VNB.t8 2030.77
R252 VNB.t22 VNB.t18 2030.77
R253 VNB.t2 VNB.t22 2030.77
R254 VNB.t6 VNB.t2 2030.77
R255 VNB.t3 VNB.t6 2030.77
R256 VNB.t7 VNB.t3 2030.77
R257 VNB.t4 VNB.t7 2030.77
R258 VNB.t5 VNB.t4 2030.77
R259 VNB.t1 VNB.t5 2030.77
R260 VNB.t0 VNB.t1 2030.77
R261 VNB.t24 VNB.t0 2030.77
R262 Y.n2 Y.n0 146.81
R263 Y.n2 Y.n1 108.41
R264 Y.n4 Y.n3 108.41
R265 Y.n6 Y.n5 108.41
R266 Y.n8 Y.n7 108.41
R267 Y.n10 Y.n9 108.41
R268 Y.n12 Y.n11 108.41
R269 Y.n14 Y.n13 108.41
R270 Y.n17 Y.n15 90.831
R271 Y.n17 Y.n16 52.431
R272 Y.n19 Y.n18 52.431
R273 Y.n21 Y.n20 52.431
R274 Y.n23 Y.n22 52.431
R275 Y.n25 Y.n24 52.431
R276 Y.n27 Y.n26 52.431
R277 Y.n29 Y.n28 52.431
R278 Y.n19 Y.n17 38.4
R279 Y.n21 Y.n19 38.4
R280 Y.n23 Y.n21 38.4
R281 Y.n25 Y.n23 38.4
R282 Y.n27 Y.n25 38.4
R283 Y.n29 Y.n27 38.4
R284 Y.n4 Y.n2 38.4
R285 Y.n6 Y.n4 38.4
R286 Y.n8 Y.n6 38.4
R287 Y.n10 Y.n8 38.4
R288 Y.n12 Y.n10 38.4
R289 Y.n14 Y.n12 38.4
R290 Y.n0 Y.t18 26.595
R291 Y.n0 Y.t31 26.595
R292 Y.n1 Y.t24 26.595
R293 Y.n1 Y.t19 26.595
R294 Y.n3 Y.t26 26.595
R295 Y.n3 Y.t17 26.595
R296 Y.n5 Y.t28 26.595
R297 Y.n5 Y.t27 26.595
R298 Y.n7 Y.t20 26.595
R299 Y.n7 Y.t29 26.595
R300 Y.n9 Y.t23 26.595
R301 Y.n9 Y.t22 26.595
R302 Y.n11 Y.t25 26.595
R303 Y.n11 Y.t16 26.595
R304 Y.n13 Y.t21 26.595
R305 Y.n13 Y.t30 26.595
R306 Y Y.n29 26.441
R307 Y.n15 Y.t10 24.923
R308 Y.n15 Y.t14 24.923
R309 Y.n16 Y.t12 24.923
R310 Y.n16 Y.t0 24.923
R311 Y.n18 Y.t11 24.923
R312 Y.n18 Y.t15 24.923
R313 Y.n20 Y.t9 24.923
R314 Y.n20 Y.t7 24.923
R315 Y.n22 Y.t8 24.923
R316 Y.n22 Y.t6 24.923
R317 Y.n24 Y.t3 24.923
R318 Y.n24 Y.t5 24.923
R319 Y.n26 Y.t2 24.923
R320 Y.n26 Y.t4 24.923
R321 Y.n28 Y.t13 24.923
R322 Y.n28 Y.t1 24.923
R323 Y Y.n14 17.132
R324 VPWR.n0 VPWR.t21 207.169
R325 VPWR.n64 VPWR.n63 174.594
R326 VPWR.n58 VPWR.n57 174.594
R327 VPWR.n52 VPWR.n51 174.594
R328 VPWR.n48 VPWR.n47 174.594
R329 VPWR.n42 VPWR.n41 174.594
R330 VPWR.n36 VPWR.n35 174.594
R331 VPWR.n30 VPWR.n29 174.594
R332 VPWR.n24 VPWR.n23 174.594
R333 VPWR.n18 VPWR.n17 174.594
R334 VPWR.n14 VPWR.n13 174.594
R335 VPWR.n8 VPWR.n7 174.594
R336 VPWR.n2 VPWR.n1 174.594
R337 VPWR.n63 VPWR.t0 26.595
R338 VPWR.n63 VPWR.t1 26.595
R339 VPWR.n57 VPWR.t7 26.595
R340 VPWR.n57 VPWR.t2 26.595
R341 VPWR.n51 VPWR.t3 26.595
R342 VPWR.n51 VPWR.t8 26.595
R343 VPWR.n47 VPWR.t5 26.595
R344 VPWR.n47 VPWR.t4 26.595
R345 VPWR.n41 VPWR.t17 26.595
R346 VPWR.n41 VPWR.t6 26.595
R347 VPWR.n35 VPWR.t19 26.595
R348 VPWR.n35 VPWR.t18 26.595
R349 VPWR.n29 VPWR.t10 26.595
R350 VPWR.n29 VPWR.t24 26.595
R351 VPWR.n23 VPWR.t13 26.595
R352 VPWR.n23 VPWR.t12 26.595
R353 VPWR.n17 VPWR.t15 26.595
R354 VPWR.n17 VPWR.t14 26.595
R355 VPWR.n13 VPWR.t22 26.595
R356 VPWR.n13 VPWR.t20 26.595
R357 VPWR.n7 VPWR.t9 26.595
R358 VPWR.n7 VPWR.t23 26.595
R359 VPWR.n1 VPWR.t16 26.595
R360 VPWR.n1 VPWR.t11 26.595
R361 VPWR.n49 VPWR.n48 15.811
R362 VPWR.n15 VPWR.n14 14.305
R363 VPWR.n19 VPWR.n18 14.305
R364 VPWR.n53 VPWR.n52 12.8
R365 VPWR.n43 VPWR.n42 9.788
R366 VPWR.n9 VPWR.n8 8.282
R367 VPWR.n25 VPWR.n24 8.282
R368 VPWR.n59 VPWR.n58 6.776
R369 VPWR.n66 VPWR.n65 4.65
R370 VPWR.n4 VPWR.n3 4.65
R371 VPWR.n6 VPWR.n5 4.65
R372 VPWR.n10 VPWR.n9 4.65
R373 VPWR.n12 VPWR.n11 4.65
R374 VPWR.n16 VPWR.n15 4.65
R375 VPWR.n20 VPWR.n19 4.65
R376 VPWR.n22 VPWR.n21 4.65
R377 VPWR.n26 VPWR.n25 4.65
R378 VPWR.n28 VPWR.n27 4.65
R379 VPWR.n32 VPWR.n31 4.65
R380 VPWR.n34 VPWR.n33 4.65
R381 VPWR.n38 VPWR.n37 4.65
R382 VPWR.n40 VPWR.n39 4.65
R383 VPWR.n44 VPWR.n43 4.65
R384 VPWR.n46 VPWR.n45 4.65
R385 VPWR.n50 VPWR.n49 4.65
R386 VPWR.n54 VPWR.n53 4.65
R387 VPWR.n56 VPWR.n55 4.65
R388 VPWR.n60 VPWR.n59 4.65
R389 VPWR.n62 VPWR.n61 4.65
R390 VPWR.n37 VPWR.n36 3.764
R391 VPWR.n3 VPWR.n2 2.258
R392 VPWR.n31 VPWR.n30 2.258
R393 VPWR.n4 VPWR.n0 1.02
R394 VPWR.n65 VPWR.n64 0.752
R395 VPWR.n6 VPWR.n4 0.119
R396 VPWR.n10 VPWR.n6 0.119
R397 VPWR.n12 VPWR.n10 0.119
R398 VPWR.n16 VPWR.n12 0.119
R399 VPWR.n20 VPWR.n16 0.119
R400 VPWR.n22 VPWR.n20 0.119
R401 VPWR.n26 VPWR.n22 0.119
R402 VPWR.n28 VPWR.n26 0.119
R403 VPWR.n32 VPWR.n28 0.119
R404 VPWR.n34 VPWR.n32 0.119
R405 VPWR.n38 VPWR.n34 0.119
R406 VPWR.n40 VPWR.n38 0.119
R407 VPWR.n44 VPWR.n40 0.119
R408 VPWR.n46 VPWR.n44 0.119
R409 VPWR.n50 VPWR.n46 0.119
R410 VPWR.n54 VPWR.n50 0.119
R411 VPWR.n56 VPWR.n54 0.119
R412 VPWR.n60 VPWR.n56 0.119
R413 VPWR.n62 VPWR.n60 0.119
R414 VPWR.n66 VPWR.n62 0.119
R415 VPWR.n67 VPWR.n66 0.119
R416 VPWR VPWR.n67 0.02
R417 VPB.t16 VPB.t21 248.598
R418 VPB.t11 VPB.t16 248.598
R419 VPB.t9 VPB.t11 248.598
R420 VPB.t23 VPB.t9 248.598
R421 VPB.t22 VPB.t23 248.598
R422 VPB.t20 VPB.t22 248.598
R423 VPB.t15 VPB.t20 248.598
R424 VPB.t14 VPB.t15 248.598
R425 VPB.t13 VPB.t14 248.598
R426 VPB.t12 VPB.t13 248.598
R427 VPB.t10 VPB.t12 248.598
R428 VPB.t24 VPB.t10 248.598
R429 VPB.t19 VPB.t24 248.598
R430 VPB.t18 VPB.t19 248.598
R431 VPB.t17 VPB.t18 248.598
R432 VPB.t6 VPB.t17 248.598
R433 VPB.t5 VPB.t6 248.598
R434 VPB.t4 VPB.t5 248.598
R435 VPB.t3 VPB.t4 248.598
R436 VPB.t8 VPB.t3 248.598
R437 VPB.t7 VPB.t8 248.598
R438 VPB.t2 VPB.t7 248.598
R439 VPB.t0 VPB.t2 248.598
R440 VPB.t1 VPB.t0 248.598
R441 VPB VPB.t1 189.408
R442 A.n0 A.t0 221.719
R443 A.n2 A.t1 221.719
R444 A.n3 A.t4 221.719
R445 A.n0 A.t3 149.419
R446 A.n2 A.t2 149.419
R447 A.n3 A.t5 149.419
R448 A.n5 A.n1 97.76
R449 A.n5 A.n4 76
R450 A.n1 A.n0 51.77
R451 A.n4 A.n2 37.488
R452 A.n4 A.n3 37.488
R453 A A.n5 33.92
C0 VPB VPWR 0.22fF
C1 VGND Y 1.76fF
C2 VGND VPWR 0.24fF
C3 VPWR Y 2.13fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__clkbuf_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__clkbuf_1 VGND VPWR X A VNB VPB
X0 VPWR.t1 a_75_212.t2 X.t0 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X1 a_75_212.t0 A.t0 VGND.t0 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X2 a_75_212.t1 A.t1 VPWR.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X3 VGND.t1 a_75_212.t3 X.t1 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
R0 a_75_212.t1 a_75_212.n1 260.844
R1 a_75_212.n0 a_75_212.t2 254.387
R2 a_75_212.n0 a_75_212.t3 211.007
R3 a_75_212.n1 a_75_212.t0 201.838
R4 a_75_212.n1 a_75_212.n0 76
R5 X.n1 X.t0 222.242
R6 X.n0 X.t1 123.653
R7 X X.n0 82.224
R8 X.n1 X 10.483
R9 X X.n1 5.504
R10 X.n0 X 5.169
R11 VPWR VPWR.n0 169.297
R12 VPWR.n0 VPWR.t0 36.158
R13 VPWR.n0 VPWR.t1 36.158
R14 VPB.t0 VPB.t1 260.436
R15 VPB VPB.t0 91.744
R16 A.n0 A.t1 260.32
R17 A.n0 A.t0 175.167
R18 A A.n0 78.133
R19 VGND VGND.n0 110.77
R20 VGND.n0 VGND.t0 33.461
R21 VGND.n0 VGND.t1 33.461
R22 VNB VNB.t0 6271.49
R23 VNB.t0 VNB.t1 2482.05
C0 X VPWR 0.14fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__clkbuf_2.ext - technology: sky130A

.subckt sky130_fd_sc_hd__clkbuf_2 A X VGND VPWR VNB VPB
X0 VPWR.t0 A.t0 a_27_47.t1 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 VPWR.t1 a_27_47.t2 X.t3 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 VGND.t0 A.t1 a_27_47.t0 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3 X.t2 a_27_47.t3 VPWR.t2 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 X.t1 a_27_47.t4 VGND.t2 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 VGND.t1 a_27_47.t5 X.t0 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
R0 A.n0 A.t0 224.982
R1 A.n0 A.t1 187.712
R2 A A.n0 77.955
R3 a_27_47.t1 a_27_47.n3 257.015
R4 a_27_47.n3 a_27_47.t0 213.169
R5 a_27_47.n0 a_27_47.t3 189.586
R6 a_27_47.n0 a_27_47.t2 189.586
R7 a_27_47.n3 a_27_47.n2 143.433
R8 a_27_47.n1 a_27_47.t5 96.4
R9 a_27_47.n1 a_27_47.t4 96.4
R10 a_27_47.n2 a_27_47.n1 35.092
R11 a_27_47.n2 a_27_47.n0 19.871
R12 VPWR.n1 VPWR.t1 547.613
R13 VPWR.n1 VPWR.n0 169.858
R14 VPWR.n0 VPWR.t2 36.445
R15 VPWR.n0 VPWR.t0 27.58
R16 VPWR VPWR.n1 0.219
R17 VPB.t0 VPB.t1 281.152
R18 VPB.t1 VPB.t2 248.598
R19 VPB VPB.t0 195.327
R20 X X.n0 331.407
R21 X X.n1 123.962
R22 X.n1 X.t0 38.571
R23 X.n1 X.t1 38.571
R24 X.n0 X.t3 26.595
R25 X.n0 X.t2 26.595
R26 VGND.n1 VGND.t1 150.351
R27 VGND.n1 VGND.n0 114.507
R28 VGND.n0 VGND.t2 52.857
R29 VGND.n0 VGND.t0 40
R30 VGND VGND.n1 0.214
R31 VNB VNB.t0 6502.94
R32 VNB.t0 VNB.t2 3073.53
R33 VNB.t2 VNB.t1 2717.65
C0 VGND X 0.17fF
C1 VPWR X 0.19fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__clkbuf_4.ext - technology: sky130A

.subckt sky130_fd_sc_hd__clkbuf_4 X A VGND VPWR VNB VPB
X0 VPWR.t4 A.t0 a_27_47.t0 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 VGND.t3 a_27_47.t2 X.t7 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 VGND.t2 a_27_47.t3 X.t6 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3 X.t3 a_27_47.t4 VPWR.t3 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 X.t5 a_27_47.t5 VGND.t1 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 VGND.t4 A.t1 a_27_47.t1 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 VPWR.t2 a_27_47.t6 X.t2 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 X.t4 a_27_47.t7 VGND.t0 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 X.t1 a_27_47.t8 VPWR.t1 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 VPWR.t0 a_27_47.t9 X.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
R0 A.n0 A.t0 238.589
R1 A.n0 A.t1 203.243
R2 A A.n0 78.011
R3 a_27_47.t0 a_27_47.n11 270.079
R4 a_27_47.n8 a_27_47.t8 223.188
R5 a_27_47.n0 a_27_47.t6 221.719
R6 a_27_47.n3 a_27_47.t4 221.719
R7 a_27_47.n7 a_27_47.t9 221.719
R8 a_27_47.n11 a_27_47.t1 211.566
R9 a_27_47.n0 a_27_47.t2 185.378
R10 a_27_47.n8 a_27_47.t7 184.766
R11 a_27_47.n6 a_27_47.t3 184.766
R12 a_27_47.n2 a_27_47.t5 184.766
R13 a_27_47.n5 a_27_47.n1 101.6
R14 a_27_47.n11 a_27_47.n10 82.445
R15 a_27_47.n5 a_27_47.n4 76
R16 a_27_47.n10 a_27_47.n9 76
R17 a_27_47.n1 a_27_47.n0 56.963
R18 a_27_47.n9 a_27_47.n8 49.076
R19 a_27_47.n4 a_27_47.n3 41.189
R20 a_27_47.n10 a_27_47.n5 25.6
R21 a_27_47.n9 a_27_47.n7 25.414
R22 a_27_47.n3 a_27_47.n2 0.876
R23 a_27_47.n7 a_27_47.n6 0.876
R24 VPWR.n1 VPWR.n0 311.574
R25 VPWR.n2 VPWR.t2 201.736
R26 VPWR.n6 VPWR.n5 165.368
R27 VPWR.n5 VPWR.t1 37.43
R28 VPWR.n0 VPWR.t3 27.58
R29 VPWR.n0 VPWR.t0 27.58
R30 VPWR.n5 VPWR.t4 27.58
R31 VPWR.n4 VPWR.n3 4.65
R32 VPWR.n7 VPWR.n6 4.01
R33 VPWR.n2 VPWR.n1 3.901
R34 VPWR.n4 VPWR.n2 0.238
R35 VPWR.n7 VPWR.n4 0.135
R36 VPWR VPWR.n7 0.125
R37 VPB.t4 VPB.t1 284.112
R38 VPB.t3 VPB.t2 254.517
R39 VPB.t0 VPB.t3 254.517
R40 VPB.t1 VPB.t0 254.517
R41 VPB VPB.t4 195.327
R42 X.n5 X.n3 354.632
R43 X.n2 X.n0 151.126
R44 X.n2 X.n1 107.761
R45 X.n5 X.n4 96.929
R46 X.n0 X.t6 40
R47 X.n0 X.t4 40
R48 X.n1 X.t7 40
R49 X.n1 X.t5 40
R50 X.n4 X.t2 27.58
R51 X.n4 X.t3 27.58
R52 X.n3 X.t0 27.58
R53 X.n3 X.t1 27.58
R54 X X.n6 19.259
R55 X.n6 X.n5 15.308
R56 X.n7 X 9.007
R57 X.n7 X.n2 6.776
R58 X.n6 X 2.707
R59 X X.n7 1.738
R60 VGND.n2 VGND.t3 154.76
R61 VGND.n1 VGND.n0 112.578
R62 VGND.n6 VGND.n5 111.118
R63 VGND.n5 VGND.t0 55.714
R64 VGND.n0 VGND.t1 40
R65 VGND.n0 VGND.t2 40
R66 VGND.n5 VGND.t4 40
R67 VGND.n4 VGND.n3 4.65
R68 VGND.n7 VGND.n6 3.996
R69 VGND.n2 VGND.n1 3.901
R70 VGND.n4 VGND.n2 0.238
R71 VGND.n7 VGND.n4 0.136
R72 VGND VGND.n7 0.125
R73 VNB VNB.t4 6502.94
R74 VNB.t4 VNB.t0 3138.24
R75 VNB.t1 VNB.t3 2782.35
R76 VNB.t2 VNB.t1 2782.35
R77 VNB.t0 VNB.t2 2782.35
C0 X VGND 0.35fF
C1 VPWR X 0.47fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__clkbuf_8.ext - technology: sky130A

.subckt sky130_fd_sc_hd__clkbuf_8 X A VGND VPWR VNB VPB
X0 VPWR.t1 A.t0 a_110_47.t1 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 VPWR.t9 a_110_47.t4 X.t15 VPB.t9 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 X.t14 a_110_47.t5 VPWR.t8 VPB.t8 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 a_110_47.t0 A.t1 VPWR.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 X.t5 a_110_47.t6 VGND.t9 VNB.t9 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 X.t13 a_110_47.t7 VPWR.t7 VPB.t7 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 VGND.t8 a_110_47.t8 X.t4 VNB.t8 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7 VPWR.t6 a_110_47.t9 X.t12 VPB.t6 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 VGND.t1 A.t2 a_110_47.t3 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9 VGND.t7 a_110_47.t10 X.t3 VNB.t7 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10 a_110_47.t2 A.t3 VGND.t0 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11 VPWR.t5 a_110_47.t11 X.t11 VPB.t5 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 X.t10 a_110_47.t12 VPWR.t4 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13 VGND.t6 a_110_47.t13 X.t2 VNB.t6 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14 VGND.t5 a_110_47.t14 X.t1 VNB.t5 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15 X.t9 a_110_47.t15 VPWR.t3 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16 X.t0 a_110_47.t16 VGND.t4 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17 VPWR.t2 a_110_47.t17 X.t8 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X18 X.t7 a_110_47.t18 VGND.t3 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19 X.t6 a_110_47.t19 VGND.t2 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
R0 A.n0 A.t0 184.766
R1 A.n1 A.t1 184.766
R2 A.n0 A.t2 146.206
R3 A.n1 A.t3 146.206
R4 A A.n1 97.608
R5 A.n1 A.n0 40.639
R6 a_110_47.n1 a_110_47.t17 212.079
R7 a_110_47.n2 a_110_47.t12 212.079
R8 a_110_47.n3 a_110_47.t9 212.079
R9 a_110_47.n5 a_110_47.t5 212.079
R10 a_110_47.n8 a_110_47.t4 212.079
R11 a_110_47.n11 a_110_47.t15 212.079
R12 a_110_47.n16 a_110_47.t11 212.079
R13 a_110_47.n17 a_110_47.t7 212.079
R14 a_110_47.n21 a_110_47.n20 170.244
R15 a_110_47.n1 a_110_47.t10 162.273
R16 a_110_47.n2 a_110_47.t16 162.273
R17 a_110_47.n3 a_110_47.t13 162.273
R18 a_110_47.n5 a_110_47.t18 162.273
R19 a_110_47.n8 a_110_47.t14 162.273
R20 a_110_47.n11 a_110_47.t19 162.273
R21 a_110_47.n16 a_110_47.t8 162.273
R22 a_110_47.n17 a_110_47.t6 162.273
R23 a_110_47.n20 a_110_47.n0 124.756
R24 a_110_47.n7 a_110_47.n4 93.408
R25 a_110_47.n19 a_110_47.n18 76
R26 a_110_47.n7 a_110_47.n6 76
R27 a_110_47.n10 a_110_47.n9 76
R28 a_110_47.n13 a_110_47.n12 76
R29 a_110_47.n15 a_110_47.n14 76
R30 a_110_47.n2 a_110_47.n1 55.269
R31 a_110_47.n3 a_110_47.n2 55.269
R32 a_110_47.n20 a_110_47.n19 43.52
R33 a_110_47.n0 a_110_47.t3 40
R34 a_110_47.n0 a_110_47.t2 40
R35 a_110_47.n4 a_110_47.n3 30.848
R36 a_110_47.n18 a_110_47.n16 28.277
R37 a_110_47.n21 a_110_47.t1 27.58
R38 a_110_47.t0 a_110_47.n21 27.58
R39 a_110_47.n18 a_110_47.n17 26.992
R40 a_110_47.n6 a_110_47.n5 19.28
R41 a_110_47.n10 a_110_47.n7 17.408
R42 a_110_47.n13 a_110_47.n10 17.408
R43 a_110_47.n15 a_110_47.n13 17.408
R44 a_110_47.n19 a_110_47.n15 17.408
R45 a_110_47.n9 a_110_47.n8 7.712
R46 a_110_47.n12 a_110_47.n11 3.856
R47 VPWR.n2 VPWR.t2 493.844
R48 VPWR.n12 VPWR.n11 317.115
R49 VPWR.n6 VPWR.n5 317.115
R50 VPWR.n1 VPWR.n0 317.115
R51 VPWR.n21 VPWR.t0 204.384
R52 VPWR.n17 VPWR.n16 180.896
R53 VPWR.n16 VPWR.t7 27.58
R54 VPWR.n16 VPWR.t1 27.58
R55 VPWR.n11 VPWR.t3 27.58
R56 VPWR.n11 VPWR.t5 27.58
R57 VPWR.n5 VPWR.t8 27.58
R58 VPWR.n5 VPWR.t9 27.58
R59 VPWR.n0 VPWR.t4 27.58
R60 VPWR.n0 VPWR.t6 27.58
R61 VPWR.n2 VPWR.n1 9.867
R62 VPWR.n4 VPWR.n3 4.65
R63 VPWR.n8 VPWR.n7 4.65
R64 VPWR.n10 VPWR.n9 4.65
R65 VPWR.n13 VPWR.n12 4.65
R66 VPWR.n15 VPWR.n14 4.65
R67 VPWR.n18 VPWR.n17 4.65
R68 VPWR.n20 VPWR.n19 4.65
R69 VPWR.n22 VPWR.n21 4.65
R70 VPWR.n7 VPWR.n6 1.505
R71 VPWR.n4 VPWR.n2 0.424
R72 VPWR.n8 VPWR.n4 0.119
R73 VPWR.n10 VPWR.n8 0.119
R74 VPWR.n13 VPWR.n10 0.119
R75 VPWR.n15 VPWR.n13 0.119
R76 VPWR.n18 VPWR.n15 0.119
R77 VPWR.n20 VPWR.n18 0.119
R78 VPWR.n22 VPWR.n20 0.119
R79 VPWR VPWR.n22 0.022
R80 VPB.t4 VPB.t2 254.517
R81 VPB.t6 VPB.t4 254.517
R82 VPB.t8 VPB.t6 254.517
R83 VPB.t9 VPB.t8 254.517
R84 VPB.t3 VPB.t9 254.517
R85 VPB.t5 VPB.t3 254.517
R86 VPB.t7 VPB.t5 254.517
R87 VPB.t1 VPB.t7 254.517
R88 VPB.t0 VPB.t1 254.517
R89 VPB VPB.t0 195.327
R90 X.n7 X.n5 187.05
R91 X.n2 X.n0 156.137
R92 X.n7 X.n6 155.05
R93 X.n9 X.n8 155.05
R94 X.n11 X.n10 151.969
R95 X.n2 X.n1 110.961
R96 X.n4 X.n3 110.961
R97 X X.n13 107.171
R98 X.n4 X.n2 45.176
R99 X.n0 X.t4 40
R100 X.n0 X.t5 40
R101 X.n1 X.t1 40
R102 X.n1 X.t6 40
R103 X.n3 X.t2 40
R104 X.n3 X.t7 40
R105 X.n13 X.t3 40
R106 X.n13 X.t0 40
R107 X.n9 X.n7 32
R108 X.n5 X.t11 27.58
R109 X.n5 X.t13 27.58
R110 X.n6 X.t15 27.58
R111 X.n6 X.t9 27.58
R112 X.n8 X.t12 27.58
R113 X.n8 X.t14 27.58
R114 X.n10 X.t8 27.58
R115 X.n10 X.t10 27.58
R116 X.n12 X.n4 27.105
R117 X.n11 X.n9 19.2
R118 X.n12 X 3.76
R119 X X.n11 2.243
R120 X X.n12 0.725
R121 VGND.n2 VGND.t7 155.887
R122 VGND.n21 VGND.t0 152.353
R123 VGND.n17 VGND.n16 114.407
R124 VGND.n1 VGND.n0 112.192
R125 VGND.n6 VGND.n5 112.192
R126 VGND.n12 VGND.n11 112.192
R127 VGND.n0 VGND.t4 40
R128 VGND.n0 VGND.t6 40
R129 VGND.n5 VGND.t3 40
R130 VGND.n5 VGND.t5 40
R131 VGND.n11 VGND.t2 40
R132 VGND.n11 VGND.t8 40
R133 VGND.n16 VGND.t9 40
R134 VGND.n16 VGND.t1 40
R135 VGND.n2 VGND.n1 9.871
R136 VGND.n22 VGND.n21 4.65
R137 VGND.n4 VGND.n3 4.65
R138 VGND.n8 VGND.n7 4.65
R139 VGND.n10 VGND.n9 4.65
R140 VGND.n13 VGND.n12 4.65
R141 VGND.n15 VGND.n14 4.65
R142 VGND.n18 VGND.n17 4.65
R143 VGND.n20 VGND.n19 4.65
R144 VGND.n7 VGND.n6 1.505
R145 VGND.n4 VGND.n2 0.42
R146 VGND.n8 VGND.n4 0.119
R147 VGND.n10 VGND.n8 0.119
R148 VGND.n13 VGND.n10 0.119
R149 VGND.n15 VGND.n13 0.119
R150 VGND.n18 VGND.n15 0.119
R151 VGND.n20 VGND.n18 0.119
R152 VGND.n22 VGND.n20 0.119
R153 VGND VGND.n22 0.022
R154 VNB VNB.t0 6502.94
R155 VNB.t4 VNB.t7 2782.35
R156 VNB.t6 VNB.t4 2782.35
R157 VNB.t3 VNB.t6 2782.35
R158 VNB.t5 VNB.t3 2782.35
R159 VNB.t2 VNB.t5 2782.35
R160 VNB.t8 VNB.t2 2782.35
R161 VNB.t9 VNB.t8 2782.35
R162 VNB.t1 VNB.t9 2782.35
R163 VNB.t0 VNB.t1 2782.35
C0 VPB VPWR 0.11fF
C1 X VGND 0.80fF
C2 VGND VPWR 0.12fF
C3 X VPWR 1.21fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__clkbuf_16.ext - technology: sky130A

.subckt sky130_fd_sc_hd__clkbuf_16 X A VGND VPWR VNB VPB
X0 VPWR.t3 A.t0 a_110_47.t7 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 VPWR.t19 a_110_47.t8 X.t18 VPB.t19 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 X.t17 a_110_47.t9 VPWR.t18 VPB.t18 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 X.t16 a_110_47.t10 VPWR.t17 VPB.t17 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 VPWR.t16 a_110_47.t11 X.t15 VPB.t16 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 VPWR.t15 a_110_47.t12 X.t14 VPB.t15 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 a_110_47.t6 A.t1 VPWR.t2 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 a_110_47.t3 A.t2 VGND.t3 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 VGND.t19 a_110_47.t13 X.t24 VNB.t19 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9 X.t23 a_110_47.t14 VGND.t18 VNB.t18 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10 VGND.t17 a_110_47.t15 X.t22 VNB.t17 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11 a_110_47.t5 A.t3 VPWR.t1 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 VGND.t2 A.t4 a_110_47.t2 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13 VGND.t16 a_110_47.t16 X.t21 VNB.t16 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14 VPWR.t14 a_110_47.t17 X.t13 VPB.t14 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 X.t12 a_110_47.t18 VPWR.t13 VPB.t13 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16 VGND.t1 A.t5 a_110_47.t1 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17 VGND.t15 a_110_47.t19 X.t20 VNB.t15 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18 VPWR.t12 a_110_47.t20 X.t11 VPB.t12 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X19 VGND.t14 a_110_47.t21 X.t19 VNB.t14 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20 X.t10 a_110_47.t22 VPWR.t11 VPB.t11 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X21 a_110_47.t0 A.t6 VGND.t0 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22 VPWR.t0 A.t7 a_110_47.t4 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X23 VPWR.t10 a_110_47.t23 X.t9 VPB.t10 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X24 VPWR.t9 a_110_47.t24 X.t8 VPB.t9 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X25 VGND.t13 a_110_47.t25 X.t31 VNB.t13 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X26 X.t7 a_110_47.t26 VPWR.t8 VPB.t8 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X27 VGND.t12 a_110_47.t27 X.t30 VNB.t12 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X28 VGND.t11 a_110_47.t28 X.t29 VNB.t11 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X29 X.t28 a_110_47.t29 VGND.t10 VNB.t10 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X30 X.t6 a_110_47.t30 VPWR.t7 VPB.t7 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X31 X.t5 a_110_47.t31 VPWR.t6 VPB.t6 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X32 X.t27 a_110_47.t32 VGND.t9 VNB.t9 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X33 VPWR.t5 a_110_47.t33 X.t4 VPB.t5 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X34 X.t3 a_110_47.t34 VPWR.t4 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X35 X.t26 a_110_47.t35 VGND.t8 VNB.t8 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X36 X.t25 a_110_47.t36 VGND.t7 VNB.t7 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X37 X.t2 a_110_47.t37 VGND.t6 VNB.t6 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X38 X.t1 a_110_47.t38 VGND.t5 VNB.t5 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X39 X.t0 a_110_47.t39 VGND.t4 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
R0 A.n0 A.t7 184.766
R1 A.n1 A.t3 184.766
R2 A.n2 A.t0 184.766
R3 A.n3 A.t1 184.766
R4 A.n0 A.t4 146.206
R5 A.n1 A.t2 146.206
R6 A.n2 A.t5 146.206
R7 A.n3 A.t6 146.206
R8 A A.n3 97.608
R9 A.n1 A.n0 40.639
R10 A.n2 A.n1 40.639
R11 A.n3 A.n2 40.639
R12 a_110_47.n1 a_110_47.t12 212.079
R13 a_110_47.n2 a_110_47.t34 212.079
R14 a_110_47.n3 a_110_47.t24 212.079
R15 a_110_47.n5 a_110_47.t18 212.079
R16 a_110_47.n8 a_110_47.t11 212.079
R17 a_110_47.n11 a_110_47.t30 212.079
R18 a_110_47.n14 a_110_47.t23 212.079
R19 a_110_47.n19 a_110_47.t22 212.079
R20 a_110_47.n22 a_110_47.t20 212.079
R21 a_110_47.n25 a_110_47.t10 212.079
R22 a_110_47.n28 a_110_47.t33 212.079
R23 a_110_47.n33 a_110_47.t26 212.079
R24 a_110_47.n36 a_110_47.t17 212.079
R25 a_110_47.n39 a_110_47.t9 212.079
R26 a_110_47.n44 a_110_47.t8 212.079
R27 a_110_47.n45 a_110_47.t31 212.079
R28 a_110_47.n50 a_110_47.n49 183.992
R29 a_110_47.n52 a_110_47.n51 180.942
R30 a_110_47.n1 a_110_47.t19 162.273
R31 a_110_47.n2 a_110_47.t29 162.273
R32 a_110_47.n3 a_110_47.t25 162.273
R33 a_110_47.n5 a_110_47.t35 162.273
R34 a_110_47.n8 a_110_47.t13 162.273
R35 a_110_47.n11 a_110_47.t37 162.273
R36 a_110_47.n14 a_110_47.t15 162.273
R37 a_110_47.n19 a_110_47.t39 162.273
R38 a_110_47.n22 a_110_47.t16 162.273
R39 a_110_47.n25 a_110_47.t14 162.273
R40 a_110_47.n28 a_110_47.t21 162.273
R41 a_110_47.n33 a_110_47.t32 162.273
R42 a_110_47.n36 a_110_47.t27 162.273
R43 a_110_47.n39 a_110_47.t36 162.273
R44 a_110_47.n44 a_110_47.t28 162.273
R45 a_110_47.n45 a_110_47.t38 162.273
R46 a_110_47.n51 a_110_47.n0 124.756
R47 a_110_47.n50 a_110_47.n48 124.756
R48 a_110_47.n7 a_110_47.n4 93.408
R49 a_110_47.n47 a_110_47.n46 76
R50 a_110_47.n7 a_110_47.n6 76
R51 a_110_47.n10 a_110_47.n9 76
R52 a_110_47.n13 a_110_47.n12 76
R53 a_110_47.n16 a_110_47.n15 76
R54 a_110_47.n18 a_110_47.n17 76
R55 a_110_47.n21 a_110_47.n20 76
R56 a_110_47.n24 a_110_47.n23 76
R57 a_110_47.n27 a_110_47.n26 76
R58 a_110_47.n30 a_110_47.n29 76
R59 a_110_47.n32 a_110_47.n31 76
R60 a_110_47.n35 a_110_47.n34 76
R61 a_110_47.n38 a_110_47.n37 76
R62 a_110_47.n41 a_110_47.n40 76
R63 a_110_47.n43 a_110_47.n42 76
R64 a_110_47.n2 a_110_47.n1 55.269
R65 a_110_47.n3 a_110_47.n2 55.269
R66 a_110_47.n51 a_110_47.n50 44.032
R67 a_110_47.n51 a_110_47.n47 43.52
R68 a_110_47.n0 a_110_47.t2 40
R69 a_110_47.n0 a_110_47.t3 40
R70 a_110_47.n48 a_110_47.t1 40
R71 a_110_47.n48 a_110_47.t0 40
R72 a_110_47.n4 a_110_47.n3 35.346
R73 a_110_47.n46 a_110_47.n44 28.277
R74 a_110_47.n49 a_110_47.t7 27.58
R75 a_110_47.n49 a_110_47.t6 27.58
R76 a_110_47.t4 a_110_47.n52 27.58
R77 a_110_47.n52 a_110_47.t5 27.58
R78 a_110_47.n46 a_110_47.n45 26.992
R79 a_110_47.n6 a_110_47.n5 23.778
R80 a_110_47.n20 a_110_47.n19 21.208
R81 a_110_47.n34 a_110_47.n33 19.28
R82 a_110_47.n10 a_110_47.n7 17.408
R83 a_110_47.n13 a_110_47.n10 17.408
R84 a_110_47.n16 a_110_47.n13 17.408
R85 a_110_47.n18 a_110_47.n16 17.408
R86 a_110_47.n21 a_110_47.n18 17.408
R87 a_110_47.n24 a_110_47.n21 17.408
R88 a_110_47.n27 a_110_47.n24 17.408
R89 a_110_47.n30 a_110_47.n27 17.408
R90 a_110_47.n32 a_110_47.n30 17.408
R91 a_110_47.n35 a_110_47.n32 17.408
R92 a_110_47.n38 a_110_47.n35 17.408
R93 a_110_47.n41 a_110_47.n38 17.408
R94 a_110_47.n43 a_110_47.n41 17.408
R95 a_110_47.n47 a_110_47.n43 17.408
R96 a_110_47.n29 a_110_47.n28 12.853
R97 a_110_47.n9 a_110_47.n8 12.21
R98 a_110_47.n15 a_110_47.n14 10.925
R99 a_110_47.n23 a_110_47.n22 10.282
R100 a_110_47.n37 a_110_47.n36 7.712
R101 a_110_47.n40 a_110_47.n39 3.856
R102 a_110_47.n26 a_110_47.n25 1.285
R103 a_110_47.n12 a_110_47.n11 0.642
R104 VPWR.n2 VPWR.t15 494.84
R105 VPWR.n16 VPWR.n15 318.361
R106 VPWR.n11 VPWR.n10 318.361
R107 VPWR.n6 VPWR.n5 318.361
R108 VPWR.n1 VPWR.n0 317.347
R109 VPWR.n31 VPWR.n30 316.869
R110 VPWR.n25 VPWR.n24 316.869
R111 VPWR.n21 VPWR.n20 316.869
R112 VPWR.n47 VPWR.t2 193.916
R113 VPWR.n43 VPWR.n42 169.026
R114 VPWR.n37 VPWR.n36 168.78
R115 VPWR.n42 VPWR.t1 27.58
R116 VPWR.n42 VPWR.t3 27.58
R117 VPWR.n0 VPWR.t4 27.58
R118 VPWR.n0 VPWR.t9 27.58
R119 VPWR.n36 VPWR.t6 27.58
R120 VPWR.n36 VPWR.t0 27.58
R121 VPWR.n30 VPWR.t18 27.58
R122 VPWR.n30 VPWR.t19 27.58
R123 VPWR.n24 VPWR.t8 27.58
R124 VPWR.n24 VPWR.t14 27.58
R125 VPWR.n20 VPWR.t17 27.58
R126 VPWR.n20 VPWR.t5 27.58
R127 VPWR.n15 VPWR.t12 27.58
R128 VPWR.n10 VPWR.t7 27.58
R129 VPWR.n10 VPWR.t10 27.58
R130 VPWR.n5 VPWR.t13 27.58
R131 VPWR.n5 VPWR.t16 27.58
R132 VPWR.n15 VPWR.t11 26.595
R133 VPWR.n26 VPWR.n25 5.851
R134 VPWR.n17 VPWR.n16 4.911
R135 VPWR.n12 VPWR.n11 4.911
R136 VPWR.n7 VPWR.n6 4.911
R137 VPWR.n4 VPWR.n3 4.65
R138 VPWR.n9 VPWR.n8 4.65
R139 VPWR.n14 VPWR.n13 4.65
R140 VPWR.n19 VPWR.n18 4.65
R141 VPWR.n23 VPWR.n22 4.65
R142 VPWR.n27 VPWR.n26 4.65
R143 VPWR.n29 VPWR.n28 4.65
R144 VPWR.n33 VPWR.n32 4.65
R145 VPWR.n35 VPWR.n34 4.65
R146 VPWR.n39 VPWR.n38 4.65
R147 VPWR.n41 VPWR.n40 4.65
R148 VPWR.n44 VPWR.n43 4.65
R149 VPWR.n46 VPWR.n45 4.65
R150 VPWR.n48 VPWR.n47 4.65
R151 VPWR.n22 VPWR.n21 4.388
R152 VPWR.n2 VPWR.n1 4.213
R153 VPWR.n32 VPWR.n31 1.462
R154 VPWR.n38 VPWR.n37 0.246
R155 VPWR.n4 VPWR.n2 0.233
R156 VPWR.n7 VPWR.n4 0.119
R157 VPWR.n9 VPWR.n7 0.119
R158 VPWR.n12 VPWR.n9 0.119
R159 VPWR.n14 VPWR.n12 0.119
R160 VPWR.n17 VPWR.n14 0.119
R161 VPWR.n19 VPWR.n17 0.119
R162 VPWR.n23 VPWR.n19 0.119
R163 VPWR.n27 VPWR.n23 0.119
R164 VPWR.n29 VPWR.n27 0.119
R165 VPWR.n33 VPWR.n29 0.119
R166 VPWR.n35 VPWR.n33 0.119
R167 VPWR.n39 VPWR.n35 0.119
R168 VPWR.n41 VPWR.n39 0.119
R169 VPWR.n44 VPWR.n41 0.119
R170 VPWR.n46 VPWR.n44 0.119
R171 VPWR.n48 VPWR.n46 0.119
R172 VPWR VPWR.n48 0.022
R173 VPB.t4 VPB.t15 254.517
R174 VPB.t9 VPB.t4 254.517
R175 VPB.t13 VPB.t9 254.517
R176 VPB.t16 VPB.t13 254.517
R177 VPB.t7 VPB.t16 254.517
R178 VPB.t10 VPB.t7 254.517
R179 VPB.t11 VPB.t10 254.517
R180 VPB.t17 VPB.t12 254.517
R181 VPB.t5 VPB.t17 254.517
R182 VPB.t8 VPB.t5 254.517
R183 VPB.t14 VPB.t8 254.517
R184 VPB.t18 VPB.t14 254.517
R185 VPB.t19 VPB.t18 254.517
R186 VPB.t6 VPB.t19 254.517
R187 VPB.t0 VPB.t6 254.517
R188 VPB.t1 VPB.t0 254.517
R189 VPB.t3 VPB.t1 254.517
R190 VPB.t2 VPB.t3 254.517
R191 VPB.t12 VPB.t11 251.557
R192 VPB VPB.t2 145.015
R193 X.n15 X.n13 187.05
R194 X.n2 X.n0 156.137
R195 X.n15 X.n14 155.05
R196 X.n17 X.n16 155.05
R197 X.n19 X.n18 155.05
R198 X.n21 X.n20 155.05
R199 X.n23 X.n22 155.05
R200 X.n25 X.n24 155.05
R201 X.n27 X.n26 151.546
R202 X.n2 X.n1 110.961
R203 X.n4 X.n3 110.961
R204 X.n8 X.n7 110.961
R205 X.n10 X.n9 110.961
R206 X.n12 X.n11 110.961
R207 X.n6 X.n5 109.954
R208 X X.n29 107.105
R209 X.n4 X.n2 45.176
R210 X.n10 X.n8 45.176
R211 X.n12 X.n10 45.176
R212 X.n6 X.n4 44.047
R213 X.n8 X.n6 44.047
R214 X.n0 X.t29 40
R215 X.n0 X.t1 40
R216 X.n1 X.t30 40
R217 X.n1 X.t25 40
R218 X.n3 X.t19 40
R219 X.n3 X.t27 40
R220 X.n5 X.t21 40
R221 X.n5 X.t23 40
R222 X.n7 X.t22 40
R223 X.n7 X.t0 40
R224 X.n9 X.t24 40
R225 X.n9 X.t2 40
R226 X.n11 X.t31 40
R227 X.n11 X.t26 40
R228 X.n29 X.t20 40
R229 X.n29 X.t28 40
R230 X.n17 X.n15 32
R231 X.n19 X.n17 32
R232 X.n23 X.n21 32
R233 X.n25 X.n23 32
R234 X.n21 X.n19 31.2
R235 X.n24 X.t8 27.58
R236 X.n24 X.t12 27.58
R237 X.n13 X.t18 27.58
R238 X.n13 X.t5 27.58
R239 X.n14 X.t13 27.58
R240 X.n14 X.t17 27.58
R241 X.n16 X.t4 27.58
R242 X.n16 X.t7 27.58
R243 X.n18 X.t11 27.58
R244 X.n18 X.t16 27.58
R245 X.n20 X.t9 27.58
R246 X.n20 X.t10 27.58
R247 X.n22 X.t15 27.58
R248 X.n22 X.t6 27.58
R249 X.n26 X.t14 27.58
R250 X.n26 X.t3 27.58
R251 X.n28 X.n12 13.176
R252 X.n27 X.n25 10.447
R253 X.n28 X 3.131
R254 X X.n27 1.757
R255 X X.n28 0.604
R256 VGND.n2 VGND.t15 153.42
R257 VGND.n46 VGND.t0 148.447
R258 VGND.n37 VGND.n36 114.407
R259 VGND.n42 VGND.n41 114.407
R260 VGND.n16 VGND.n15 113.397
R261 VGND.n21 VGND.n20 113.397
R262 VGND.n6 VGND.n5 112.98
R263 VGND.n11 VGND.n10 112.98
R264 VGND.n1 VGND.n0 112.192
R265 VGND.n25 VGND.n24 112.192
R266 VGND.n31 VGND.n30 112.192
R267 VGND.n0 VGND.t10 40
R268 VGND.n0 VGND.t13 40
R269 VGND.n5 VGND.t8 40
R270 VGND.n5 VGND.t19 40
R271 VGND.n10 VGND.t6 40
R272 VGND.n10 VGND.t17 40
R273 VGND.n15 VGND.t16 40
R274 VGND.n20 VGND.t18 40
R275 VGND.n20 VGND.t14 40
R276 VGND.n24 VGND.t9 40
R277 VGND.n24 VGND.t12 40
R278 VGND.n30 VGND.t7 40
R279 VGND.n30 VGND.t11 40
R280 VGND.n36 VGND.t5 40
R281 VGND.n36 VGND.t2 40
R282 VGND.n41 VGND.t3 40
R283 VGND.n41 VGND.t1 40
R284 VGND.n15 VGND.t4 38.571
R285 VGND.n26 VGND.n25 6.023
R286 VGND.n47 VGND.n46 4.65
R287 VGND.n4 VGND.n3 4.65
R288 VGND.n7 VGND.n6 4.65
R289 VGND.n9 VGND.n8 4.65
R290 VGND.n12 VGND.n11 4.65
R291 VGND.n14 VGND.n13 4.65
R292 VGND.n17 VGND.n16 4.65
R293 VGND.n19 VGND.n18 4.65
R294 VGND.n23 VGND.n22 4.65
R295 VGND.n27 VGND.n26 4.65
R296 VGND.n29 VGND.n28 4.65
R297 VGND.n33 VGND.n32 4.65
R298 VGND.n35 VGND.n34 4.65
R299 VGND.n38 VGND.n37 4.65
R300 VGND.n40 VGND.n39 4.65
R301 VGND.n43 VGND.n42 4.65
R302 VGND.n45 VGND.n44 4.65
R303 VGND.n22 VGND.n21 4.517
R304 VGND.n2 VGND.n1 3.953
R305 VGND.n32 VGND.n31 1.505
R306 VGND.n4 VGND.n2 0.242
R307 VGND.n7 VGND.n4 0.119
R308 VGND.n9 VGND.n7 0.119
R309 VGND.n12 VGND.n9 0.119
R310 VGND.n14 VGND.n12 0.119
R311 VGND.n17 VGND.n14 0.119
R312 VGND.n19 VGND.n17 0.119
R313 VGND.n23 VGND.n19 0.119
R314 VGND.n27 VGND.n23 0.119
R315 VGND.n29 VGND.n27 0.119
R316 VGND.n33 VGND.n29 0.119
R317 VGND.n35 VGND.n33 0.119
R318 VGND.n38 VGND.n35 0.119
R319 VGND.n40 VGND.n38 0.119
R320 VGND.n43 VGND.n40 0.119
R321 VGND.n45 VGND.n43 0.119
R322 VGND.n47 VGND.n45 0.119
R323 VGND VGND.n47 0.022
R324 VNB VNB.t0 4302.94
R325 VNB.t10 VNB.t15 2782.35
R326 VNB.t13 VNB.t10 2782.35
R327 VNB.t8 VNB.t13 2782.35
R328 VNB.t19 VNB.t8 2782.35
R329 VNB.t6 VNB.t19 2782.35
R330 VNB.t17 VNB.t6 2782.35
R331 VNB.t4 VNB.t17 2782.35
R332 VNB.t18 VNB.t16 2782.35
R333 VNB.t14 VNB.t18 2782.35
R334 VNB.t9 VNB.t14 2782.35
R335 VNB.t12 VNB.t9 2782.35
R336 VNB.t7 VNB.t12 2782.35
R337 VNB.t11 VNB.t7 2782.35
R338 VNB.t5 VNB.t11 2782.35
R339 VNB.t2 VNB.t5 2782.35
R340 VNB.t3 VNB.t2 2782.35
R341 VNB.t1 VNB.t3 2782.35
R342 VNB.t0 VNB.t1 2782.35
R343 VNB.t16 VNB.t4 2750
C0 VGND X 1.57fF
C1 VGND VPWR 0.21fF
C2 VPWR X 2.31fF
C3 VPB VPWR 0.19fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__clkdlybuf4s15_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__clkdlybuf4s15_1 VGND VPWR A X VNB VPB
X0 VPWR.t1 A.t0 a_27_47.t0 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_282_47.t0 a_27_47.t2 VGND.t2 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 X.t0 a_394_47.t2 VGND.t0 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3 VGND.t3 a_282_47.t2 a_394_47.t0 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 X.t1 a_394_47.t3 VPWR.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 a_282_47.t1 a_27_47.t3 VPWR.t2 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=820000u l=150000u
X6 VGND.t1 A.t1 a_27_47.t1 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7 VPWR.t3 a_282_47.t3 a_394_47.t1 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=820000u l=150000u
R0 A.n0 A.t0 236.179
R1 A.n0 A.t1 206.091
R2 A A.n0 87.851
R3 a_27_47.n0 a_27_47.t3 250.639
R4 a_27_47.t0 a_27_47.n1 225.505
R5 a_27_47.n1 a_27_47.t1 180.776
R6 a_27_47.n1 a_27_47.n0 140.266
R7 a_27_47.n0 a_27_47.t2 139.779
R8 VPWR.n2 VPWR.n1 174.111
R9 VPWR.n2 VPWR.n0 168.571
R10 VPWR.n0 VPWR.t3 112.888
R11 VPWR.n1 VPWR.t2 110.653
R12 VPWR.n0 VPWR.t0 33.528
R13 VPWR.n1 VPWR.t1 29.521
R14 VPWR VPWR.n2 0.151
R15 VPB.t2 VPB.t3 577.102
R16 VPB.t3 VPB.t0 509.034
R17 VPB.t1 VPB.t2 509.034
R18 VPB VPB.t1 195.327
R19 VGND.n2 VGND.n1 111.347
R20 VGND.n2 VGND.n0 111.121
R21 VGND.n1 VGND.t2 95.076
R22 VGND.n0 VGND.t3 90.461
R23 VGND.n0 VGND.t0 51.735
R24 VGND.n1 VGND.t1 43.581
R25 VGND VGND.n2 0.15
R26 a_282_47.n0 a_282_47.t3 239.392
R27 a_282_47.t1 a_282_47.n1 232.41
R28 a_282_47.n0 a_282_47.t2 141.386
R29 a_282_47.n1 a_282_47.t0 108.239
R30 a_282_47.n1 a_282_47.n0 87.409
R31 VNB VNB.t1 6502.94
R32 VNB.t2 VNB.t3 4714.29
R33 VNB.t1 VNB.t2 4116.88
R34 VNB.t3 VNB.t0 4044.51
R35 a_394_47.n1 a_394_47.t0 248.651
R36 a_394_47.t1 a_394_47.n1 241.811
R37 a_394_47.n0 a_394_47.t3 235.302
R38 a_394_47.n0 a_394_47.t2 201.709
R39 a_394_47.n1 a_394_47.n0 76
R40 X.n1 X.t1 174.565
R41 X X.t0 133.996
R42 X X.n0 12.243
R43 X.n1 X 9.187
R44 X.n0 X 6.678
R45 X.n0 X 3.989
R46 X X.n1 2.088
C0 VGND X 0.10fF
C1 VPWR X 0.19fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__clkdlybuf4s15_2.ext - technology: sky130A

.subckt sky130_fd_sc_hd__clkdlybuf4s15_2 A X VPWR VGND VNB VPB
X0 VPWR.t2 A.t0 a_27_47.t1 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 VGND.t1 a_362_333.t2 X.t1 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 VPWR.t0 a_228_47.t2 a_362_333.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=820000u l=150000u
X3 VGND.t2 A.t1 a_27_47.t0 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 X.t3 a_362_333.t3 VPWR.t1 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 X.t0 a_362_333.t4 VGND.t0 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 VPWR.t3 a_362_333.t5 X.t2 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 VGND.t3 a_228_47.t3 a_362_333.t1 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 a_228_47.t1 a_27_47.t2 VPWR.t4 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=820000u l=150000u
X9 a_228_47.t0 a_27_47.t3 VGND.t4 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
R0 A.n0 A.t0 241.142
R1 A.n0 A.t1 205.796
R2 A.n1 A.n0 76
R3 A.n1 A 7.761
R4 A A.n1 1.497
R5 a_27_47.n0 a_27_47.t2 270.357
R6 a_27_47.t1 a_27_47.n1 262.333
R7 a_27_47.n1 a_27_47.t0 203.526
R8 a_27_47.n0 a_27_47.t3 169.137
R9 a_27_47.n1 a_27_47.n0 89.552
R10 VPWR.n2 VPWR.n1 308.79
R11 VPWR.n12 VPWR.n11 308.79
R12 VPWR.n0 VPWR.t3 242.35
R13 VPWR.n1 VPWR.t0 117.719
R14 VPWR.n11 VPWR.t4 54.054
R15 VPWR.n1 VPWR.t1 49.657
R16 VPWR.n11 VPWR.t2 47.254
R17 VPWR.n4 VPWR.n3 4.65
R18 VPWR.n6 VPWR.n5 4.65
R19 VPWR.n8 VPWR.n7 4.65
R20 VPWR.n10 VPWR.n9 4.65
R21 VPWR.n13 VPWR.n12 4.056
R22 VPWR.n3 VPWR.n2 1.505
R23 VPWR.n4 VPWR.n0 0.213
R24 VPWR.n13 VPWR.n10 0.134
R25 VPWR VPWR.n13 0.124
R26 VPWR.n6 VPWR.n4 0.119
R27 VPWR.n8 VPWR.n6 0.119
R28 VPWR.n10 VPWR.n8 0.119
R29 VPB.t4 VPB.t0 642.211
R30 VPB.t0 VPB.t1 509.034
R31 VPB.t2 VPB.t4 346.261
R32 VPB.t1 VPB.t3 254.517
R33 VPB VPB.t2 195.327
R34 a_362_333.t0 a_362_333.n3 281.168
R35 a_362_333.n3 a_362_333.t1 242.712
R36 a_362_333.n0 a_362_333.t5 221.719
R37 a_362_333.n1 a_362_333.t3 221.719
R38 a_362_333.n0 a_362_333.t2 186.373
R39 a_362_333.n1 a_362_333.t4 186.373
R40 a_362_333.n3 a_362_333.n2 91.435
R41 a_362_333.n2 a_362_333.n0 74.977
R42 a_362_333.n2 a_362_333.n1 1.785
R43 X.n3 X.n2 145.63
R44 X X.n0 97.154
R45 X.n0 X.t1 40
R46 X.n0 X.t0 40
R47 X.n2 X.t2 27.58
R48 X.n2 X.t3 27.58
R49 X X.n1 8
R50 X.n3 X 5.395
R51 X X.n3 3.585
R52 X.n1 X 2.625
R53 X.n1 X 1.066
R54 VGND.n0 VGND.t1 216.848
R55 VGND.n1 VGND.t3 126.857
R56 VGND.n12 VGND.n11 108.79
R57 VGND.n2 VGND.n1 108.015
R58 VGND.n1 VGND.t0 62.857
R59 VGND.n11 VGND.t2 55.714
R60 VGND.n11 VGND.t4 51.889
R61 VGND.n4 VGND.n3 4.65
R62 VGND.n6 VGND.n5 4.65
R63 VGND.n8 VGND.n7 4.65
R64 VGND.n10 VGND.n9 4.65
R65 VGND.n13 VGND.n12 4.037
R66 VGND.n3 VGND.n2 1.505
R67 VGND.n4 VGND.n0 0.212
R68 VGND.n13 VGND.n10 0.135
R69 VGND VGND.n13 0.124
R70 VGND.n6 VGND.n4 0.119
R71 VGND.n8 VGND.n6 0.119
R72 VGND.n10 VGND.n8 0.119
R73 VNB VNB.t2 6502.94
R74 VNB.t4 VNB.t3 5246.15
R75 VNB.t3 VNB.t0 4796.06
R76 VNB.t0 VNB.t1 2782.35
R77 VNB.t2 VNB.t4 2714.84
R78 a_228_47.n0 a_228_47.t2 250.639
R79 a_228_47.t1 a_228_47.n1 237.798
R80 a_228_47.n1 a_228_47.t0 173.328
R81 a_228_47.n0 a_228_47.t3 149.419
R82 a_228_47.n1 a_228_47.n0 66.055
C0 X VGND 0.20fF
C1 VPWR VGND 0.11fF
C2 VPWR X 0.30fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__clkdlybuf4s18_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__clkdlybuf4s18_1 VPWR VGND A X VNB VPB
X0 VPWR.t0 A.t0 a_27_47.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 X.t0 a_394_47.t2 VGND.t3 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 VGND.t2 a_282_47.t2 a_394_47.t0 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=180000u
X3 X.t1 a_394_47.t3 VPWR.t3 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 a_282_47.t1 a_27_47.t2 VPWR.t1 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=820000u l=180000u
X5 VGND.t0 A.t1 a_27_47.t1 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 a_282_47.t0 a_27_47.t3 VGND.t1 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=180000u
X7 VPWR.t2 a_282_47.t3 a_394_47.t1 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=820000u l=180000u
R0 A.n0 A.t0 227.415
R1 A.n0 A.t1 206.091
R2 A A.n0 87.377
R3 a_27_47.t0 a_27_47.n1 225.06
R4 a_27_47.n0 a_27_47.t2 187.443
R5 a_27_47.n1 a_27_47.t1 180.31
R6 a_27_47.n1 a_27_47.n0 130.397
R7 a_27_47.n0 a_27_47.t3 124.515
R8 VPWR.n2 VPWR.n0 169.792
R9 VPWR.n2 VPWR.n1 168.21
R10 VPWR.n1 VPWR.t1 112.267
R11 VPWR.n0 VPWR.t2 108.627
R12 VPWR.n1 VPWR.t0 36.856
R13 VPWR.n0 VPWR.t3 36.263
R14 VPWR VPWR.n2 0.151
R15 VPB.t1 VPB.t2 594.859
R16 VPB.t2 VPB.t3 500.155
R17 VPB.t0 VPB.t1 500.155
R18 VPB VPB.t0 195.327
R19 a_394_47.t1 a_394_47.n1 258.74
R20 a_394_47.n1 a_394_47.t0 248.651
R21 a_394_47.n0 a_394_47.t3 227.415
R22 a_394_47.n0 a_394_47.t2 205.214
R23 a_394_47.n1 a_394_47.n0 76
R24 VGND.n2 VGND.n1 111.347
R25 VGND.n2 VGND.n0 111.121
R26 VGND.n1 VGND.t1 89.538
R27 VGND.n0 VGND.t2 84.923
R28 VGND.n0 VGND.t3 51.735
R29 VGND.n1 VGND.t0 47.12
R30 VGND VGND.n2 0.15
R31 X.n1 X.t1 174
R32 X X.t0 134.015
R33 X X.n0 12.515
R34 X.n1 X 8.94
R35 X.n0 X 6.826
R36 X.n0 X 4.042
R37 X X.n1 2.771
R38 VNB VNB.t0 6502.94
R39 VNB.t1 VNB.t2 4859.34
R40 VNB.t2 VNB.t3 3971.98
R41 VNB.t0 VNB.t1 3971.98
R42 a_282_47.t1 a_282_47.n1 231.386
R43 a_282_47.n0 a_282_47.t3 201.836
R44 a_282_47.n0 a_282_47.t2 132.549
R45 a_282_47.n1 a_282_47.t0 108.239
R46 a_282_47.n1 a_282_47.n0 76.014
C0 X VPWR 0.14fF
C1 X VGND 0.12fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__clkdlybuf4s18_2.ext - technology: sky130A

.subckt sky130_fd_sc_hd__clkdlybuf4s18_2 A X VGND VPWR VNB VPB
X0 a_227_47.t0 a_27_47.t2 VGND.t4 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=180000u
X1 VGND.t1 a_334_47.t2 X.t1 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 VGND.t0 a_227_47.t2 a_334_47.t0 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=180000u
X3 VPWR.t0 a_227_47.t3 a_334_47.t1 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=820000u l=180000u
X4 VPWR.t3 A.t0 a_27_47.t0 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 X.t0 a_334_47.t3 VGND.t2 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 VGND.t3 A.t1 a_27_47.t1 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7 X.t3 a_334_47.t4 VPWR.t2 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 a_227_47.t1 a_27_47.t3 VPWR.t4 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=820000u l=180000u
X9 VPWR.t1 a_334_47.t5 X.t2 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
R0 a_27_47.t0 a_27_47.n1 230.252
R1 a_27_47.n0 a_27_47.t3 228.583
R2 a_27_47.n1 a_27_47.t1 184.54
R3 a_27_47.n0 a_27_47.t2 144.233
R4 a_27_47.n1 a_27_47.n0 76
R5 VGND.n2 VGND.t1 184.019
R6 VGND.n10 VGND.n9 108.015
R7 VGND.n1 VGND.n0 106.337
R8 VGND.n0 VGND.t2 71.428
R9 VGND.n9 VGND.t3 55.714
R10 VGND.n0 VGND.t0 44.571
R11 VGND.n9 VGND.t4 43.911
R12 VGND.n4 VGND.n3 4.65
R13 VGND.n6 VGND.n5 4.65
R14 VGND.n8 VGND.n7 4.65
R15 VGND.n2 VGND.n1 4.065
R16 VGND.n11 VGND.n10 4.037
R17 VGND.n4 VGND.n2 0.202
R18 VGND.n11 VGND.n8 0.135
R19 VGND VGND.n11 0.124
R20 VGND.n6 VGND.n4 0.119
R21 VGND.n8 VGND.n6 0.119
R22 a_227_47.t1 a_227_47.n1 230.545
R23 a_227_47.n0 a_227_47.t3 208.865
R24 a_227_47.n1 a_227_47.t0 161.652
R25 a_227_47.n0 a_227_47.t2 124.515
R26 a_227_47.n1 a_227_47.n0 82.727
R27 VNB VNB.t3 6502.94
R28 VNB.t4 VNB.t0 4738.46
R29 VNB.t0 VNB.t2 3032.47
R30 VNB.t2 VNB.t1 2782.35
R31 VNB.t3 VNB.t4 2618.14
R32 a_334_47.t1 a_334_47.n3 253.235
R33 a_334_47.n0 a_334_47.t5 221.719
R34 a_334_47.n1 a_334_47.t4 221.719
R35 a_334_47.n0 a_334_47.t2 186.373
R36 a_334_47.n1 a_334_47.t3 186.373
R37 a_334_47.n3 a_334_47.t0 183.726
R38 a_334_47.n3 a_334_47.n2 92.188
R39 a_334_47.n2 a_334_47.n0 74.977
R40 a_334_47.n2 a_334_47.n1 1.785
R41 X.n1 X.n0 146.395
R42 X.n3 X.n2 92.5
R43 X X.n3 88.933
R44 X.n2 X.t1 40
R45 X.n2 X.t0 40
R46 X.n0 X.t2 27.58
R47 X.n0 X.t3 27.58
R48 X X.n1 7.611
R49 X.n1 X 2.357
R50 X.n3 X 0.287
R51 VPWR.n2 VPWR.t1 219.843
R52 VPWR.n10 VPWR.n9 165.571
R53 VPWR.n1 VPWR.n0 161.626
R54 VPWR.n0 VPWR.t0 56.457
R55 VPWR.n0 VPWR.t2 54.462
R56 VPWR.n9 VPWR.t3 47.254
R57 VPWR.n9 VPWR.t4 45.646
R58 VPWR.n4 VPWR.n3 4.65
R59 VPWR.n6 VPWR.n5 4.65
R60 VPWR.n8 VPWR.n7 4.65
R61 VPWR.n11 VPWR.n10 4.056
R62 VPWR.n2 VPWR.n1 4.055
R63 VPWR.n4 VPWR.n2 0.204
R64 VPWR.n11 VPWR.n8 0.134
R65 VPWR VPWR.n11 0.124
R66 VPWR.n6 VPWR.n4 0.119
R67 VPWR.n8 VPWR.n6 0.119
R68 VPB.t4 VPB.t0 580.062
R69 VPB.t0 VPB.t2 378.816
R70 VPB.t3 VPB.t4 334.423
R71 VPB.t2 VPB.t1 254.517
R72 VPB VPB.t3 195.327
R73 A.n0 A.t0 240.01
R74 A.n0 A.t1 204.664
R75 A A.n0 90.586
C0 X VGND 0.18fF
C1 VPWR X 0.33fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__clkdlybuf4s25_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__clkdlybuf4s25_1 A X VPWR VGND VNB VPB
X0 a_244_47.t1 a_27_47.t2 VPWR.t1 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=820000u l=250000u
X1 VPWR.t0 a_244_47.t2 a_355_47.t1 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=820000u l=250000u
X2 X.t1 a_355_47.t2 VPWR.t3 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 VPWR.t2 A.t0 a_27_47.t0 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 VGND.t0 A.t1 a_27_47.t1 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 VGND.t2 a_244_47.t3 a_355_47.t0 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=250000u
X6 X.t0 a_355_47.t3 VGND.t3 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7 a_244_47.t0 a_27_47.t3 VGND.t1 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=250000u
R0 a_27_47.t0 a_27_47.n1 224.619
R1 a_27_47.n1 a_27_47.t1 179.134
R2 a_27_47.n0 a_27_47.t2 165.006
R3 a_27_47.n0 a_27_47.t3 104.274
R4 a_27_47.n1 a_27_47.n0 76
R5 VPWR.n2 VPWR.n1 168.067
R6 VPWR.n2 VPWR.n0 159.449
R7 VPWR.n0 VPWR.t0 93.695
R8 VPWR.n1 VPWR.t1 50.451
R9 VPWR.n0 VPWR.t3 49.657
R10 VPWR.n1 VPWR.t2 46.053
R11 VPWR VPWR.n2 0.15
R12 a_244_47.t1 a_244_47.n1 227.592
R13 a_244_47.n1 a_244_47.t0 193.434
R14 a_244_47.n0 a_244_47.t2 150.384
R15 a_244_47.n0 a_244_47.t3 89.652
R16 a_244_47.n1 a_244_47.n0 85.708
R17 VPB.t0 VPB.t1 633.333
R18 VPB.t1 VPB.t3 479.439
R19 VPB.t2 VPB.t0 364.018
R20 VPB VPB.t2 195.327
R21 a_355_47.t1 a_355_47.n1 267.314
R22 a_355_47.n0 a_355_47.t2 241.534
R23 a_355_47.n0 a_355_47.t3 206.188
R24 a_355_47.n1 a_355_47.t0 196.313
R25 a_355_47.n1 a_355_47.n0 76
R26 X.n0 X.t1 173.887
R27 X X.t0 133.051
R28 X X.n0 5.861
R29 X.n1 X 5.028
R30 X X.n1 4.208
R31 X.n1 X 2.742
R32 X.n0 X 1.887
R33 A.n0 A.t0 235.978
R34 A.n0 A.t1 200.632
R35 A A.n0 84.881
R36 VGND.n2 VGND.n0 111.407
R37 VGND.n2 VGND.n1 97.917
R38 VGND.n1 VGND.t2 72
R39 VGND.n0 VGND.t0 54.285
R40 VGND.n1 VGND.t3 51.735
R41 VGND.n0 VGND.t1 48.615
R42 VGND VGND.n2 0.148
R43 VNB VNB.t0 6502.94
R44 VNB.t1 VNB.t2 5173.63
R45 VNB.t2 VNB.t3 3802.75
R46 VNB.t0 VNB.t1 2870.23
C0 X VGND 0.16fF
C1 X VPWR 0.16fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__clkdlybuf4s25_2.ext - technology: sky130A

.subckt sky130_fd_sc_hd__clkdlybuf4s25_2 X A VPWR VGND VNB VPB
X0 X.t3 a_331_47.t2 VGND.t4 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1 VPWR.t1 A.t0 a_27_47.t0 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 VGND.t0 a_225_47.t2 a_331_47.t0 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=250000u
X3 VPWR.t3 a_331_47.t3 X.t1 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 VGND.t1 A.t1 a_27_47.t1 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 VPWR.t0 a_225_47.t3 a_331_47.t1 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=820000u l=250000u
X6 a_225_47.t0 a_27_47.t2 VGND.t2 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=250000u
X7 X.t0 a_331_47.t4 VPWR.t2 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 a_225_47.t1 a_27_47.t3 VPWR.t4 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=820000u l=250000u
X9 VGND.t3 a_331_47.t5 X.t2 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
R0 a_331_47.t1 a_331_47.n2 298.082
R1 a_331_47.n2 a_331_47.t0 224.779
R2 a_331_47.n0 a_331_47.t3 207.259
R3 a_331_47.n1 a_331_47.t4 207.259
R4 a_331_47.n0 a_331_47.t5 173.52
R5 a_331_47.n1 a_331_47.t2 173.52
R6 a_331_47.n2 a_331_47.n1 83.467
R7 a_331_47.n1 a_331_47.n0 67.887
R8 VGND.n2 VGND.t3 171.46
R9 VGND.n10 VGND.n9 107.433
R10 VGND.n1 VGND.n0 107.239
R11 VGND.n0 VGND.t4 54.285
R12 VGND.n9 VGND.t1 54.285
R13 VGND.n0 VGND.t0 25.934
R14 VGND.n9 VGND.t2 25.934
R15 VGND.n2 VGND.n1 8.954
R16 VGND.n4 VGND.n3 4.65
R17 VGND.n6 VGND.n5 4.65
R18 VGND.n8 VGND.n7 4.65
R19 VGND.n11 VGND.n10 4.024
R20 VGND.n4 VGND.n2 0.211
R21 VGND.n11 VGND.n8 0.135
R22 VGND VGND.n11 0.125
R23 VGND.n6 VGND.n4 0.119
R24 VGND.n8 VGND.n6 0.119
R25 X.n3 X.n2 144.679
R26 X.n1 X.n0 92.5
R27 X.n0 X.t3 61.428
R28 X.n2 X.t0 42.355
R29 X.n0 X.t2 38.571
R30 X.n2 X.t1 26.595
R31 X X.n1 14.845
R32 X.n3 X 6.576
R33 X X.n3 6.526
R34 X.n1 X 0.984
R35 VNB VNB.t1 6502.94
R36 VNB.t2 VNB.t0 5028.57
R37 VNB.t4 VNB.t3 3235.29
R38 VNB.t0 VNB.t4 2497.1
R39 VNB.t1 VNB.t2 2497.1
R40 A.n0 A.t0 236.179
R41 A.n0 A.t1 196.451
R42 A.n1 A.n0 76
R43 A.n1 A 8.897
R44 A A.n1 1.717
R45 a_27_47.t0 a_27_47.n1 237.494
R46 a_27_47.n1 a_27_47.t1 195.609
R47 a_27_47.n0 a_27_47.t3 170.254
R48 a_27_47.n0 a_27_47.t2 109.522
R49 a_27_47.n1 a_27_47.n0 76
R50 VPWR.n10 VPWR.n9 307.239
R51 VPWR.n2 VPWR.t3 210.944
R52 VPWR.n1 VPWR.n0 164.214
R53 VPWR.n0 VPWR.t2 42.449
R54 VPWR.n9 VPWR.t1 42.449
R55 VPWR.n0 VPWR.t0 32.432
R56 VPWR.n9 VPWR.t4 32.432
R57 VPWR.n2 VPWR.n1 8.954
R58 VPWR.n4 VPWR.n3 4.65
R59 VPWR.n6 VPWR.n5 4.65
R60 VPWR.n8 VPWR.n7 4.65
R61 VPWR.n11 VPWR.n10 4.024
R62 VPWR.n4 VPWR.n2 0.212
R63 VPWR.n11 VPWR.n8 0.135
R64 VPWR VPWR.n11 0.125
R65 VPWR.n6 VPWR.n4 0.119
R66 VPWR.n8 VPWR.n6 0.119
R67 VPB.t4 VPB.t0 615.576
R68 VPB.t0 VPB.t2 310.747
R69 VPB.t1 VPB.t4 310.747
R70 VPB.t2 VPB.t3 295.95
R71 VPB VPB.t1 195.327
R72 a_225_47.t1 a_225_47.n1 269.016
R73 a_225_47.n0 a_225_47.t3 144.6
R74 a_225_47.n1 a_225_47.t0 140.403
R75 a_225_47.n0 a_225_47.t2 83.868
R76 a_225_47.n1 a_225_47.n0 67.726
C0 X VPWR 0.25fF
C1 X VGND 0.15fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__clkdlybuf4s50_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__clkdlybuf4s50_1 A X VGND VPWR VNB VPB
X0 a_283_47.t0 a_27_47.t2 VPWR.t3 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=820000u l=500000u
X1 VPWR.t0 A.t0 a_27_47.t0 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 VPWR.t1 a_283_47.t2 a_390_47.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=820000u l=500000u
X3 VGND.t0 a_283_47.t3 a_390_47.t1 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=500000u
X4 X.t0 a_390_47.t2 VPWR.t2 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 VGND.t1 A.t1 a_27_47.t1 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 a_283_47.t1 a_27_47.t3 VGND.t2 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=500000u
X7 X.t1 a_390_47.t3 VGND.t3 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
R0 a_27_47.t0 a_27_47.n1 227.285
R1 a_27_47.n1 a_27_47.t1 181.702
R2 a_27_47.n0 a_27_47.t2 88.206
R3 a_27_47.n1 a_27_47.n0 76
R4 a_27_47.n0 a_27_47.t3 57.84
R5 VPWR.n2 VPWR.n0 169.406
R6 VPWR.n2 VPWR.n1 168.942
R7 VPWR.n1 VPWR.t0 47.254
R8 VPWR.n0 VPWR.t2 41.248
R9 VPWR.n1 VPWR.t3 36.036
R10 VPWR.n0 VPWR.t1 33.634
R11 VPWR VPWR.n2 0.149
R12 a_283_47.t0 a_283_47.n1 211.09
R13 a_283_47.n1 a_283_47.t1 145.217
R14 a_283_47.n1 a_283_47.n0 118.656
R15 a_283_47.n0 a_283_47.t2 88.206
R16 a_283_47.n0 a_283_47.t3 57.84
R17 VPB.t3 VPB.t0 769.47
R18 VPB.t1 VPB.t3 405.451
R19 VPB.t0 VPB.t2 384.735
R20 VPB VPB.t1 195.327
R21 A.n0 A.t0 237.556
R22 A.n0 A.t1 203.128
R23 A A.n0 89.097
R24 a_390_47.n0 a_390_47.t2 241.534
R25 a_390_47.t0 a_390_47.n1 235.568
R26 a_390_47.n0 a_390_47.t3 206.188
R27 a_390_47.n1 a_390_47.t1 164.154
R28 a_390_47.n1 a_390_47.n0 98.496
R29 VGND.n2 VGND.n0 113.206
R30 VGND.n2 VGND.n1 112.76
R31 VGND.n1 VGND.t1 55.714
R32 VGND.n0 VGND.t3 52.857
R33 VGND.n1 VGND.t2 34.505
R34 VGND.n0 VGND.t0 27.362
R35 VGND VGND.n2 0.148
R36 VNB VNB.t1 6502.94
R37 VNB.t2 VNB.t0 6285.71
R38 VNB.t1 VNB.t2 3198.35
R39 VNB.t0 VNB.t3 3101.5
R40 X.n0 X.t0 176.863
R41 X.n1 X.t1 136.785
R42 X X.n1 12.879
R43 X X.n0 8.09
R44 X.n0 X 2.609
R45 X.n1 X 0.316
C0 X VGND 0.13fF
C1 VPWR X 0.13fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__clkdlybuf4s50_2.ext - technology: sky130A

.subckt sky130_fd_sc_hd__clkdlybuf4s50_2 A X VGND VPWR VNB VPB
X0 VPWR.t4 a_283_47.t2 a_390_47.t1 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=820000u l=500000u
X1 a_283_47.t1 a_27_47.t2 VPWR.t3 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=820000u l=500000u
X2 VPWR.t2 a_390_47.t2 X.t3 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 VPWR.t0 A.t0 a_27_47.t1 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 X.t2 a_390_47.t3 VPWR.t1 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 VGND.t4 a_283_47.t3 a_390_47.t0 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=500000u
X6 VGND.t3 A.t1 a_27_47.t0 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7 VGND.t2 a_390_47.t4 X.t1 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 a_283_47.t0 a_27_47.t3 VGND.t0 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=500000u
X9 X.t0 a_390_47.t5 VGND.t1 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
R0 a_283_47.t1 a_283_47.n1 228.87
R1 a_283_47.n1 a_283_47.t0 148.288
R2 a_283_47.n1 a_283_47.n0 120.01
R3 a_283_47.n0 a_283_47.t2 88.206
R4 a_283_47.n0 a_283_47.t3 57.84
R5 a_390_47.n1 a_390_47.t3 308.479
R6 a_390_47.n1 a_390_47.t5 273.133
R7 a_390_47.t1 a_390_47.n2 238.792
R8 a_390_47.n0 a_390_47.t2 221.719
R9 a_390_47.n0 a_390_47.t4 186.373
R10 a_390_47.n2 a_390_47.t0 166.589
R11 a_390_47.n2 a_390_47.n1 95.2
R12 a_390_47.n1 a_390_47.n0 86.581
R13 VPWR.n2 VPWR.t2 227.105
R14 VPWR.n1 VPWR.n0 165.571
R15 VPWR.n12 VPWR.n11 165.571
R16 VPWR.n11 VPWR.t0 47.254
R17 VPWR.n0 VPWR.t1 42.449
R18 VPWR.n11 VPWR.t3 36.036
R19 VPWR.n0 VPWR.t4 33.634
R20 VPWR.n4 VPWR.n3 4.65
R21 VPWR.n6 VPWR.n5 4.65
R22 VPWR.n8 VPWR.n7 4.65
R23 VPWR.n10 VPWR.n9 4.65
R24 VPWR.n13 VPWR.n12 4.056
R25 VPWR.n2 VPWR.n1 4.047
R26 VPWR.n4 VPWR.n2 0.203
R27 VPWR.n13 VPWR.n10 0.134
R28 VPWR VPWR.n13 0.124
R29 VPWR.n6 VPWR.n4 0.119
R30 VPWR.n8 VPWR.n6 0.119
R31 VPWR.n10 VPWR.n8 0.119
R32 VPB.t3 VPB.t4 766.51
R33 VPB.t0 VPB.t3 405.451
R34 VPB.t4 VPB.t1 387.694
R35 VPB.t1 VPB.t2 251.557
R36 VPB VPB.t0 195.327
R37 a_27_47.t1 a_27_47.n1 234.987
R38 a_27_47.n1 a_27_47.t0 189.188
R39 a_27_47.n0 a_27_47.t2 88.206
R40 a_27_47.n0 a_27_47.t3 57.84
R41 a_27_47.n1 a_27_47.n0 38
R42 X.n1 X.n0 146.322
R43 X.n4 X.n3 92.5
R44 X.n3 X.t0 40
R45 X.n3 X.t1 38.571
R46 X.n0 X.t2 27.58
R47 X.n0 X.t3 26.595
R48 X X.n4 10.659
R49 X X.n1 7.451
R50 X.n2 X 7.418
R51 X X.n2 3.885
R52 X.n2 X 2.472
R53 X.n1 X 2.402
R54 X.n4 X 1.309
R55 A.n0 A.t0 235.762
R56 A.n0 A.t1 200.416
R57 A A.n0 86.057
R58 VGND.n2 VGND.t2 195.503
R59 VGND.n12 VGND.n11 108.984
R60 VGND.n1 VGND.n0 108.015
R61 VGND.n11 VGND.t3 55.714
R62 VGND.n0 VGND.t1 54.285
R63 VGND.n11 VGND.t0 34.505
R64 VGND.n0 VGND.t4 27.362
R65 VGND.n4 VGND.n3 4.65
R66 VGND.n6 VGND.n5 4.65
R67 VGND.n8 VGND.n7 4.65
R68 VGND.n10 VGND.n9 4.65
R69 VGND.n2 VGND.n1 4.047
R70 VGND.n13 VGND.n12 4.037
R71 VGND.n4 VGND.n2 0.203
R72 VGND.n13 VGND.n10 0.135
R73 VGND VGND.n13 0.124
R74 VGND.n6 VGND.n4 0.119
R75 VGND.n8 VGND.n6 0.119
R76 VGND.n10 VGND.n8 0.119
R77 VNB VNB.t3 6502.94
R78 VNB.t0 VNB.t4 6261.54
R79 VNB.t3 VNB.t0 3198.35
R80 VNB.t4 VNB.t1 3115.34
R81 VNB.t1 VNB.t2 2750
C0 X VGND 0.17fF
C1 VPWR VGND 0.10fF
C2 VPWR X 0.25fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__clkinv_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__clkinv_1 Y A VGND VPWR VNB VPB
X0 Y.t2 A.t0 VPWR.t1 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X1 VGND.t0 A.t1 Y.t0 VNB sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 VPWR.t0 A.t2 Y.t1 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
R0 A.n0 A.t2 231.907
R1 A.n1 A.t0 231.36
R2 A A.n1 207.012
R3 A.n0 A.t1 170.306
R4 A.n1 A.n0 54.062
R5 VPWR.n0 VPWR.t1 271.758
R6 VPWR.n0 VPWR.t0 263.248
R7 VPWR VPWR.n0 0.126
R8 Y Y.n0 165.967
R9 Y Y.t0 143.953
R10 Y.n0 Y.t1 31.66
R11 Y.n0 Y.t2 31.66
R12 VPB.t1 VPB.t0 248.598
R13 VPB VPB.t1 192.367
R14 VGND VGND.t0 154.376
C0 Y VGND 0.15fF
C1 VPWR Y 0.35fF
C2 A Y 0.16fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__clkinv_2.ext - technology: sky130A

.subckt sky130_fd_sc_hd__clkinv_2 Y A VPWR VGND VNB VPB
X0 Y.t4 A.t0 VGND.t1 VNB sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1 Y.t2 A.t1 VPWR.t2 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 VPWR.t1 A.t2 Y.t1 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 VGND.t0 A.t3 Y.t3 VNB sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 VPWR.t0 A.t4 Y.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
R0 A.n0 A.t4 221.719
R1 A.n3 A.t1 221.719
R2 A.n7 A.t2 218.506
R3 A.n0 A.t3 189.05
R4 A.n2 A.t0 183.16
R5 A.n8 A.n7 105.086
R6 A.n6 A.n5 76
R7 A.n1 A.n0 63.278
R8 A.n6 A.n3 45.617
R9 A.n7 A.n6 27.957
R10 A.n5 A.n4 19.342
R11 A.n8 A 16.213
R12 A.n2 A.n1 10.328
R13 A A.n8 9.955
R14 A.n4 A 3.697
R15 A.n5 A 3.128
R16 A.n3 A.n2 2.582
R17 VGND.n0 VGND.t1 155.166
R18 VGND.n0 VGND.t0 150.198
R19 VGND VGND.n0 0.242
R20 Y.n2 Y.t1 289.254
R21 Y.n2 Y.n1 165.503
R22 Y.n3 Y.n0 130.205
R23 Y.n0 Y.t3 40
R24 Y.n0 Y.t4 40
R25 Y.n1 Y.t0 27.58
R26 Y.n1 Y.t2 27.58
R27 Y Y.n2 20.006
R28 Y.n3 Y 13.485
R29 Y Y.n3 2.057
R30 VPWR.n1 VPWR.t0 202.855
R31 VPWR.n1 VPWR.n0 174.156
R32 VPWR.n0 VPWR.t2 27.58
R33 VPWR.n0 VPWR.t1 27.58
R34 VPWR VPWR.n1 0.234
R35 VPB.t2 VPB.t0 254.517
R36 VPB.t1 VPB.t2 254.517
R37 VPB VPB.t1 207.165
C0 Y VGND 0.22fF
C1 Y VPWR 0.48fF
C2 Y A 0.28fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__clkinv_4.ext - technology: sky130A

.subckt sky130_fd_sc_hd__clkinv_4 A Y VPWR VGND VNB VPB
X0 Y.t7 A.t0 VPWR.t1 VPB.t5 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 VGND.t3 A.t1 Y.t1 VNB sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 VGND.t2 A.t2 Y.t0 VNB sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3 VPWR.t0 A.t3 Y.t6 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 VPWR.t5 A.t4 Y.t5 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 Y.t9 A.t5 VGND.t1 VNB sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 Y.t4 A.t6 VPWR.t4 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 Y.t8 A.t7 VGND.t0 VNB sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 Y.t3 A.t8 VPWR.t3 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 VPWR.t2 A.t9 Y.t2 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
R0 A.n0 A.t4 276.167
R1 A.n6 A.t6 247.604
R2 A.n2 A.t0 221.719
R3 A.n5 A.t9 221.719
R4 A.n13 A.t8 221.719
R5 A.n7 A.t3 221.719
R6 A.n2 A.t1 186.373
R7 A.n5 A.t5 186.373
R8 A.n13 A.t2 186.373
R9 A.n7 A.t7 186.373
R10 A.n1 A.n0 76
R11 A.n4 A.n3 76
R12 A.n15 A.n14 76
R13 A.n12 A.n11 76
R14 A.n10 A.n8 76
R15 A.n12 A.n8 60.696
R16 A.n14 A.n13 54.448
R17 A.n7 A.n6 50.877
R18 A.n3 A.n2 38.381
R19 A.n14 A.n5 22.314
R20 A.n4 A.n1 19.342
R21 A.n10 A.n9 19.342
R22 A A.n15 17.351
R23 A.n11 A 15.644
R24 A.n11 A 10.524
R25 A.n8 A.n7 9.818
R26 A.n15 A 8.817
R27 A.n13 A.n12 6.248
R28 A.n1 A 4.835
R29 A A.n10 3.697
R30 A.n9 A 3.128
R31 A A.n4 1.991
R32 VPWR.n2 VPWR.t5 194.268
R33 VPWR.n10 VPWR.t4 192.315
R34 VPWR.n6 VPWR.n5 170.749
R35 VPWR.n1 VPWR.n0 170.749
R36 VPWR.n5 VPWR.t3 27.58
R37 VPWR.n5 VPWR.t0 27.58
R38 VPWR.n0 VPWR.t1 27.58
R39 VPWR.n0 VPWR.t2 27.58
R40 VPWR.n4 VPWR.n3 4.65
R41 VPWR.n7 VPWR.n6 4.65
R42 VPWR.n9 VPWR.n8 4.65
R43 VPWR.n11 VPWR.n10 4.65
R44 VPWR.n2 VPWR.n1 3.948
R45 VPWR.n4 VPWR.n2 0.241
R46 VPWR.n7 VPWR.n4 0.119
R47 VPWR.n9 VPWR.n7 0.119
R48 VPWR.n11 VPWR.n9 0.119
R49 VPWR VPWR.n11 0.022
R50 Y.n5 Y.n4 165.877
R51 Y.n7 Y.n6 165.877
R52 Y.n9 Y.n8 165.503
R53 Y.n5 Y.n3 137.035
R54 Y.n1 Y.n0 110.821
R55 Y.n3 Y.n2 110.469
R56 Y.n10 Y.n1 51.952
R57 Y.n7 Y.n5 45.552
R58 Y.n3 Y.n1 45.176
R59 Y.n9 Y.n7 45.176
R60 Y.n0 Y.t1 40
R61 Y.n0 Y.t9 40
R62 Y.n2 Y.t0 40
R63 Y.n2 Y.t8 40
R64 Y.n4 Y.t6 27.58
R65 Y.n4 Y.t4 27.58
R66 Y.n6 Y.t2 27.58
R67 Y.n6 Y.t3 27.58
R68 Y.n8 Y.t5 27.58
R69 Y.n8 Y.t7 27.58
R70 Y Y.n9 23.466
R71 Y.n10 Y 12.586
R72 Y Y.n10 1.92
R73 VPB.t5 VPB.t3 254.517
R74 VPB.t0 VPB.t5 254.517
R75 VPB.t1 VPB.t0 254.517
R76 VPB.t4 VPB.t1 254.517
R77 VPB.t2 VPB.t4 254.517
R78 VPB VPB.t2 219.003
R79 VGND.n2 VGND.t3 152.681
R80 VGND.n5 VGND.t0 149.422
R81 VGND.n1 VGND.n0 111.7
R82 VGND.n0 VGND.t1 40
R83 VGND.n0 VGND.t2 40
R84 VGND.n4 VGND.n3 4.65
R85 VGND.n6 VGND.n5 4.01
R86 VGND.n2 VGND.n1 3.921
R87 VGND.n4 VGND.n2 0.23
R88 VGND.n6 VGND.n4 0.135
R89 VGND VGND.n6 0.125
C0 Y VGND 0.52fF
C1 VPWR Y 0.90fF
C2 A Y 1.20fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__clkinv_8.ext - technology: sky130A

.subckt sky130_fd_sc_hd__clkinv_8 Y A VGND VPWR VNB VPB
X0 Y.t16 A.t0 VGND.t3 VNB sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1 VPWR.t11 A.t1 Y.t19 VPB.t11 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 Y.t15 A.t2 VGND.t2 VNB sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3 Y.t14 A.t3 VGND.t1 VNB sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 Y.t8 A.t4 VPWR.t10 VPB.t10 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 VPWR.t9 A.t5 Y.t7 VPB.t9 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 VPWR.t8 A.t6 Y.t6 VPB.t8 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 Y.t13 A.t7 VGND.t0 VNB sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 Y.t5 A.t8 VPWR.t7 VPB.t7 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 VGND.t7 A.t9 Y.t12 VNB sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10 Y.t4 A.t10 VPWR.t6 VPB.t6 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 VPWR.t5 A.t11 Y.t3 VPB.t5 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 VGND.t6 A.t12 Y.t11 VNB sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13 VPWR.t4 A.t13 Y.t2 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14 Y.t1 A.t14 VPWR.t3 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 VGND.t5 A.t15 Y.t10 VNB sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16 VPWR.t2 A.t16 Y.t0 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17 Y.t18 A.t17 VPWR.t1 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X18 Y.t17 A.t18 VPWR.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X19 VGND.t4 A.t19 Y.t9 VNB sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
R0 A.n5 A.t11 225.91
R1 A.n41 A.t18 205.372
R2 A.n6 A.t8 192.799
R3 A.n4 A.t13 192.799
R4 A.n13 A.t14 192.799
R5 A.n15 A.t16 192.799
R6 A.n22 A.t17 192.799
R7 A.n2 A.t1 192.799
R8 A.n29 A.t4 192.799
R9 A.n32 A.t6 192.799
R10 A.n0 A.t10 192.799
R11 A.n40 A.t5 192.799
R12 A.n33 A.t0 117.286
R13 A.n31 A.t15 117.286
R14 A.n28 A.t7 117.286
R15 A.n23 A.t12 117.286
R16 A.n3 A.t3 117.286
R17 A.n16 A.t9 117.286
R18 A.n12 A.t2 117.286
R19 A.n7 A.t19 117.286
R20 A.n9 A.n8 76
R21 A.n11 A.n10 76
R22 A.n18 A.n17 76
R23 A.n21 A.n20 76
R24 A.n25 A.n24 76
R25 A.n27 A.n26 76
R26 A.n35 A.n34 76
R27 A.n37 A.n36 76
R28 A.n39 A.n38 76
R29 A.n42 A.n41 76
R30 A.n38 A.n37 28.5
R31 A.n23 A.n22 24.309
R32 A.n41 A.n40 22.633
R33 A.n27 A.n2 21.375
R34 A.n7 A.n6 20.956
R35 A.n11 A.n4 19.699
R36 A.n34 A.n33 18.86
R37 A.n14 A.n3 17.184
R38 A.n20 A.n19 17.066
R39 A.n35 A.n1 17.066
R40 A.n42 A.n39 17.066
R41 A.n26 A 16.564
R42 A A.n18 15.56
R43 A.n30 A.n29 14.669
R44 A.n10 A 13.552
R45 A.n13 A.n12 13.412
R46 A.n17 A.n13 12.993
R47 A.n16 A.n15 12.573
R48 A.n25 A 12.549
R49 A.n36 A 11.545
R50 A.n36 A 11.545
R51 A.n21 A.n3 11.316
R52 A.n31 A.n30 11.316
R53 A A.n25 10.541
R54 A.n29 A.n28 10.059
R55 A.n17 A.n16 9.64
R56 A.n10 A 9.537
R57 A.n32 A.n31 9.22
R58 A.n8 A.n4 8.801
R59 A.n33 A.n0 8.382
R60 A.n34 A.n32 7.963
R61 A.n18 A 7.529
R62 A.n24 A.n2 7.125
R63 A.n26 A 6.525
R64 A.n15 A.n14 6.286
R65 A A.n35 5.521
R66 A.n39 A 5.521
R67 A.n8 A.n7 5.448
R68 A.n20 A 4.517
R69 A.n24 A.n23 3.772
R70 A.n28 A.n27 3.772
R71 A A.n9 3.513
R72 A.n6 A.n5 2.095
R73 A.n12 A.n11 2.095
R74 A.n19 A 1.505
R75 A.n37 A.n0 1.257
R76 A A.n1 0.501
R77 A A.n42 0.501
R78 A.n22 A.n21 0.419
R79 VGND.n3 VGND.t4 151.62
R80 VGND.n0 VGND.t3 147.627
R81 VGND.n2 VGND.n1 107.627
R82 VGND.n7 VGND.n6 107.627
R83 VGND.n12 VGND.n11 107.627
R84 VGND.n1 VGND.t2 40
R85 VGND.n1 VGND.t7 40
R86 VGND.n6 VGND.t1 40
R87 VGND.n6 VGND.t6 40
R88 VGND.n11 VGND.t0 40
R89 VGND.n11 VGND.t5 40
R90 VGND.n5 VGND.n4 4.65
R91 VGND.n8 VGND.n7 4.65
R92 VGND.n10 VGND.n9 4.65
R93 VGND.n13 VGND.n12 4.65
R94 VGND.n15 VGND.n14 4.65
R95 VGND.n16 VGND.n0 4.013
R96 VGND.n3 VGND.n2 3.923
R97 VGND.n5 VGND.n3 0.31
R98 VGND VGND.n16 0.241
R99 VGND.n16 VGND.n15 0.137
R100 VGND.n8 VGND.n5 0.119
R101 VGND.n10 VGND.n8 0.119
R102 VGND.n13 VGND.n10 0.119
R103 VGND.n15 VGND.n13 0.119
R104 Y.n9 Y.n7 172.799
R105 Y.n9 Y.n8 171.181
R106 Y.n11 Y.n10 167.091
R107 Y.n19 Y.n18 167.091
R108 Y.n15 Y.n14 166.669
R109 Y.n13 Y.n12 166.266
R110 Y.n17 Y.n16 165.877
R111 Y.n1 Y.n0 115.068
R112 Y.n3 Y.n2 115.068
R113 Y.n5 Y.n4 115.068
R114 Y.n7 Y.n6 115.068
R115 Y.n20 Y.n1 65.129
R116 Y.n3 Y.n1 50.447
R117 Y.n5 Y.n3 50.447
R118 Y.n7 Y.n5 50.447
R119 Y.n11 Y.n9 45.176
R120 Y.n13 Y.n11 45.176
R121 Y.n17 Y.n15 44.8
R122 Y.n19 Y.n17 44.423
R123 Y.n15 Y.n13 44.047
R124 Y.n0 Y.t9 40
R125 Y.n0 Y.t15 40
R126 Y.n2 Y.t12 40
R127 Y.n2 Y.t14 40
R128 Y.n4 Y.t11 40
R129 Y.n4 Y.t13 40
R130 Y.n6 Y.t10 40
R131 Y.n6 Y.t16 40
R132 Y.n8 Y.t7 26.595
R133 Y.n8 Y.t17 26.595
R134 Y.n10 Y.t6 26.595
R135 Y.n10 Y.t4 26.595
R136 Y.n12 Y.t19 26.595
R137 Y.n12 Y.t8 26.595
R138 Y.n14 Y.t0 26.595
R139 Y.n14 Y.t18 26.595
R140 Y.n16 Y.t2 26.595
R141 Y.n16 Y.t1 26.595
R142 Y.n18 Y.t3 26.595
R143 Y.n18 Y.t5 26.595
R144 Y Y.n19 17.163
R145 Y.n20 Y 15.407
R146 Y Y.n20 0.711
R147 VPWR.n2 VPWR.t5 201.444
R148 VPWR.n25 VPWR.t0 197.344
R149 VPWR.n10 VPWR.n9 172.242
R150 VPWR.n1 VPWR.n0 171.725
R151 VPWR.n6 VPWR.n5 171.228
R152 VPWR.n21 VPWR.n20 170.749
R153 VPWR.n16 VPWR.n15 170.749
R154 VPWR.n20 VPWR.t9 27.58
R155 VPWR.n20 VPWR.t6 26.595
R156 VPWR.n15 VPWR.t10 26.595
R157 VPWR.n15 VPWR.t8 26.595
R158 VPWR.n9 VPWR.t1 26.595
R159 VPWR.n9 VPWR.t11 26.595
R160 VPWR.n5 VPWR.t3 26.595
R161 VPWR.n5 VPWR.t2 26.595
R162 VPWR.n0 VPWR.t7 26.595
R163 VPWR.n0 VPWR.t4 26.595
R164 VPWR.n11 VPWR.n10 6.023
R165 VPWR.n4 VPWR.n3 4.65
R166 VPWR.n8 VPWR.n7 4.65
R167 VPWR.n12 VPWR.n11 4.65
R168 VPWR.n14 VPWR.n13 4.65
R169 VPWR.n17 VPWR.n16 4.65
R170 VPWR.n19 VPWR.n18 4.65
R171 VPWR.n22 VPWR.n21 4.65
R172 VPWR.n24 VPWR.n23 4.65
R173 VPWR.n26 VPWR.n25 4.65
R174 VPWR.n2 VPWR.n1 3.716
R175 VPWR.n7 VPWR.n6 3.388
R176 VPWR.n4 VPWR.n2 0.237
R177 VPWR.n8 VPWR.n4 0.119
R178 VPWR.n12 VPWR.n8 0.119
R179 VPWR.n14 VPWR.n12 0.119
R180 VPWR.n17 VPWR.n14 0.119
R181 VPWR.n19 VPWR.n17 0.119
R182 VPWR.n22 VPWR.n19 0.119
R183 VPWR.n24 VPWR.n22 0.119
R184 VPWR.n26 VPWR.n24 0.119
R185 VPWR VPWR.n26 0.02
R186 VPB.t9 VPB.t6 251.557
R187 VPB.t7 VPB.t5 248.598
R188 VPB.t4 VPB.t7 248.598
R189 VPB.t3 VPB.t4 248.598
R190 VPB.t2 VPB.t3 248.598
R191 VPB.t1 VPB.t2 248.598
R192 VPB.t11 VPB.t1 248.598
R193 VPB.t10 VPB.t11 248.598
R194 VPB.t8 VPB.t10 248.598
R195 VPB.t6 VPB.t8 248.598
R196 VPB.t0 VPB.t9 248.598
R197 VPB VPB.t0 189.408
C0 VGND Y 0.93fF
C1 VGND VPWR 0.14fF
C2 VPWR Y 1.76fF
C3 A Y 2.37fF
C4 VPB VPWR 0.13fF
C5 VPB A 0.14fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__clkinv_16.ext - technology: sky130A

.subckt sky130_fd_sc_hd__clkinv_16 Y A VGND VPWR VNB VPB
X0 VGND.t15 A.t0 Y.t15 VNB sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1 Y.t29 A.t1 VPWR.t23 VPB.t23 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 VPWR.t22 A.t2 Y.t28 VPB.t22 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 Y.t27 A.t3 VPWR.t21 VPB.t21 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 VGND.t14 A.t4 Y.t14 VNB sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 VPWR.t20 A.t5 Y.t26 VPB.t20 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 Y.t13 A.t6 VGND.t13 VNB sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7 VGND.t12 A.t7 Y.t12 VNB sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 VPWR.t19 A.t8 Y.t25 VPB.t19 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 VPWR.t18 A.t9 Y.t8 VPB.t18 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 Y.t11 A.t10 VGND.t11 VNB sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11 Y.t7 A.t11 VPWR.t17 VPB.t17 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 VPWR.t16 A.t12 Y.t6 VPB.t16 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13 VGND.t10 A.t13 Y.t10 VNB sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14 Y.t5 A.t14 VPWR.t15 VPB.t15 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 VPWR.t14 A.t15 Y.t4 VPB.t14 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16 Y.t3 A.t16 VPWR.t13 VPB.t13 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17 Y.t2 A.t17 VPWR.t12 VPB.t12 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X18 Y.t9 A.t18 VGND.t9 VNB sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19 VGND.t8 A.t19 Y.t24 VNB sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20 Y.t23 A.t20 VGND.t7 VNB sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21 VGND.t6 A.t21 Y.t22 VNB sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22 Y.t1 A.t22 VPWR.t11 VPB.t11 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X23 VPWR.t10 A.t23 Y.t0 VPB.t10 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X24 Y.t39 A.t24 VPWR.t9 VPB.t9 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X25 Y.t38 A.t25 VPWR.t8 VPB.t8 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X26 VPWR.t7 A.t26 Y.t37 VPB.t7 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X27 Y.t21 A.t27 VGND.t5 VNB sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X28 Y.t36 A.t28 VPWR.t6 VPB.t6 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X29 VPWR.t5 A.t29 Y.t35 VPB.t5 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X30 VPWR.t4 A.t30 Y.t34 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X31 Y.t20 A.t31 VGND.t4 VNB sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X32 VGND.t3 A.t32 Y.t19 VNB sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X33 VPWR.t3 A.t33 Y.t33 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X34 Y.t18 A.t34 VGND.t2 VNB sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X35 Y.t32 A.t35 VPWR.t2 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X36 Y.t17 A.t36 VGND.t1 VNB sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X37 VPWR.t1 A.t37 Y.t31 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X38 Y.t30 A.t38 VPWR.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X39 VGND.t0 A.t39 Y.t16 VNB sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
R0 A.n3 A.t30 218.104
R1 A.n33 A.t14 218.104
R2 A.n4 A.t28 204.046
R3 A.n6 A.t29 204.046
R4 A.n26 A.t17 204.046
R5 A.n24 A.t5 204.046
R6 A.n23 A.t38 204.046
R7 A.n22 A.t26 204.046
R8 A.n21 A.t16 204.046
R9 A.n20 A.t15 204.046
R10 A.n19 A.t3 204.046
R11 A.n18 A.t37 204.046
R12 A.n17 A.t25 204.046
R13 A.n44 A.t12 204.046
R14 A.n45 A.t24 204.046
R15 A.n46 A.t2 204.046
R16 A.n47 A.t35 204.046
R17 A.n48 A.t23 204.046
R18 A.n49 A.t11 204.046
R19 A.n50 A.t9 204.046
R20 A.n51 A.t1 204.046
R21 A.n38 A.t33 204.046
R22 A.n40 A.t22 204.046
R23 A.n34 A.t8 204.046
R24 A.n24 A.t0 175.126
R25 A.n23 A.t10 175.126
R26 A.n22 A.t4 175.126
R27 A.n21 A.t18 175.126
R28 A.n20 A.t7 175.126
R29 A.n19 A.t20 175.126
R30 A.n18 A.t32 175.126
R31 A.n17 A.t27 175.126
R32 A.n44 A.t39 175.126
R33 A.n45 A.t34 175.126
R34 A.n46 A.t13 175.126
R35 A.n47 A.t6 175.126
R36 A.n48 A.t19 175.126
R37 A.n49 A.t31 175.126
R38 A.n50 A.t21 175.126
R39 A.n51 A.t36 175.126
R40 A.n36 A.n33 87.452
R41 A.n45 A.n44 78.325
R42 A.n36 A.n35 76
R43 A.n46 A.n45 62.258
R44 A.n24 A.n23 57.572
R45 A.n23 A.n22 57.572
R46 A.n22 A.n21 57.572
R47 A.n21 A.n20 57.572
R48 A.n20 A.n19 57.572
R49 A.n19 A.n18 57.572
R50 A.n18 A.n17 57.572
R51 A.n47 A.n46 57.572
R52 A.n48 A.n47 57.572
R53 A.n49 A.n48 57.572
R54 A.n50 A.n49 57.572
R55 A.n51 A.n50 57.572
R56 A.n4 A.n3 43.513
R57 A.n9 A.n5 38.158
R58 A.n41 A.n40 35.48
R59 A.n25 A.n24 34.141
R60 A.n54 A.n51 26.108
R61 A.n26 A.n25 23.43
R62 A.n41 A.n38 22.091
R63 A.n27 A.n26 21.422
R64 A.n42 A.n37 11.452
R65 A.n37 A.n36 11.452
R66 A.n16 A.n15 10.711
R67 A.n40 A.n39 10.041
R68 A.n10 A.n9 9.3
R69 A.n28 A.n27 9.3
R70 A.n55 A.n54 9.3
R71 A.n42 A.n41 8.286
R72 A.n54 A.n53 8.033
R73 A.n11 A.n0 7.806
R74 A.n9 A.n8 7.363
R75 A.n43 A.n32 6.435
R76 A.n7 A.n6 6.025
R77 A.n31 A.n30 4.65
R78 A.n8 A.n7 4.016
R79 A.n53 A.n52 3.347
R80 A.n43 A.n42 3.341
R81 A.n55 A.n43 3.33
R82 A.n14 A.n13 2.694
R83 A.n30 A.n29 2.694
R84 A.n12 A.n11 2.106
R85 A.n5 A.n4 2.008
R86 A.n35 A.n34 2.008
R87 A.n10 A.n2 1.852
R88 A.n11 A.n10 1.401
R89 A A.n57 1.178
R90 A.n2 A.n1 1.01
R91 A A.n55 0.842
R92 A.n57 A.n56 0.842
R93 A.n27 A.n16 0.669
R94 A.n28 A.n14 0.168
R95 A.n30 A.n28 0.168
R96 A.n32 A.n31 0.043
R97 A.n31 A.n12 0.002
R98 Y.n20 Y.n18 194.947
R99 Y.n10 Y.n8 158.161
R100 Y.n20 Y.n19 157.811
R101 Y.n3 Y.n2 157.157
R102 Y.n31 Y.n29 154.444
R103 Y.n5 Y.n4 154.376
R104 Y.n13 Y.n12 154.011
R105 Y.n22 Y.n21 153.778
R106 Y.n24 Y.n23 153.778
R107 Y.n26 Y.n25 153.778
R108 Y.n28 Y.n27 153.778
R109 Y.n7 Y.n6 147.682
R110 Y.n10 Y.n9 147.464
R111 Y.n3 Y.n1 146.381
R112 Y.n11 Y.n0 144.233
R113 Y.n28 Y.n14 142.164
R114 Y.n26 Y.n15 142.164
R115 Y.n24 Y.n16 142.164
R116 Y.n22 Y.n17 142.164
R117 Y Y.n30 128.998
R118 Y.n30 Y.t16 75.714
R119 Y.n29 Y.t39 53.19
R120 Y.n30 Y.t18 48.571
R121 Y.n24 Y.n22 44.032
R122 Y.n26 Y.n24 44.032
R123 Y.n28 Y.n26 44.032
R124 Y.n5 Y.n3 43.93
R125 Y.n22 Y.n20 43.58
R126 Y.n14 Y.t19 40
R127 Y.n14 Y.t21 40
R128 Y.n15 Y.t12 40
R129 Y.n15 Y.t23 40
R130 Y.n16 Y.t14 40
R131 Y.n16 Y.t9 40
R132 Y.n17 Y.t15 40
R133 Y.n17 Y.t11 40
R134 Y.n6 Y.t22 40
R135 Y.n6 Y.t17 40
R136 Y.n9 Y.t24 40
R137 Y.n9 Y.t20 40
R138 Y.n0 Y.t10 40
R139 Y.n0 Y.t13 40
R140 Y.n31 Y.n28 39.424
R141 Y.n31 Y.n13 39.29
R142 Y.n11 Y.n10 37.12
R143 Y.n10 Y.n7 36.864
R144 Y.n29 Y.t6 32.505
R145 Y.n27 Y.t31 27.58
R146 Y.n27 Y.t38 27.58
R147 Y.n25 Y.t4 27.58
R148 Y.n25 Y.t27 27.58
R149 Y.n23 Y.t37 27.58
R150 Y.n23 Y.t3 27.58
R151 Y.n21 Y.t26 27.58
R152 Y.n21 Y.t30 27.58
R153 Y.n18 Y.t34 27.58
R154 Y.n18 Y.t36 27.58
R155 Y.n19 Y.t35 27.58
R156 Y.n19 Y.t2 27.58
R157 Y.n1 Y.t25 27.58
R158 Y.n1 Y.t5 27.58
R159 Y.n2 Y.t33 27.58
R160 Y.n2 Y.t1 27.58
R161 Y.n4 Y.t8 27.58
R162 Y.n4 Y.t29 27.58
R163 Y.n8 Y.t0 27.58
R164 Y.n8 Y.t7 27.58
R165 Y.n12 Y.t28 27.58
R166 Y.n12 Y.t32 27.58
R167 Y Y.n31 3.84
R168 Y.n31 Y 3.242
R169 Y.n7 Y.n5 0.406
R170 Y.n13 Y.n11 0.135
R171 VGND.n1 VGND.t15 157.105
R172 VGND.n0 VGND.t1 153.596
R173 VGND.n13 VGND.n12 117.815
R174 VGND.n3 VGND.n2 113.994
R175 VGND.n9 VGND.n8 113.994
R176 VGND.n19 VGND.n18 113.994
R177 VGND.n26 VGND.n25 113.994
R178 VGND.n30 VGND.n29 113.994
R179 VGND.n36 VGND.n35 113.994
R180 VGND.n25 VGND.t10 47.142
R181 VGND.n25 VGND.t2 42.857
R182 VGND.n2 VGND.t11 40
R183 VGND.n2 VGND.t14 40
R184 VGND.n8 VGND.t9 40
R185 VGND.n8 VGND.t12 40
R186 VGND.n12 VGND.t7 40
R187 VGND.n12 VGND.t3 40
R188 VGND.n18 VGND.t5 40
R189 VGND.n18 VGND.t0 40
R190 VGND.n29 VGND.t13 40
R191 VGND.n29 VGND.t8 40
R192 VGND.n35 VGND.t4 40
R193 VGND.n35 VGND.t6 40
R194 VGND.n14 VGND.n13 7.152
R195 VGND.n27 VGND.n26 7.152
R196 VGND.n10 VGND.n9 6.023
R197 VGND.n31 VGND.n30 4.894
R198 VGND.n5 VGND.n4 4.65
R199 VGND.n7 VGND.n6 4.65
R200 VGND.n11 VGND.n10 4.65
R201 VGND.n15 VGND.n14 4.65
R202 VGND.n17 VGND.n16 4.65
R203 VGND.n20 VGND.n19 4.65
R204 VGND.n22 VGND.n21 4.65
R205 VGND.n24 VGND.n23 4.65
R206 VGND.n28 VGND.n27 4.65
R207 VGND.n32 VGND.n31 4.65
R208 VGND.n34 VGND.n33 4.65
R209 VGND.n38 VGND.n37 4.65
R210 VGND.n40 VGND.n39 4.65
R211 VGND.n41 VGND.n0 3.838
R212 VGND.n4 VGND.n3 1.505
R213 VGND.n5 VGND.n1 0.577
R214 VGND VGND.n41 0.477
R215 VGND.n37 VGND.n36 0.376
R216 VGND.n41 VGND.n40 0.142
R217 VGND.n7 VGND.n5 0.119
R218 VGND.n11 VGND.n7 0.119
R219 VGND.n15 VGND.n11 0.119
R220 VGND.n17 VGND.n15 0.119
R221 VGND.n20 VGND.n17 0.119
R222 VGND.n22 VGND.n20 0.119
R223 VGND.n24 VGND.n22 0.119
R224 VGND.n28 VGND.n24 0.119
R225 VGND.n32 VGND.n28 0.119
R226 VGND.n34 VGND.n32 0.119
R227 VGND.n38 VGND.n34 0.119
R228 VGND.n40 VGND.n38 0.119
R229 VPWR.n2 VPWR.t4 199.659
R230 VPWR.n50 VPWR.n49 169.471
R231 VPWR.n38 VPWR.n37 169.471
R232 VPWR.n34 VPWR.n33 169.471
R233 VPWR.n21 VPWR.n20 169.471
R234 VPWR.n17 VPWR.n16 169.471
R235 VPWR.n11 VPWR.n10 169.471
R236 VPWR.n6 VPWR.n5 169.471
R237 VPWR.n1 VPWR.n0 169.471
R238 VPWR.n27 VPWR.n26 169.053
R239 VPWR.n55 VPWR.n54 169.026
R240 VPWR.n44 VPWR.n43 169.026
R241 VPWR.n59 VPWR.t15 151.121
R242 VPWR.n33 VPWR.t22 31.52
R243 VPWR.n33 VPWR.t9 30.535
R244 VPWR.n26 VPWR.t8 28.565
R245 VPWR.n54 VPWR.t11 27.58
R246 VPWR.n54 VPWR.t19 27.58
R247 VPWR.n49 VPWR.t23 27.58
R248 VPWR.n49 VPWR.t3 27.58
R249 VPWR.n43 VPWR.t17 27.58
R250 VPWR.n43 VPWR.t18 27.58
R251 VPWR.n37 VPWR.t2 27.58
R252 VPWR.n37 VPWR.t10 27.58
R253 VPWR.n20 VPWR.t21 27.58
R254 VPWR.n20 VPWR.t1 27.58
R255 VPWR.n16 VPWR.t13 27.58
R256 VPWR.n16 VPWR.t14 27.58
R257 VPWR.n10 VPWR.t0 27.58
R258 VPWR.n10 VPWR.t7 27.58
R259 VPWR.n5 VPWR.t12 27.58
R260 VPWR.n5 VPWR.t20 27.58
R261 VPWR.n0 VPWR.t6 27.58
R262 VPWR.n0 VPWR.t5 27.58
R263 VPWR.n26 VPWR.t16 26.595
R264 VPWR.n35 VPWR.n34 7.152
R265 VPWR.n18 VPWR.n17 6.4
R266 VPWR.n39 VPWR.n38 5.27
R267 VPWR.n4 VPWR.n3 4.65
R268 VPWR.n7 VPWR.n6 4.65
R269 VPWR.n9 VPWR.n8 4.65
R270 VPWR.n13 VPWR.n12 4.65
R271 VPWR.n15 VPWR.n14 4.65
R272 VPWR.n19 VPWR.n18 4.65
R273 VPWR.n23 VPWR.n22 4.65
R274 VPWR.n25 VPWR.n24 4.65
R275 VPWR.n28 VPWR.n27 4.65
R276 VPWR.n30 VPWR.n29 4.65
R277 VPWR.n32 VPWR.n31 4.65
R278 VPWR.n36 VPWR.n35 4.65
R279 VPWR.n40 VPWR.n39 4.65
R280 VPWR.n42 VPWR.n41 4.65
R281 VPWR.n46 VPWR.n45 4.65
R282 VPWR.n48 VPWR.n47 4.65
R283 VPWR.n51 VPWR.n50 4.65
R284 VPWR.n53 VPWR.n52 4.65
R285 VPWR.n56 VPWR.n55 4.65
R286 VPWR.n58 VPWR.n57 4.65
R287 VPWR.n60 VPWR.n59 4.65
R288 VPWR.n22 VPWR.n21 4.517
R289 VPWR.n2 VPWR.n1 3.84
R290 VPWR.n12 VPWR.n11 1.882
R291 VPWR.n45 VPWR.n44 0.752
R292 VPWR.n4 VPWR.n2 0.24
R293 VPWR.n7 VPWR.n4 0.119
R294 VPWR.n9 VPWR.n7 0.119
R295 VPWR.n13 VPWR.n9 0.119
R296 VPWR.n15 VPWR.n13 0.119
R297 VPWR.n19 VPWR.n15 0.119
R298 VPWR.n23 VPWR.n19 0.119
R299 VPWR.n25 VPWR.n23 0.119
R300 VPWR.n28 VPWR.n25 0.119
R301 VPWR.n30 VPWR.n28 0.119
R302 VPWR.n32 VPWR.n30 0.119
R303 VPWR.n36 VPWR.n32 0.119
R304 VPWR.n40 VPWR.n36 0.119
R305 VPWR.n42 VPWR.n40 0.119
R306 VPWR.n46 VPWR.n42 0.119
R307 VPWR.n48 VPWR.n46 0.119
R308 VPWR.n51 VPWR.n48 0.119
R309 VPWR.n53 VPWR.n51 0.119
R310 VPWR.n56 VPWR.n53 0.119
R311 VPWR.n58 VPWR.n56 0.119
R312 VPWR.n60 VPWR.n58 0.119
R313 VPWR VPWR.n60 0.022
R314 VPB.t9 VPB.t16 346.261
R315 VPB.t22 VPB.t9 275.233
R316 VPB.t6 VPB.t4 254.517
R317 VPB.t5 VPB.t6 254.517
R318 VPB.t12 VPB.t5 254.517
R319 VPB.t20 VPB.t12 254.517
R320 VPB.t0 VPB.t20 254.517
R321 VPB.t7 VPB.t0 254.517
R322 VPB.t13 VPB.t7 254.517
R323 VPB.t14 VPB.t13 254.517
R324 VPB.t21 VPB.t14 254.517
R325 VPB.t1 VPB.t21 254.517
R326 VPB.t8 VPB.t1 254.517
R327 VPB.t16 VPB.t8 254.517
R328 VPB.t2 VPB.t22 254.517
R329 VPB.t10 VPB.t2 254.517
R330 VPB.t17 VPB.t10 254.517
R331 VPB.t18 VPB.t17 254.517
R332 VPB.t23 VPB.t18 254.517
R333 VPB.t3 VPB.t23 254.517
R334 VPB.t11 VPB.t3 254.517
R335 VPB.t19 VPB.t11 254.517
R336 VPB.t15 VPB.t19 254.517
R337 VPB VPB.t15 201.246
C0 VPWR Y 3.28fF
C1 A Y 0.96fF
C2 A VPWR 0.47fF
C3 VPB VPWR 0.22fF
C4 VPB A 0.32fF
C5 Y VGND 1.38fF
C6 VPWR VGND 0.12fF
C7 A VGND 0.71fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__clkinvlp_2.ext - technology: sky130A

.subckt sky130_fd_sc_hd__clkinvlp_2 VGND VPWR Y A VNB VPB
X0 Y.t2 A.t0 a_150_67.t0 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=550000u l=150000u
X1 VPWR.t1 A.t1 Y.t1 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=250000u
X2 a_150_67.t1 A.t2 VGND.t0 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=550000u l=150000u
X3 Y.t0 A.t3 VPWR.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=250000u
R0 A.n0 A.t1 189.265
R1 A.n2 A.t3 140.941
R2 A.n1 A.t2 130.163
R3 A.n0 A.t0 122.106
R4 A A.n2 83.068
R5 A.n1 A.n0 77.923
R6 A.n2 A.n1 6.072
R7 a_150_67.t0 a_150_67.t1 52.363
R8 Y Y.n0 167.649
R9 Y.n1 Y.t2 123.045
R10 Y.n0 Y.t1 27.58
R11 Y.n0 Y.t0 27.58
R12 Y Y.n1 3.877
R13 Y.n1 Y 3.124
R14 VNB VNB.t0 10770.2
R15 VNB.t0 VNB.t1 2118.52
R16 VPWR.n0 VPWR.t0 195.132
R17 VPWR.n0 VPWR.t1 178.059
R18 VPWR VPWR.n0 0.079
R19 VPB.t0 VPB.t1 313.707
R20 VPB VPB.t0 301.869
R21 VGND VGND.t0 150.24
C0 Y VGND 0.15fF
C1 VPWR Y 0.27fF
C2 A Y 0.10fF
C3 A VPWR 0.11fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__clkinvlp_4.ext - technology: sky130A

.subckt sky130_fd_sc_hd__clkinvlp_4 A Y VPWR VGND VNB VPB
X0 Y.t5 A.t0 VPWR.t3 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=250000u
X1 VGND.t0 A.t1 a_268_47.t0 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=550000u l=150000u
X2 Y.t4 A.t2 VPWR.t2 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=250000u
X3 Y.t1 A.t3 a_110_47.t1 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=550000u l=150000u
X4 VPWR.t1 A.t4 Y.t3 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=250000u
X5 a_110_47.t0 A.t5 VGND.t1 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=550000u l=150000u
X6 a_268_47.t1 A.t6 Y.t0 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=550000u l=150000u
X7 VPWR.t0 A.t7 Y.t2 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=250000u
R0 A.n0 A.t7 198.817
R1 A.n6 A.t5 155.846
R2 A.n4 A.t3 155.846
R3 A.n2 A.t6 155.846
R4 A.n0 A.t1 155.846
R5 A.n1 A.t2 127.248
R6 A.n3 A.t4 127.248
R7 A.n5 A.t0 127.248
R8 A A.n6 101.439
R9 A.n2 A.n1 46.739
R10 A.n5 A.n4 45.278
R11 A.n4 A.n3 32.133
R12 A.n3 A.n2 30.672
R13 A.n6 A.n5 7.303
R14 A.n1 A.n0 5.842
R15 VPWR.n0 VPWR.t0 150.756
R16 VPWR.n7 VPWR.t3 146.852
R17 VPWR.n2 VPWR.n1 119.569
R18 VPWR.n1 VPWR.t2 27.58
R19 VPWR.n1 VPWR.t1 27.58
R20 VPWR.n4 VPWR.n3 4.65
R21 VPWR.n6 VPWR.n5 4.65
R22 VPWR.n8 VPWR.n7 4.65
R23 VPWR.n3 VPWR.n2 0.376
R24 VPWR.n4 VPWR.n0 0.25
R25 VPWR.n6 VPWR.n4 0.119
R26 VPWR.n8 VPWR.n6 0.119
R27 VPWR VPWR.n8 0.022
R28 Y.n5 Y.n4 292.5
R29 Y.n3 Y.n0 156.625
R30 Y.n6 Y.n5 146.903
R31 Y.n2 Y.n1 95.361
R32 Y.n1 Y.t0 30.545
R33 Y.n1 Y.t1 30.545
R34 Y.n5 Y.t3 27.58
R35 Y.n5 Y.t5 27.58
R36 Y.n0 Y.t2 27.58
R37 Y.n0 Y.t4 27.58
R38 Y Y.n2 10.666
R39 Y Y.n3 10.311
R40 Y.n6 Y 9.547
R41 Y.n4 Y 6.577
R42 Y.n4 Y 5.511
R43 Y Y.n6 2.5
R44 Y.n3 Y 1.777
R45 Y.n2 Y 1.422
R46 VPB.t2 VPB.t0 313.707
R47 VPB.t1 VPB.t2 313.707
R48 VPB.t3 VPB.t1 313.707
R49 VPB VPB.t3 224.922
R50 a_268_47.t0 a_268_47.t1 45.818
R51 VGND.n0 VGND.t0 147.702
R52 VGND.n0 VGND.t1 143.599
R53 VGND VGND.n0 0.048
R54 VNB VNB.t1 6248.51
R55 VNB.t2 VNB.t0 2335.8
R56 VNB.t0 VNB.t3 1955.56
R57 VNB.t1 VNB.t2 1955.56
R58 a_110_47.t0 a_110_47.t1 45.818
C0 A VPWR 0.10fF
C1 Y VPWR 0.75fF
C2 Y A 0.16fF
C3 Y VGND 0.26fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__conb_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__conb_1 LO HI VPB VNB VGND VPWR
R0 HI VPWR sky130_fd_pr__res_generic_po w=480000u l=45000u
R1 VGND LO sky130_fd_pr__res_generic_po w=480000u l=45000u
C0 HI VGND 0.20fF
C1 HI LO 0.14fF
C2 VPWR LO 0.30fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__decap_3.ext - technology: sky130A

.subckt sky130_fd_sc_hd__decap_3 VPWR VGND VNB VPB
X0 VPWR.t1 VGND.t2 VPWR.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=870000u l=590000u
X1 VGND.t1 VPWR.t2 VGND.t0 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=550000u l=590000u
R0 VGND.n1 VGND.t2 183.08
R1 VGND.n0 VGND.t0 123.916
R2 VGND.n2 VGND.t1 121.954
R3 VGND.n3 VGND.n2 5.067
R4 VGND.n3 VGND.n0 1.644
R5 VGND.n2 VGND.n1 1.182
R6 VGND VGND.n3 0.022
R7 VPWR.n1 VPWR.t0 234.553
R8 VPWR.n4 VPWR.t1 234.553
R9 VPWR.n0 VPWR.t2 166.281
R10 VPWR.n3 VPWR.n1 5.073
R11 VPWR.n5 VPWR.n4 4.954
R12 VPWR.n3 VPWR.n2 4.65
R13 VPWR.n1 VPWR.n0 0.863
R14 VPWR.n5 VPWR.n3 0.119
R15 VPWR VPWR.n5 0.022
R16 VPB VPB.t0 315.767
R17 VNB VNB.t0 7416.41
C0 VGND VPWR 0.44fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__decap_4.ext - technology: sky130A

.subckt sky130_fd_sc_hd__decap_4 VGND VPWR VNB VPB
X0 VPWR.t1 VGND.t2 VPWR.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X1 VGND.t1 VPWR.t2 VGND.t0 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
R0 VGND.n0 VGND.t2 142.306
R1 VGND.n1 VGND.t0 124.813
R2 VGND.n2 VGND.t1 121.954
R3 VGND.n1 VGND.n0 5.732
R4 VGND.n3 VGND.n2 5.058
R5 VGND.n3 VGND.n1 0.657
R6 VGND VGND.n3 0.022
R7 VPWR.n0 VPWR.t0 242.133
R8 VPWR.n6 VPWR.t1 242.133
R9 VPWR.n1 VPWR.t2 134.961
R10 VPWR.n3 VPWR.n0 5.073
R11 VPWR.n7 VPWR.n6 4.954
R12 VPWR.n3 VPWR.n2 4.65
R13 VPWR.n5 VPWR.n4 4.65
R14 VPWR.n2 VPWR.n1 2.336
R15 VPWR.n5 VPWR.n3 0.119
R16 VPWR.n7 VPWR.n5 0.119
R17 VPWR VPWR.n7 0.022
R18 VPB VPB.t0 458.722
R19 VNB VNB.t0 8665.79
C0 VGND VPWR 0.67fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__decap_6.ext - technology: sky130A

.subckt sky130_fd_sc_hd__decap_6 VPWR VGND VNB VPB
X0 VPWR.t1 VGND.t2 VPWR.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.97e+06u
X1 VGND.t1 VPWR.t2 VGND.t0 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=550000u l=1.97e+06u
R0 VGND.n1 VGND.t0 125.217
R1 VGND.n0 VGND.t1 121.954
R2 VGND.n0 VGND.t2 83.894
R3 VGND.n1 VGND.n0 3.853
R4 VGND VGND.n1 0.465
R5 VPWR.n1 VPWR.t0 243.707
R6 VPWR.n8 VPWR.t1 242.133
R7 VPWR.n0 VPWR.t2 91.339
R8 VPWR.n9 VPWR.n8 4.954
R9 VPWR.n3 VPWR.n2 4.65
R10 VPWR.n5 VPWR.n4 4.65
R11 VPWR.n7 VPWR.n6 4.65
R12 VPWR.n3 VPWR.n1 1.794
R13 VPWR.n1 VPWR.n0 1.442
R14 VPWR.n5 VPWR.n3 0.119
R15 VPWR.n7 VPWR.n5 0.119
R16 VPWR.n9 VPWR.n7 0.119
R17 VPWR VPWR.n9 0.022
R18 VPB VPB.t0 730.996
R19 VNB VNB.t0 11164.6
C0 VGND VPWR 1.12fF
C1 VPB VPWR 0.10fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__decap_8.ext - technology: sky130A

.subckt sky130_fd_sc_hd__decap_8 VPWR VGND VNB VPB
X0 VPWR.t1 VGND.t2 VPWR.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=870000u l=2.89e+06u
X1 VGND.t1 VPWR.t2 VGND.t0 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=550000u l=2.89e+06u
R0 VGND.n1 VGND.t0 125.437
R1 VGND.n10 VGND.t1 121.954
R2 VGND.n4 VGND.n3 76
R3 VGND.n2 VGND.t2 34.296
R4 VGND.n11 VGND.n10 4.913
R5 VGND.n3 VGND.n2 4.857
R6 VGND.n6 VGND.n5 4.65
R7 VGND.n9 VGND.n8 4.65
R8 VGND.n1 VGND.n0 3.466
R9 VGND.n8 VGND.n7 1.139
R10 VGND.n5 VGND.n4 0.832
R11 VGND.n6 VGND.n1 0.235
R12 VGND.n9 VGND.n6 0.119
R13 VGND.n11 VGND.n9 0.119
R14 VGND VGND.n11 0.022
R15 VPWR.n18 VPWR.t1 242.133
R16 VPWR.n0 VPWR.t0 242.133
R17 VPWR.n6 VPWR.n5 76
R18 VPWR.n4 VPWR.t2 50.505
R19 VPWR.n5 VPWR.n4 7.118
R20 VPWR.n3 VPWR.n0 4.984
R21 VPWR.n19 VPWR.n18 4.954
R22 VPWR.n3 VPWR.n2 4.65
R23 VPWR.n8 VPWR.n7 4.65
R24 VPWR.n11 VPWR.n10 4.65
R25 VPWR.n13 VPWR.n12 4.65
R26 VPWR.n15 VPWR.n14 4.65
R27 VPWR.n17 VPWR.n16 4.65
R28 VPWR.n2 VPWR.n1 0.934
R29 VPWR.n7 VPWR.n6 0.539
R30 VPWR.n10 VPWR.n9 0.143
R31 VPWR.n8 VPWR.n3 0.119
R32 VPWR.n11 VPWR.n8 0.119
R33 VPWR.n13 VPWR.n11 0.119
R34 VPWR.n15 VPWR.n13 0.119
R35 VPWR.n17 VPWR.n15 0.119
R36 VPWR.n19 VPWR.n17 0.119
R37 VPWR VPWR.n19 0.022
R38 VPB VPB.t0 1003.27
R39 VNB VNB.t0 13663.3
C0 VPB VPWR 0.13fF
C1 VPB VGND 0.12fF
C2 VGND VPWR 1.57fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__decap_12.ext - technology: sky130A

.subckt sky130_fd_sc_hd__decap_12 VGND VPWR VNB VPB
X0 VPWR.t1 VGND.t2 VPWR.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=870000u l=4.73e+06u
X1 VGND.t1 VPWR.t2 VGND.t0 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=550000u l=4.73e+06u
R0 VGND.n2 VGND.t0 125.719
R1 VGND.n17 VGND.t1 121.954
R2 VGND.n1 VGND.n0 76
R3 VGND.n6 VGND.n5 76
R4 VGND.n11 VGND.n10 76
R5 VGND.n9 VGND.t2 68.698
R6 VGND.n10 VGND.n9 31.477
R7 VGND.n18 VGND.n17 4.913
R8 VGND.n4 VGND.n3 4.65
R9 VGND.n8 VGND.n7 4.65
R10 VGND.n13 VGND.n12 4.65
R11 VGND.n16 VGND.n15 4.65
R12 VGND.n2 VGND.n1 3.42
R13 VGND.n7 VGND.n6 2.016
R14 VGND.n15 VGND.n14 1.139
R15 VGND.n12 VGND.n11 0.438
R16 VGND.n4 VGND.n2 0.187
R17 VGND.n8 VGND.n4 0.119
R18 VGND.n13 VGND.n8 0.119
R19 VGND.n16 VGND.n13 0.119
R20 VGND.n18 VGND.n16 0.119
R21 VGND VGND.n18 0.022
R22 VPWR.n29 VPWR.t1 242.133
R23 VPWR.n0 VPWR.t0 242.133
R24 VPWR.n4 VPWR.t2 107.792
R25 VPWR.n16 VPWR.n15 76
R26 VPWR.n6 VPWR.n5 76
R27 VPWR.n12 VPWR.n11 76
R28 VPWR.n5 VPWR.n4 30.493
R29 VPWR.n3 VPWR.n0 4.984
R30 VPWR.n30 VPWR.n29 4.954
R31 VPWR.n3 VPWR.n2 4.65
R32 VPWR.n8 VPWR.n7 4.65
R33 VPWR.n10 VPWR.n9 4.65
R34 VPWR.n14 VPWR.n13 4.65
R35 VPWR.n18 VPWR.n17 4.65
R36 VPWR.n20 VPWR.n19 4.65
R37 VPWR.n22 VPWR.n21 4.65
R38 VPWR.n24 VPWR.n23 4.65
R39 VPWR.n26 VPWR.n25 4.65
R40 VPWR.n28 VPWR.n27 4.65
R41 VPWR.n13 VPWR.n12 1.51
R42 VPWR.n2 VPWR.n1 0.791
R43 VPWR.n7 VPWR.n6 0.503
R44 VPWR.n17 VPWR.n16 0.215
R45 VPWR.n8 VPWR.n3 0.119
R46 VPWR.n10 VPWR.n8 0.119
R47 VPWR.n14 VPWR.n10 0.119
R48 VPWR.n18 VPWR.n14 0.119
R49 VPWR.n20 VPWR.n18 0.119
R50 VPWR.n22 VPWR.n20 0.119
R51 VPWR.n24 VPWR.n22 0.119
R52 VPWR.n26 VPWR.n24 0.119
R53 VPWR.n28 VPWR.n26 0.119
R54 VPWR.n30 VPWR.n28 0.119
R55 VPWR VPWR.n30 0.022
R56 VPB VPB.t0 1547.82
R57 VNB VNB.t0 -7851.29
C0 VGND VPWR 2.47fF
C1 VPB VPWR 0.20fF
C2 VPB VGND 0.18fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__dfbbn_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__dfbbn_1 RESET_B VGND CLK_N SET_B Q VPWR D Q_N VNB VPB
X0 a_791_47.t0 SET_B.t0 VGND.t1 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1 a_1555_47.t0 SET_B.t1 VGND.t0 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 VPWR.t7 RESET_B.t0 a_941_21.t1 VPB.t11 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X3 a_1415_315.t0 SET_B.t2 VPWR.t1 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 a_791_47.t1 a_941_21.t2 a_647_21.t3 VNB.t9 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X5 VGND.t7 a_1415_315.t4 a_1363_47.t0 VNB.t13 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 a_1340_413.t1 a_27_47.t2 a_1256_413.t0 VPB.t18 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7 VPWR.t6 CLK_N.t0 a_27_47.t0 VPB.t8 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X8 a_381_47.t1 D.t0 VPWR.t13 VPB.t19 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9 a_473_413.t3 a_193_47.t2 a_381_47.t3 VNB.t8 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X10 a_1555_47.t2 a_941_21.t3 a_1415_315.t3 VNB.t10 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X11 VPWR.t10 a_1415_315.t5 a_2136_47.t0 VPB.t14 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X12 a_1256_413.t2 a_193_47.t3 a_1112_329.t1 VPB.t9 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13 a_581_47.t1 a_27_47.t3 a_473_413.t1 VNB.t17 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X14 a_647_21.t1 a_473_413.t4 a_791_47.t2 VNB.t11 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X15 a_647_21.t0 SET_B.t3 VPWR.t2 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16 VPWR.t9 a_941_21.t4 a_891_329.t0 VPB.t13 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X17 a_557_413.t1 a_193_47.t4 a_473_413.t2 VPB.t17 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18 a_193_47.t1 a_27_47.t4 VGND.t10 VNB.t18 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19 Q.t0 a_2136_47.t2 VPWR.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X20 a_473_413.t0 a_27_47.t5 a_381_47.t0 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21 a_891_329.t1 a_473_413.t5 a_647_21.t2 VPB.t10 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X22 Q_N.t0 a_1415_315.t6 VPWR.t4 VPB.t6 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X23 VGND.t6 RESET_B.t1 a_941_21.t0 VNB.t12 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24 Q.t1 a_2136_47.t3 VGND.t2 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X25 VPWR.t11 a_647_21.t4 a_557_413.t0 VPB.t15 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X26 a_1112_329.t0 a_647_21.t5 VPWR.t12 VPB.t16 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X27 VGND.t8 a_647_21.t6 a_581_47.t0 VNB.t14 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X28 VGND.t3 a_1415_315.t7 a_2136_47.t1 VNB.t5 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X29 a_193_47.t0 a_27_47.t6 VPWR.t3 VPB.t5 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X30 VPWR.t8 a_941_21.t5 a_1672_329.t1 VPB.t12 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X31 VPWR.t5 a_1415_315.t8 a_1340_413.t0 VPB.t7 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X32 a_1363_47.t1 a_193_47.t5 a_1256_413.t3 VNB.t16 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X33 Q_N.t1 a_1415_315.t9 VGND.t4 VNB.t6 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X34 a_381_47.t2 D.t1 VGND.t11 VNB.t19 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X35 a_1159_47.t0 a_647_21.t7 VGND.t9 VNB.t15 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X36 a_1672_329.t0 a_1256_413.t4 a_1415_315.t1 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X37 VGND.t5 CLK_N.t1 a_27_47.t1 VNB.t7 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X38 a_1256_413.t1 a_27_47.t7 a_1159_47.t1 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X39 a_1415_315.t2 a_1256_413.t5 a_1555_47.t1 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
R0 SET_B.n0 SET_B.t3 396.831
R1 SET_B.n3 SET_B.t2 391.565
R2 SET_B.n3 SET_B.t1 137.943
R3 SET_B.n0 SET_B.t0 134.063
R4 SET_B SET_B.n6 13.6
R5 SET_B.n5 SET_B.n3 12.711
R6 SET_B.n1 SET_B.n0 6.985
R7 SET_B.n6 SET_B.n5 6.318
R8 SET_B.n6 SET_B.n1 2.521
R9 SET_B.n2 SET_B 2.521
R10 SET_B.n6 SET_B.n2 0.775
R11 SET_B.n5 SET_B.n4 0.001
R12 VGND.n24 VGND.t9 187.166
R13 VGND.n43 VGND.t11 144.772
R14 VGND.n34 VGND.n33 113.205
R15 VGND.n3 VGND.n0 112.777
R16 VGND.n2 VGND.n1 108.447
R17 VGND.n48 VGND.n47 107.239
R18 VGND.n13 VGND.n12 106.678
R19 VGND.n33 VGND.t8 81.428
R20 VGND.n12 VGND.t7 57.142
R21 VGND.n0 VGND.t3 54.285
R22 VGND.n1 VGND.t6 54.285
R23 VGND.n12 VGND.t0 38.571
R24 VGND.n33 VGND.t1 38.571
R25 VGND.n47 VGND.t10 38.571
R26 VGND.n47 VGND.t5 38.571
R27 VGND.n0 VGND.t2 25.934
R28 VGND.n1 VGND.t4 25.934
R29 VGND.n35 VGND.n34 16.564
R30 VGND.n5 VGND.n4 4.65
R31 VGND.n7 VGND.n6 4.65
R32 VGND.n9 VGND.n8 4.65
R33 VGND.n11 VGND.n10 4.65
R34 VGND.n15 VGND.n14 4.65
R35 VGND.n17 VGND.n16 4.65
R36 VGND.n19 VGND.n18 4.65
R37 VGND.n21 VGND.n20 4.65
R38 VGND.n23 VGND.n22 4.65
R39 VGND.n26 VGND.n25 4.65
R40 VGND.n28 VGND.n27 4.65
R41 VGND.n30 VGND.n29 4.65
R42 VGND.n32 VGND.n31 4.65
R43 VGND.n36 VGND.n35 4.65
R44 VGND.n38 VGND.n37 4.65
R45 VGND.n40 VGND.n39 4.65
R46 VGND.n42 VGND.n41 4.65
R47 VGND.n44 VGND.n43 4.65
R48 VGND.n46 VGND.n45 4.65
R49 VGND.n3 VGND.n2 3.969
R50 VGND.n49 VGND.n48 3.932
R51 VGND.n25 VGND.n24 2.635
R52 VGND.n14 VGND.n13 1.129
R53 VGND.n5 VGND.n3 0.146
R54 VGND.n49 VGND.n46 0.137
R55 VGND VGND.n49 0.123
R56 VGND.n7 VGND.n5 0.119
R57 VGND.n9 VGND.n7 0.119
R58 VGND.n11 VGND.n9 0.119
R59 VGND.n15 VGND.n11 0.119
R60 VGND.n17 VGND.n15 0.119
R61 VGND.n19 VGND.n17 0.119
R62 VGND.n21 VGND.n19 0.119
R63 VGND.n23 VGND.n21 0.119
R64 VGND.n26 VGND.n23 0.119
R65 VGND.n28 VGND.n26 0.119
R66 VGND.n30 VGND.n28 0.119
R67 VGND.n32 VGND.n30 0.119
R68 VGND.n36 VGND.n32 0.119
R69 VGND.n38 VGND.n36 0.119
R70 VGND.n40 VGND.n38 0.119
R71 VGND.n42 VGND.n40 0.119
R72 VGND.n44 VGND.n42 0.119
R73 VGND.n46 VGND.n44 0.119
R74 a_791_47.t1 a_791_47.n0 283.512
R75 a_791_47.n0 a_791_47.t2 42.946
R76 a_791_47.n0 a_791_47.t0 38.571
R77 VNB.t18 VNB.t19 6082.35
R78 VNB.t10 VNB.t12 4595.56
R79 VNB.t9 VNB.t15 4595.56
R80 VNB.t6 VNB.t5 4545.05
R81 VNB VNB.t7 4270.59
R82 VNB.t14 VNB.t1 3688.24
R83 VNB.t8 VNB.t17 3397.06
R84 VNB.t15 VNB.t4 3162.68
R85 VNB.t13 VNB.t0 3138.24
R86 VNB.t17 VNB.t14 3105.88
R87 VNB.t16 VNB.t13 3073.53
R88 VNB.t19 VNB.t8 3073.53
R89 VNB.t0 VNB.t2 2774.44
R90 VNB.t4 VNB.t16 2717.65
R91 VNB.t7 VNB.t18 2717.65
R92 VNB.t1 VNB.t11 2304.58
R93 VNB.t5 VNB.t3 2296.7
R94 VNB.t12 VNB.t6 2248.62
R95 VNB.t2 VNB.t10 2053.33
R96 VNB.t11 VNB.t9 2053.33
R97 a_1555_47.n0 a_1555_47.t2 277.452
R98 a_1555_47.t1 a_1555_47.n0 60.579
R99 a_1555_47.n0 a_1555_47.t0 38.571
R100 RESET_B.n0 RESET_B.t1 202.557
R101 RESET_B.n0 RESET_B.t0 173.636
R102 RESET_B RESET_B.n0 78.109
R103 a_941_21.t1 a_941_21.n3 445.092
R104 a_941_21.n1 a_941_21.t3 211.734
R105 a_941_21.n0 a_941_21.t2 210.472
R106 a_941_21.n1 a_941_21.t5 205.308
R107 a_941_21.n0 a_941_21.t4 204.046
R108 a_941_21.n2 a_941_21.t0 197.012
R109 a_941_21.n3 a_941_21.n0 126.517
R110 a_941_21.n2 a_941_21.n1 76
R111 a_941_21.n3 a_941_21.n2 9.431
R112 VPWR.n6 VPWR.t8 500.865
R113 VPWR.n1 VPWR.n0 440.25
R114 VPWR.n44 VPWR.t13 373.849
R115 VPWR.n49 VPWR.n48 311.893
R116 VPWR.n36 VPWR.n35 306.984
R117 VPWR.n14 VPWR.n13 292.5
R118 VPWR.n3 VPWR.n2 173.128
R119 VPWR.n28 VPWR.n27 164.214
R120 VPWR.n13 VPWR.t5 121.952
R121 VPWR.n13 VPWR.t1 91.464
R122 VPWR.n35 VPWR.t2 91.464
R123 VPWR.n27 VPWR.t12 86.773
R124 VPWR.n35 VPWR.t11 86.773
R125 VPWR.n0 VPWR.t7 63.101
R126 VPWR.n2 VPWR.t10 58.484
R127 VPWR.n48 VPWR.t3 41.554
R128 VPWR.n48 VPWR.t6 41.554
R129 VPWR.n27 VPWR.t9 38.696
R130 VPWR.n2 VPWR.t0 31.83
R131 VPWR.n0 VPWR.t4 28.032
R132 VPWR.n5 VPWR.n4 4.65
R133 VPWR.n8 VPWR.n7 4.65
R134 VPWR.n10 VPWR.n9 4.65
R135 VPWR.n12 VPWR.n11 4.65
R136 VPWR.n16 VPWR.n15 4.65
R137 VPWR.n18 VPWR.n17 4.65
R138 VPWR.n20 VPWR.n19 4.65
R139 VPWR.n22 VPWR.n21 4.65
R140 VPWR.n24 VPWR.n23 4.65
R141 VPWR.n26 VPWR.n25 4.65
R142 VPWR.n30 VPWR.n29 4.65
R143 VPWR.n32 VPWR.n31 4.65
R144 VPWR.n34 VPWR.n33 4.65
R145 VPWR.n37 VPWR.n36 4.65
R146 VPWR.n39 VPWR.n38 4.65
R147 VPWR.n41 VPWR.n40 4.65
R148 VPWR.n43 VPWR.n42 4.65
R149 VPWR.n45 VPWR.n44 4.65
R150 VPWR.n47 VPWR.n46 4.65
R151 VPWR.n3 VPWR.n1 4.611
R152 VPWR.n50 VPWR.n49 3.932
R153 VPWR.n29 VPWR.n28 3.388
R154 VPWR.n7 VPWR.n6 2.676
R155 VPWR.n15 VPWR.n14 2.443
R156 VPWR.n5 VPWR.n3 0.144
R157 VPWR.n50 VPWR.n47 0.137
R158 VPWR VPWR.n50 0.123
R159 VPWR.n8 VPWR.n5 0.119
R160 VPWR.n10 VPWR.n8 0.119
R161 VPWR.n12 VPWR.n10 0.119
R162 VPWR.n16 VPWR.n12 0.119
R163 VPWR.n18 VPWR.n16 0.119
R164 VPWR.n20 VPWR.n18 0.119
R165 VPWR.n22 VPWR.n20 0.119
R166 VPWR.n24 VPWR.n22 0.119
R167 VPWR.n26 VPWR.n24 0.119
R168 VPWR.n30 VPWR.n26 0.119
R169 VPWR.n32 VPWR.n30 0.119
R170 VPWR.n34 VPWR.n32 0.119
R171 VPWR.n37 VPWR.n34 0.119
R172 VPWR.n39 VPWR.n37 0.119
R173 VPWR.n41 VPWR.n39 0.119
R174 VPWR.n43 VPWR.n41 0.119
R175 VPWR.n45 VPWR.n43 0.119
R176 VPWR.n47 VPWR.n45 0.119
R177 VPB.t12 VPB.t11 559.345
R178 VPB.t6 VPB.t14 556.386
R179 VPB.t5 VPB.t19 556.386
R180 VPB.t16 VPB.t9 426.168
R181 VPB.t13 VPB.t16 405.451
R182 VPB.t7 VPB.t2 358.099
R183 VPB.t17 VPB.t15 355.14
R184 VPB.t1 VPB.t10 319.626
R185 VPB.t2 VPB.t3 313.707
R186 VPB.t15 VPB.t1 313.707
R187 VPB.t18 VPB.t7 310.747
R188 VPB.t11 VPB.t6 287.071
R189 VPB.t14 VPB.t0 281.152
R190 VPB.t19 VPB.t4 272.274
R191 VPB.t9 VPB.t18 248.598
R192 VPB.t10 VPB.t13 248.598
R193 VPB.t4 VPB.t17 248.598
R194 VPB.t8 VPB.t5 248.598
R195 VPB.t3 VPB.t12 213.084
R196 VPB VPB.t8 142.056
R197 a_1415_315.n4 a_1415_315.t4 383.24
R198 a_1415_315.n6 a_1415_315.n5 301.911
R199 a_1415_315.n2 a_1415_315.t6 268.312
R200 a_1415_315.n3 a_1415_315.n2 236.062
R201 a_1415_315.n1 a_1415_315.t5 231.942
R202 a_1415_315.n2 a_1415_315.t9 222.789
R203 a_1415_315.n3 a_1415_315.n0 179.668
R204 a_1415_315.n1 a_1415_315.t7 164.463
R205 a_1415_315.n2 a_1415_315.n1 151.74
R206 a_1415_315.n4 a_1415_315.t8 139.027
R207 a_1415_315.n5 a_1415_315.n4 128.841
R208 a_1415_315.n6 a_1415_315.t0 91.464
R209 a_1415_315.t1 a_1415_315.n6 57.457
R210 a_1415_315.n5 a_1415_315.n3 36.894
R211 a_1415_315.n0 a_1415_315.t3 25.312
R212 a_1415_315.n0 a_1415_315.t2 25.312
R213 a_647_21.n5 a_647_21.t6 387.959
R214 a_647_21.n2 a_647_21.t5 299.91
R215 a_647_21.n7 a_647_21.n6 292.5
R216 a_647_21.n2 a_647_21.t7 167.627
R217 a_647_21.n5 a_647_21.t4 143.746
R218 a_647_21.n4 a_647_21.n2 139.816
R219 a_647_21.n6 a_647_21.n5 114.656
R220 a_647_21.n0 a_647_21.t0 110.226
R221 a_647_21.n4 a_647_21.n3 109.954
R222 a_647_21.n6 a_647_21.n4 81.172
R223 a_647_21.t2 a_647_21.n1 63.321
R224 a_647_21.t2 a_647_21.n7 63.321
R225 a_647_21.n3 a_647_21.t3 25.312
R226 a_647_21.n3 a_647_21.t1 25.312
R227 a_647_21.n1 a_647_21.n0 9.38
R228 a_1363_47.t0 a_1363_47.t1 93.059
R229 a_27_47.n2 a_27_47.t5 538.597
R230 a_27_47.t0 a_27_47.n5 279.118
R231 a_27_47.n1 a_27_47.t2 272.021
R232 a_27_47.n0 a_27_47.t6 262.942
R233 a_27_47.n0 a_27_47.t4 227.596
R234 a_27_47.n1 a_27_47.t7 209.695
R235 a_27_47.n4 a_27_47.t1 174.068
R236 a_27_47.n2 a_27_47.t3 135.786
R237 a_27_47.n5 a_27_47.n0 76
R238 a_27_47.n5 a_27_47.n4 21.426
R239 a_27_47.n3 a_27_47.n1 11.94
R240 a_27_47.n3 a_27_47.n2 10.203
R241 a_27_47.n4 a_27_47.n3 6.591
R242 a_1256_413.n3 a_1256_413.n2 399.793
R243 a_1256_413.n1 a_1256_413.t4 236.933
R244 a_1256_413.n1 a_1256_413.t5 191.945
R245 a_1256_413.n2 a_1256_413.n0 180.236
R246 a_1256_413.n2 a_1256_413.n1 159.918
R247 a_1256_413.t0 a_1256_413.n3 63.321
R248 a_1256_413.n3 a_1256_413.t2 63.321
R249 a_1256_413.n0 a_1256_413.t3 45
R250 a_1256_413.n0 a_1256_413.t1 45
R251 a_1340_413.t0 a_1340_413.t1 175.892
R252 CLK_N.n0 CLK_N.t0 272.06
R253 CLK_N.n0 CLK_N.t1 236.714
R254 CLK_N.n1 CLK_N.n0 76
R255 CLK_N CLK_N.n1 7.68
R256 CLK_N.n1 CLK_N 4.754
R257 D.n0 D.t0 331.508
R258 D.n0 D.t1 209.401
R259 D.n1 D.n0 76
R260 D.n1 D 8.585
R261 D D.n1 2.029
R262 a_381_47.n1 a_381_47.n0 574.144
R263 a_381_47.t0 a_381_47.n1 82.083
R264 a_381_47.n0 a_381_47.t3 63.333
R265 a_381_47.n1 a_381_47.t1 63.321
R266 a_381_47.n0 a_381_47.t2 29.726
R267 a_193_47.n0 a_193_47.t5 534.467
R268 a_193_47.n1 a_193_47.t2 238.651
R269 a_193_47.n1 a_193_47.t4 231.324
R270 a_193_47.n3 a_193_47.t1 210.124
R271 a_193_47.n0 a_193_47.t3 137.933
R272 a_193_47.t0 a_193_47.n3 121.825
R273 a_193_47.n2 a_193_47.n0 12.947
R274 a_193_47.n2 a_193_47.n1 4.65
R275 a_193_47.n3 a_193_47.n2 2.663
R276 a_473_413.n3 a_473_413.n2 415.031
R277 a_473_413.n1 a_473_413.t4 216.899
R278 a_473_413.n1 a_473_413.t5 210.473
R279 a_473_413.n2 a_473_413.n0 196.424
R280 a_473_413.n2 a_473_413.n1 140.828
R281 a_473_413.n0 a_473_413.t1 63.333
R282 a_473_413.n3 a_473_413.t2 63.321
R283 a_473_413.t0 a_473_413.n3 63.321
R284 a_473_413.n0 a_473_413.t3 61.666
R285 a_2136_47.n0 a_2136_47.t2 239.038
R286 a_2136_47.t0 a_2136_47.n1 237.868
R287 a_2136_47.n0 a_2136_47.t3 166.738
R288 a_2136_47.n1 a_2136_47.t1 150.778
R289 a_2136_47.n1 a_2136_47.n0 99.078
R290 a_1112_329.t0 a_1112_329.t1 236.868
R291 a_581_47.t0 a_581_47.t1 93.516
R292 a_891_329.t0 a_891_329.t1 63.321
R293 a_557_413.t0 a_557_413.t1 211.071
R294 Q.n1 Q.t0 207.372
R295 Q.n0 Q.t1 117.423
R296 Q Q.n0 67.692
R297 Q.n1 Q 9.019
R298 Q Q.n1 7.458
R299 Q.n0 Q 6.646
R300 Q_N.n1 Q_N.t0 207.566
R301 Q_N.n0 Q_N.t1 117.423
R302 Q_N Q_N.n0 79.437
R303 Q_N.n1 Q_N 8.185
R304 Q_N Q_N.n1 6.859
R305 Q_N.n0 Q_N 5.614
R306 a_1672_329.t0 a_1672_329.t1 49.25
R307 a_1159_47.n0 a_1159_47.t1 108.333
R308 a_1159_47.n1 a_1159_47.n0 67.2
R309 a_1159_47.n0 a_1159_47.t0 13.143
C0 SET_B VGND 0.39fF
C1 VPB VPWR 0.25fF
C2 VGND Q_N 0.12fF
C3 VPWR Q 0.14fF
C4 VPWR VGND 0.12fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__dfbbn_2.ext - technology: sky130A

.subckt sky130_fd_sc_hd__dfbbn_2 RESET_B VGND CLK_N SET_B Q VPWR D Q_N VNB VPB
X0 a_790_47.t0 SET_B.t0 VGND.t12 VNB.t17 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1 a_790_47.t1 a_944_21.t2 a_650_21.t0 VNB.t18 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X2 Q_N.t3 a_1431_21.t4 VPWR.t3 VPB.t5 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 a_894_329.t1 a_476_47.t4 a_650_21.t2 VPB.t20 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X4 a_476_47.t0 a_27_47.t2 a_381_47.t3 VPB.t13 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 VGND.t6 a_650_21.t4 a_584_47.t0 VNB.t11 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 VPWR.t9 a_2236_47.t2 Q.t3 VPB.t10 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 VPWR.t8 a_650_21.t5 a_560_413.t0 VPB.t8 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 a_1547_47.t0 a_944_21.t3 a_1431_21.t0 VNB.t19 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X9 VPWR.t11 CLK_N.t0 a_27_47.t0 VPB.t12 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X10 Q.t2 a_2236_47.t3 VPWR.t10 VPB.t11 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 a_381_47.t0 D.t0 VPWR.t6 VPB.t6 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12 a_1115_329.t0 a_650_21.t6 VPWR.t7 VPB.t7 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X13 a_476_47.t2 a_193_47.t2 a_381_47.t2 VNB.t9 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X14 a_584_47.t1 a_27_47.t3 a_476_47.t1 VNB.t6 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X15 VPWR.t0 a_944_21.t4 a_894_329.t0 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X16 a_1162_47.t0 a_650_21.t7 VGND.t4 VNB.t5 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X17 VGND.t7 a_1431_21.t5 Q_N.t1 VNB.t12 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X18 Q.t1 a_2236_47.t4 VGND.t1 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X19 VGND.t8 a_1431_21.t6 a_2236_47.t0 VNB.t13 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20 a_193_47.t0 a_27_47.t4 VGND.t5 VNB.t7 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21 VPWR.t15 RESET_B.t0 a_944_21.t0 VPB.t21 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X22 Q_N.t0 a_1431_21.t7 VGND.t9 VNB.t14 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X23 VPWR.t4 a_1431_21.t8 a_1343_413.t0 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24 VPWR.t1 a_944_21.t5 a_1665_329.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X25 VGND.t10 a_1431_21.t9 a_1366_47.t1 VNB.t15 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X26 VGND.t2 a_2236_47.t5 Q.t0 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X27 a_1431_21.t3 SET_B.t1 VPWR.t13 VPB.t19 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X28 VPWR.t5 a_1431_21.t10 Q_N.t2 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X29 a_1366_47.t0 a_193_47.t3 a_1257_47.t1 VNB.t10 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X30 a_1665_329.t1 a_1257_47.t4 a_1431_21.t1 VPB.t9 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X31 a_1257_47.t3 a_27_47.t5 a_1162_47.t1 VNB.t8 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X32 a_193_47.t1 a_27_47.t6 VPWR.t12 VPB.t14 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X33 a_1343_413.t1 a_27_47.t7 a_1257_47.t2 VPB.t15 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X34 a_1547_47.t2 SET_B.t2 VGND.t11 VNB.t16 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X35 a_650_21.t3 a_476_47.t5 a_790_47.t2 VNB.t20 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X36 a_1257_47.t0 a_193_47.t4 a_1115_329.t1 VPB.t16 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X37 a_381_47.t1 D.t1 VGND.t0 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X38 a_1431_21.t2 a_1257_47.t5 a_1547_47.t1 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X39 a_650_21.t1 SET_B.t3 VPWR.t14 VPB.t18 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X40 VPWR.t2 a_1431_21.t11 a_2236_47.t1 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X41 VGND.t13 RESET_B.t1 a_944_21.t1 VNB.t21 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X42 a_560_413.t1 a_193_47.t5 a_476_47.t3 VPB.t17 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X43 VGND.t3 CLK_N.t1 a_27_47.t1 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
R0 SET_B.n0 SET_B.t3 397.142
R1 SET_B.n3 SET_B.t1 394.428
R2 SET_B.n0 SET_B.t0 134.984
R3 SET_B.n3 SET_B.t2 134.495
R4 SET_B SET_B.n6 13.6
R5 SET_B.n5 SET_B.n3 13.011
R6 SET_B.n1 SET_B.n0 6.954
R7 SET_B.n6 SET_B.n5 6.318
R8 SET_B.n6 SET_B.n1 2.521
R9 SET_B.n2 SET_B 2.521
R10 SET_B.n6 SET_B.n2 0.775
R11 SET_B.n5 SET_B.n4 0.001
R12 VGND.n30 VGND.t4 188.008
R13 VGND.n51 VGND.t0 145.376
R14 VGND.n42 VGND.n41 113.205
R15 VGND.n2 VGND.t2 110.775
R16 VGND.n21 VGND.n20 110.223
R17 VGND.n1 VGND.n0 108.988
R18 VGND.n56 VGND.n55 107.239
R19 VGND.n5 VGND.t7 103.996
R20 VGND.n41 VGND.t6 75.714
R21 VGND.n10 VGND.n9 64.275
R22 VGND.n9 VGND.t13 57.796
R23 VGND.n0 VGND.t8 54.285
R24 VGND.n20 VGND.t10 41.428
R25 VGND.n20 VGND.t11 38.571
R26 VGND.n41 VGND.t12 38.571
R27 VGND.n55 VGND.t5 38.571
R28 VGND.n55 VGND.t3 38.571
R29 VGND.n0 VGND.t1 25.934
R30 VGND.n9 VGND.t9 24.765
R31 VGND.n43 VGND.n42 16.188
R32 VGND.n4 VGND.n3 4.65
R33 VGND.n6 VGND.n5 4.65
R34 VGND.n8 VGND.n7 4.65
R35 VGND.n11 VGND.n10 4.65
R36 VGND.n13 VGND.n12 4.65
R37 VGND.n15 VGND.n14 4.65
R38 VGND.n17 VGND.n16 4.65
R39 VGND.n19 VGND.n18 4.65
R40 VGND.n23 VGND.n22 4.65
R41 VGND.n25 VGND.n24 4.65
R42 VGND.n27 VGND.n26 4.65
R43 VGND.n29 VGND.n28 4.65
R44 VGND.n32 VGND.n31 4.65
R45 VGND.n34 VGND.n33 4.65
R46 VGND.n36 VGND.n35 4.65
R47 VGND.n38 VGND.n37 4.65
R48 VGND.n40 VGND.n39 4.65
R49 VGND.n44 VGND.n43 4.65
R50 VGND.n46 VGND.n45 4.65
R51 VGND.n48 VGND.n47 4.65
R52 VGND.n50 VGND.n49 4.65
R53 VGND.n52 VGND.n51 4.65
R54 VGND.n54 VGND.n53 4.65
R55 VGND.n31 VGND.n30 4.517
R56 VGND.n22 VGND.n21 4.141
R57 VGND.n57 VGND.n56 3.932
R58 VGND.n2 VGND.n1 3.724
R59 VGND.n4 VGND.n2 0.252
R60 VGND.n57 VGND.n54 0.137
R61 VGND VGND.n57 0.121
R62 VGND.n6 VGND.n4 0.119
R63 VGND.n8 VGND.n6 0.119
R64 VGND.n11 VGND.n8 0.119
R65 VGND.n13 VGND.n11 0.119
R66 VGND.n15 VGND.n13 0.119
R67 VGND.n17 VGND.n15 0.119
R68 VGND.n19 VGND.n17 0.119
R69 VGND.n23 VGND.n19 0.119
R70 VGND.n25 VGND.n23 0.119
R71 VGND.n27 VGND.n25 0.119
R72 VGND.n29 VGND.n27 0.119
R73 VGND.n32 VGND.n29 0.119
R74 VGND.n34 VGND.n32 0.119
R75 VGND.n36 VGND.n34 0.119
R76 VGND.n38 VGND.n36 0.119
R77 VGND.n40 VGND.n38 0.119
R78 VGND.n44 VGND.n40 0.119
R79 VGND.n46 VGND.n44 0.119
R80 VGND.n48 VGND.n46 0.119
R81 VGND.n50 VGND.n48 0.119
R82 VGND.n52 VGND.n50 0.119
R83 VGND.n54 VGND.n52 0.119
R84 a_790_47.t1 a_790_47.n0 278.793
R85 a_790_47.n0 a_790_47.t2 49.151
R86 a_790_47.n0 a_790_47.t0 38.571
R87 VNB.t7 VNB.t0 6082.35
R88 VNB.t12 VNB.t13 4738.46
R89 VNB.t19 VNB.t21 4693.33
R90 VNB.t18 VNB.t5 4595.56
R91 VNB VNB.t4 4238.23
R92 VNB.t11 VNB.t17 3558.82
R93 VNB.t8 VNB.t10 3526.47
R94 VNB.t9 VNB.t6 3494.12
R95 VNB.t6 VNB.t11 3105.88
R96 VNB.t16 VNB.t1 3097.97
R97 VNB.t10 VNB.t15 3073.53
R98 VNB.t0 VNB.t9 3073.53
R99 VNB.t15 VNB.t16 2782.35
R100 VNB.t4 VNB.t7 2717.65
R101 VNB.t17 VNB.t20 2349.76
R102 VNB.t21 VNB.t14 2296.97
R103 VNB.t13 VNB.t2 2296.7
R104 VNB.t5 VNB.t8 2280.14
R105 VNB.t1 VNB.t19 2053.33
R106 VNB.t20 VNB.t18 2053.33
R107 VNB.t2 VNB.t3 2030.77
R108 VNB.t14 VNB.t12 2030.77
R109 a_944_21.t0 a_944_21.n3 441.973
R110 a_944_21.n1 a_944_21.t3 211.734
R111 a_944_21.n0 a_944_21.t2 210.472
R112 a_944_21.n1 a_944_21.t5 207.402
R113 a_944_21.n0 a_944_21.t4 204.046
R114 a_944_21.n2 a_944_21.t1 194.506
R115 a_944_21.n3 a_944_21.n0 126.544
R116 a_944_21.n2 a_944_21.n1 76
R117 a_944_21.n3 a_944_21.n2 9.774
R118 a_650_21.n5 a_650_21.t4 387.959
R119 a_650_21.n2 a_650_21.t6 299.91
R120 a_650_21.n7 a_650_21.n6 292.5
R121 a_650_21.n2 a_650_21.t7 167.627
R122 a_650_21.n5 a_650_21.t5 143.746
R123 a_650_21.n4 a_650_21.n2 139.816
R124 a_650_21.n6 a_650_21.n5 114.656
R125 a_650_21.n0 a_650_21.t1 110.226
R126 a_650_21.n4 a_650_21.n3 109.954
R127 a_650_21.n6 a_650_21.n4 81.172
R128 a_650_21.t2 a_650_21.n1 63.321
R129 a_650_21.t2 a_650_21.n7 63.321
R130 a_650_21.n3 a_650_21.t0 25.312
R131 a_650_21.n3 a_650_21.t3 25.312
R132 a_650_21.n1 a_650_21.n0 9.38
R133 a_1431_21.n5 a_1431_21.t9 387.206
R134 a_1431_21.n2 a_1431_21.t4 308.479
R135 a_1431_21.n7 a_1431_21.n6 301.911
R136 a_1431_21.n2 a_1431_21.t7 236.179
R137 a_1431_21.n4 a_1431_21.n2 231.623
R138 a_1431_21.n0 a_1431_21.t11 231.473
R139 a_1431_21.n1 a_1431_21.t10 221.719
R140 a_1431_21.n4 a_1431_21.n3 183.133
R141 a_1431_21.n0 a_1431_21.t6 163.994
R142 a_1431_21.n1 a_1431_21.n0 151.74
R143 a_1431_21.n1 a_1431_21.t5 149.419
R144 a_1431_21.n5 a_1431_21.t8 142.993
R145 a_1431_21.n6 a_1431_21.n5 128.841
R146 a_1431_21.n7 a_1431_21.t3 91.464
R147 a_1431_21.n2 a_1431_21.n1 85.688
R148 a_1431_21.t1 a_1431_21.n7 32.833
R149 a_1431_21.n6 a_1431_21.n4 30.494
R150 a_1431_21.n3 a_1431_21.t0 25.312
R151 a_1431_21.n3 a_1431_21.t2 25.312
R152 VPWR.n15 VPWR.t1 500.865
R153 VPWR.n10 VPWR.n9 440.25
R154 VPWR.n53 VPWR.t6 374.644
R155 VPWR.n58 VPWR.n57 311.893
R156 VPWR.n45 VPWR.n44 306.984
R157 VPWR.n23 VPWR.n22 292.5
R158 VPWR.n1 VPWR.n0 168.939
R159 VPWR.n5 VPWR.t5 164.708
R160 VPWR.n37 VPWR.n36 164.214
R161 VPWR.n2 VPWR.t9 155.131
R162 VPWR.n22 VPWR.t13 91.464
R163 VPWR.n22 VPWR.t4 91.464
R164 VPWR.n44 VPWR.t14 91.464
R165 VPWR.n36 VPWR.t7 86.773
R166 VPWR.n44 VPWR.t8 86.773
R167 VPWR.n9 VPWR.t15 63.101
R168 VPWR.n0 VPWR.t2 58.484
R169 VPWR.n36 VPWR.t0 43.386
R170 VPWR.n57 VPWR.t12 41.554
R171 VPWR.n57 VPWR.t11 41.554
R172 VPWR.n0 VPWR.t10 31.83
R173 VPWR.n9 VPWR.t3 27.786
R174 VPWR.n4 VPWR.n3 4.65
R175 VPWR.n6 VPWR.n5 4.65
R176 VPWR.n8 VPWR.n7 4.65
R177 VPWR.n12 VPWR.n11 4.65
R178 VPWR.n14 VPWR.n13 4.65
R179 VPWR.n17 VPWR.n16 4.65
R180 VPWR.n19 VPWR.n18 4.65
R181 VPWR.n21 VPWR.n20 4.65
R182 VPWR.n25 VPWR.n24 4.65
R183 VPWR.n27 VPWR.n26 4.65
R184 VPWR.n29 VPWR.n28 4.65
R185 VPWR.n31 VPWR.n30 4.65
R186 VPWR.n33 VPWR.n32 4.65
R187 VPWR.n35 VPWR.n34 4.65
R188 VPWR.n39 VPWR.n38 4.65
R189 VPWR.n41 VPWR.n40 4.65
R190 VPWR.n43 VPWR.n42 4.65
R191 VPWR.n46 VPWR.n45 4.65
R192 VPWR.n48 VPWR.n47 4.65
R193 VPWR.n50 VPWR.n49 4.65
R194 VPWR.n52 VPWR.n51 4.65
R195 VPWR.n54 VPWR.n53 4.65
R196 VPWR.n56 VPWR.n55 4.65
R197 VPWR.n38 VPWR.n37 4.517
R198 VPWR.n59 VPWR.n58 3.932
R199 VPWR.n2 VPWR.n1 3.724
R200 VPWR.n16 VPWR.n15 3.49
R201 VPWR.n24 VPWR.n23 2.094
R202 VPWR.n11 VPWR.n10 0.349
R203 VPWR.n4 VPWR.n2 0.252
R204 VPWR.n59 VPWR.n56 0.137
R205 VPWR VPWR.n59 0.121
R206 VPWR.n6 VPWR.n4 0.119
R207 VPWR.n8 VPWR.n6 0.119
R208 VPWR.n12 VPWR.n8 0.119
R209 VPWR.n14 VPWR.n12 0.119
R210 VPWR.n17 VPWR.n14 0.119
R211 VPWR.n19 VPWR.n17 0.119
R212 VPWR.n21 VPWR.n19 0.119
R213 VPWR.n25 VPWR.n21 0.119
R214 VPWR.n27 VPWR.n25 0.119
R215 VPWR.n29 VPWR.n27 0.119
R216 VPWR.n31 VPWR.n29 0.119
R217 VPWR.n33 VPWR.n31 0.119
R218 VPWR.n35 VPWR.n33 0.119
R219 VPWR.n39 VPWR.n35 0.119
R220 VPWR.n41 VPWR.n39 0.119
R221 VPWR.n43 VPWR.n41 0.119
R222 VPWR.n46 VPWR.n43 0.119
R223 VPWR.n48 VPWR.n46 0.119
R224 VPWR.n50 VPWR.n48 0.119
R225 VPWR.n52 VPWR.n50 0.119
R226 VPWR.n54 VPWR.n52 0.119
R227 VPWR.n56 VPWR.n54 0.119
R228 Q_N.n3 Q_N.n2 142.9
R229 Q_N.n1 Q_N.n0 92.5
R230 Q_N Q_N.n1 80.819
R231 Q_N.n2 Q_N.t2 26.595
R232 Q_N.n2 Q_N.t3 26.595
R233 Q_N.n0 Q_N.t1 24.923
R234 Q_N.n0 Q_N.t0 24.923
R235 Q_N.n3 Q_N 8.895
R236 Q_N Q_N.n3 7.456
R237 Q_N.n1 Q_N 6.153
R238 VPB.t0 VPB.t21 603.738
R239 VPB.t3 VPB.t2 580.062
R240 VPB.t14 VPB.t6 556.386
R241 VPB.t7 VPB.t16 426.168
R242 VPB.t1 VPB.t7 417.289
R243 VPB.t17 VPB.t8 355.14
R244 VPB.t15 VPB.t4 349.221
R245 VPB.t4 VPB.t19 319.626
R246 VPB.t18 VPB.t20 319.626
R247 VPB.t8 VPB.t18 313.707
R248 VPB.t21 VPB.t5 287.071
R249 VPB.t19 VPB.t9 284.112
R250 VPB.t2 VPB.t11 281.152
R251 VPB.t6 VPB.t13 281.152
R252 VPB.t11 VPB.t10 248.598
R253 VPB.t5 VPB.t3 248.598
R254 VPB.t16 VPB.t15 248.598
R255 VPB.t13 VPB.t17 248.598
R256 VPB.t12 VPB.t14 248.598
R257 VPB.t20 VPB.t1 236.76
R258 VPB.t9 VPB.t0 213.084
R259 VPB VPB.t12 139.096
R260 a_476_47.n3 a_476_47.n2 413.812
R261 a_476_47.n1 a_476_47.t5 216.899
R262 a_476_47.n1 a_476_47.t4 210.473
R263 a_476_47.n2 a_476_47.n0 195.144
R264 a_476_47.n2 a_476_47.n1 142.333
R265 a_476_47.n0 a_476_47.t2 66.666
R266 a_476_47.n0 a_476_47.t1 63.333
R267 a_476_47.n3 a_476_47.t3 63.321
R268 a_476_47.t0 a_476_47.n3 63.321
R269 a_894_329.t0 a_894_329.t1 58.63
R270 a_27_47.n2 a_27_47.t2 538.588
R271 a_27_47.t0 a_27_47.n5 274.6
R272 a_27_47.n1 a_27_47.t7 267.397
R273 a_27_47.n0 a_27_47.t6 263.171
R274 a_27_47.n0 a_27_47.t4 227.825
R275 a_27_47.n1 a_27_47.t5 207.297
R276 a_27_47.n4 a_27_47.t1 168.595
R277 a_27_47.n2 a_27_47.t3 135.791
R278 a_27_47.n5 a_27_47.n0 76
R279 a_27_47.n5 a_27_47.n4 21.426
R280 a_27_47.n3 a_27_47.n2 10.055
R281 a_27_47.n3 a_27_47.n1 7.532
R282 a_27_47.n4 a_27_47.n3 6.59
R283 a_381_47.n1 a_381_47.n0 572.005
R284 a_381_47.n1 a_381_47.t3 89.119
R285 a_381_47.n0 a_381_47.t2 63.333
R286 a_381_47.t0 a_381_47.n1 63.321
R287 a_381_47.n0 a_381_47.t1 29.726
R288 a_584_47.t0 a_584_47.t1 93.516
R289 a_2236_47.t1 a_2236_47.n2 244.259
R290 a_2236_47.n0 a_2236_47.t2 212.079
R291 a_2236_47.n1 a_2236_47.t3 212.079
R292 a_2236_47.n2 a_2236_47.t0 155.416
R293 a_2236_47.n0 a_2236_47.t5 139.779
R294 a_2236_47.n1 a_2236_47.t4 139.779
R295 a_2236_47.n2 a_2236_47.n1 110.33
R296 a_2236_47.n1 a_2236_47.n0 61.345
R297 Q.n3 Q.n2 142.612
R298 Q.n1 Q.n0 92.5
R299 Q Q.n1 76.565
R300 Q.n2 Q.t3 26.595
R301 Q.n2 Q.t2 26.595
R302 Q.n0 Q.t0 24.923
R303 Q.n0 Q.t1 24.923
R304 Q.n3 Q 10.168
R305 Q Q.n3 8.276
R306 Q.n1 Q 7.513
R307 a_560_413.t0 a_560_413.t1 211.071
R308 a_1547_47.t0 a_1547_47.n0 274.441
R309 a_1547_47.n0 a_1547_47.t2 64.285
R310 a_1547_47.n0 a_1547_47.t1 49.151
R311 CLK_N.n0 CLK_N.t0 269.919
R312 CLK_N.n0 CLK_N.t1 234.573
R313 CLK_N.n1 CLK_N.n0 76
R314 CLK_N CLK_N.n1 7.571
R315 CLK_N.n1 CLK_N 4.687
R316 D.n0 D.t0 331.508
R317 D.n0 D.t1 209.401
R318 D.n1 D.n0 76
R319 D.n1 D 8.585
R320 D D.n1 2.029
R321 a_1115_329.t0 a_1115_329.t1 236.868
R322 a_193_47.n0 a_193_47.t3 534.467
R323 a_193_47.n1 a_193_47.t2 237.504
R324 a_193_47.n1 a_193_47.t5 231.324
R325 a_193_47.n3 a_193_47.t0 208.379
R326 a_193_47.n0 a_193_47.t4 137.933
R327 a_193_47.t1 a_193_47.n3 121.759
R328 a_193_47.n2 a_193_47.n0 12.947
R329 a_193_47.n2 a_193_47.n1 4.65
R330 a_193_47.n3 a_193_47.n2 2.685
R331 a_1162_47.n1 a_1162_47.n0 67.2
R332 a_1162_47.n0 a_1162_47.t1 66.666
R333 a_1162_47.n0 a_1162_47.t0 13.143
R334 RESET_B.n0 RESET_B.t1 201.872
R335 RESET_B.n0 RESET_B.t0 172.951
R336 RESET_B RESET_B.n0 78
R337 a_1343_413.t0 a_1343_413.t1 206.38
R338 a_1665_329.t0 a_1665_329.t1 49.25
R339 a_1366_47.t1 a_1366_47.t0 93.059
R340 a_1257_47.n3 a_1257_47.n2 399.793
R341 a_1257_47.n1 a_1257_47.t4 241.535
R342 a_1257_47.n1 a_1257_47.t5 196.547
R343 a_1257_47.n2 a_1257_47.n0 183.436
R344 a_1257_47.n2 a_1257_47.n1 159.918
R345 a_1257_47.n0 a_1257_47.t3 70
R346 a_1257_47.n3 a_1257_47.t2 63.321
R347 a_1257_47.t0 a_1257_47.n3 63.321
R348 a_1257_47.n0 a_1257_47.t1 61.666
C0 VGND SET_B 0.36fF
C1 VGND Q 0.15fF
C2 VGND Q_N 0.21fF
C3 VPWR Q 0.25fF
C4 VPWR Q_N 0.18fF
C5 VPWR VPB 0.27fF
C6 VPWR VGND 0.18fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__dfbbp_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__dfbbp_1 RESET_B VGND CLK SET_B Q VPWR D Q_N VNB VPB
X0 a_788_47.t1 a_942_21.t2 a_648_21.t2 VNB.t7 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1 VPWR.t10 RESET_B.t0 a_942_21.t0 VPB.t14 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X2 VGND.t1 a_1429_21.t4 a_1364_47.t0 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3 VPWR.t2 a_942_21.t3 a_1663_329.t1 VPB.t5 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X4 VPWR.t0 CLK.t0 a_27_47.t0 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X5 a_381_47.t0 D.t0 VPWR.t1 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 VPWR.t11 a_1429_21.t5 a_1341_413.t0 VPB.t17 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7 a_474_413.t3 a_27_47.t2 a_381_47.t3 VNB.t8 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X8 a_1545_47.t1 a_942_21.t4 a_1429_21.t2 VNB.t6 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X9 VPWR.t12 a_1429_21.t6 a_2136_47.t0 VPB.t18 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X10 a_582_47.t0 a_193_47.t2 a_474_413.t0 VNB.t16 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X11 a_1429_21.t3 SET_B.t0 VPWR.t8 VPB.t12 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12 a_648_21.t0 a_474_413.t4 a_788_47.t0 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X13 a_1341_413.t1 a_193_47.t3 a_1255_47.t0 VPB.t15 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14 a_1663_329.t0 a_1255_47.t4 a_1429_21.t0 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X15 a_1160_47.t1 a_648_21.t4 VGND.t7 VNB.t13 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X16 a_193_47.t1 a_27_47.t3 VGND.t5 VNB.t9 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17 a_1255_47.t3 a_27_47.t4 a_1113_329.t1 VPB.t6 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18 Q.t0 a_2136_47.t2 VPWR.t5 VPB.t9 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X19 a_648_21.t3 SET_B.t1 VPWR.t9 VPB.t13 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20 a_788_47.t2 SET_B.t2 VGND.t9 VNB.t14 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21 Q_N.t0 a_1429_21.t7 VPWR.t13 VPB.t19 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X22 VGND.t11 RESET_B.t1 a_942_21.t1 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23 Q.t1 a_2136_47.t3 VGND.t6 VNB.t11 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X24 VPWR.t3 a_942_21.t5 a_892_329.t0 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X25 a_558_413.t1 a_27_47.t5 a_474_413.t2 VPB.t7 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X26 VGND.t8 a_648_21.t5 a_582_47.t1 VNB.t12 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X27 a_892_329.t1 a_474_413.t5 a_648_21.t1 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X28 VGND.t2 a_1429_21.t8 a_2136_47.t1 VNB.t18 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X29 a_193_47.t0 a_27_47.t6 VPWR.t4 VPB.t8 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X30 a_474_413.t1 a_193_47.t4 a_381_47.t2 VPB.t16 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X31 a_1364_47.t1 a_27_47.t7 a_1255_47.t2 VNB.t10 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X32 a_1255_47.t1 a_193_47.t5 a_1160_47.t0 VNB.t17 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X33 Q_N.t1 a_1429_21.t9 VGND.t0 VNB.t19 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X34 a_1545_47.t2 SET_B.t3 VGND.t10 VNB.t15 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X35 VPWR.t6 a_648_21.t6 a_558_413.t0 VPB.t11 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X36 a_381_47.t1 D.t1 VGND.t4 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X37 a_1113_329.t0 a_648_21.t7 VPWR.t7 VPB.t10 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X38 VGND.t3 CLK.t1 a_27_47.t1 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X39 a_1429_21.t1 a_1255_47.t5 a_1545_47.t0 VNB.t5 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
R0 a_942_21.t0 a_942_21.n3 447.663
R1 a_942_21.n1 a_942_21.t4 211.734
R2 a_942_21.n0 a_942_21.t2 210.472
R3 a_942_21.n1 a_942_21.t3 207.402
R4 a_942_21.n0 a_942_21.t5 204.046
R5 a_942_21.n2 a_942_21.t1 189.295
R6 a_942_21.n3 a_942_21.n0 126.544
R7 a_942_21.n2 a_942_21.n1 76
R8 a_942_21.n3 a_942_21.n2 9.774
R9 a_648_21.n5 a_648_21.t5 387.959
R10 a_648_21.n2 a_648_21.t7 299.91
R11 a_648_21.n7 a_648_21.n6 292.5
R12 a_648_21.n2 a_648_21.t4 167.627
R13 a_648_21.n5 a_648_21.t6 143.746
R14 a_648_21.n4 a_648_21.n2 139.816
R15 a_648_21.n6 a_648_21.n5 114.656
R16 a_648_21.n0 a_648_21.t3 110.226
R17 a_648_21.n4 a_648_21.n3 109.954
R18 a_648_21.n6 a_648_21.n4 81.172
R19 a_648_21.t1 a_648_21.n1 63.321
R20 a_648_21.t1 a_648_21.n7 63.321
R21 a_648_21.n3 a_648_21.t2 25.312
R22 a_648_21.n3 a_648_21.t0 25.312
R23 a_648_21.n1 a_648_21.n0 9.38
R24 a_788_47.n0 a_788_47.t1 283.852
R25 a_788_47.t0 a_788_47.n0 49.151
R26 a_788_47.n0 a_788_47.t2 38.571
R27 VNB.t9 VNB.t4 6082.35
R28 VNB.t6 VNB.t3 4595.56
R29 VNB.t7 VNB.t13 4595.56
R30 VNB.t19 VNB.t18 4545.05
R31 VNB VNB.t1 4238.23
R32 VNB.t12 VNB.t14 3558.82
R33 VNB.t17 VNB.t10 3526.47
R34 VNB.t8 VNB.t16 3429.41
R35 VNB.t16 VNB.t12 3105.88
R36 VNB.t15 VNB.t5 3097.97
R37 VNB.t10 VNB.t2 3073.53
R38 VNB.t4 VNB.t8 3073.53
R39 VNB.t2 VNB.t15 2782.35
R40 VNB.t1 VNB.t9 2717.65
R41 VNB.t14 VNB.t0 2349.76
R42 VNB.t18 VNB.t11 2296.7
R43 VNB.t13 VNB.t17 2280.14
R44 VNB.t3 VNB.t19 2248.62
R45 VNB.t5 VNB.t6 2053.33
R46 VNB.t0 VNB.t7 2053.33
R47 RESET_B.n0 RESET_B.t1 208.013
R48 RESET_B.n0 RESET_B.t0 179.092
R49  RESET_B.n0 79.06
R50  RESET_B 2.226
R51 VPWR.n6 VPWR.t2 500.865
R52 VPWR.n1 VPWR.n0 440.25
R53 VPWR.n44 VPWR.t1 374.106
R54 VPWR.n49 VPWR.n48 311.893
R55 VPWR.n36 VPWR.n35 306.984
R56 VPWR.n14 VPWR.n13 292.5
R57 VPWR.n3 VPWR.n2 172.733
R58 VPWR.n28 VPWR.n27 164.214
R59 VPWR.n13 VPWR.t8 91.464
R60 VPWR.n13 VPWR.t11 91.464
R61 VPWR.n35 VPWR.t9 91.464
R62 VPWR.n27 VPWR.t7 86.773
R63 VPWR.n35 VPWR.t6 86.773
R64 VPWR.n0 VPWR.t10 63.101
R65 VPWR.n2 VPWR.t12 58.484
R66 VPWR.n48 VPWR.t4 41.554
R67 VPWR.n48 VPWR.t0 41.554
R68 VPWR.n27 VPWR.t3 38.696
R69 VPWR.n2 VPWR.t5 31.83
R70 VPWR.n0 VPWR.t13 28.032
R71 VPWR.n5 VPWR.n4 4.65
R72 VPWR.n8 VPWR.n7 4.65
R73 VPWR.n10 VPWR.n9 4.65
R74 VPWR.n12 VPWR.n11 4.65
R75 VPWR.n16 VPWR.n15 4.65
R76 VPWR.n18 VPWR.n17 4.65
R77 VPWR.n20 VPWR.n19 4.65
R78 VPWR.n22 VPWR.n21 4.65
R79 VPWR.n24 VPWR.n23 4.65
R80 VPWR.n26 VPWR.n25 4.65
R81 VPWR.n30 VPWR.n29 4.65
R82 VPWR.n32 VPWR.n31 4.65
R83 VPWR.n34 VPWR.n33 4.65
R84 VPWR.n37 VPWR.n36 4.65
R85 VPWR.n39 VPWR.n38 4.65
R86 VPWR.n41 VPWR.n40 4.65
R87 VPWR.n43 VPWR.n42 4.65
R88 VPWR.n45 VPWR.n44 4.65
R89 VPWR.n47 VPWR.n46 4.65
R90 VPWR.n3 VPWR.n1 4.611
R91 VPWR.n50 VPWR.n49 3.932
R92 VPWR.n29 VPWR.n28 3.764
R93 VPWR.n7 VPWR.n6 3.723
R94 VPWR.n15 VPWR.n14 2.327
R95 VPWR.n5 VPWR.n3 0.144
R96 VPWR.n50 VPWR.n47 0.137
R97 VPWR VPWR.n50 0.121
R98 VPWR.n8 VPWR.n5 0.119
R99 VPWR.n10 VPWR.n8 0.119
R100 VPWR.n12 VPWR.n10 0.119
R101 VPWR.n16 VPWR.n12 0.119
R102 VPWR.n18 VPWR.n16 0.119
R103 VPWR.n20 VPWR.n18 0.119
R104 VPWR.n22 VPWR.n20 0.119
R105 VPWR.n24 VPWR.n22 0.119
R106 VPWR.n26 VPWR.n24 0.119
R107 VPWR.n30 VPWR.n26 0.119
R108 VPWR.n32 VPWR.n30 0.119
R109 VPWR.n34 VPWR.n32 0.119
R110 VPWR.n37 VPWR.n34 0.119
R111 VPWR.n39 VPWR.n37 0.119
R112 VPWR.n41 VPWR.n39 0.119
R113 VPWR.n43 VPWR.n41 0.119
R114 VPWR.n45 VPWR.n43 0.119
R115 VPWR.n47 VPWR.n45 0.119
R116 VPB.t5 VPB.t14 585.981
R117 VPB.t19 VPB.t18 556.386
R118 VPB.t8 VPB.t2 556.386
R119 VPB.t10 VPB.t6 426.168
R120 VPB.t4 VPB.t10 405.451
R121 VPB.t7 VPB.t11 355.14
R122 VPB.t15 VPB.t17 349.221
R123 VPB.t17 VPB.t12 319.626
R124 VPB.t13 VPB.t0 319.626
R125 VPB.t11 VPB.t13 313.707
R126 VPB.t14 VPB.t19 287.071
R127 VPB.t12 VPB.t3 284.112
R128 VPB.t18 VPB.t9 281.152
R129 VPB.t2 VPB.t16 275.233
R130 VPB.t6 VPB.t15 248.598
R131 VPB.t0 VPB.t4 248.598
R132 VPB.t16 VPB.t7 248.598
R133 VPB.t1 VPB.t8 248.598
R134 VPB.t3 VPB.t5 213.084
R135 VPB VPB.t1 139.096
R136 a_1429_21.n5 a_1429_21.t4 387.206
R137 a_1429_21.n7 a_1429_21.n6 301.911
R138 a_1429_21.n1 a_1429_21.t7 300.445
R139 a_1429_21.n0 a_1429_21.t6 231.473
R140 a_1429_21.n4 a_1429_21.n2 229.012
R141 a_1429_21.n1 a_1429_21.t9 228.145
R142 a_1429_21.n4 a_1429_21.n3 183.133
R143 a_1429_21.n0 a_1429_21.t8 163.994
R144 a_1429_21.n2 a_1429_21.n0 153.525
R145 a_1429_21.n5 a_1429_21.t5 142.993
R146 a_1429_21.n6 a_1429_21.n5 128.841
R147 a_1429_21.n7 a_1429_21.t3 91.464
R148 a_1429_21.t0 a_1429_21.n7 32.833
R149 a_1429_21.n6 a_1429_21.n4 30.494
R150 a_1429_21.n3 a_1429_21.t2 25.312
R151 a_1429_21.n3 a_1429_21.t1 25.312
R152 a_1429_21.n2 a_1429_21.n1 0.892
R153 a_1364_47.t0 a_1364_47.t1 93.059
R154 VGND.n24 VGND.t7 188.008
R155 VGND.n43 VGND.t4 144.968
R156 VGND.n34 VGND.n33 113.205
R157 VGND.n3 VGND.n0 112.777
R158 VGND.n13 VGND.n12 110.223
R159 VGND.n2 VGND.n1 107.239
R160 VGND.n48 VGND.n47 107.239
R161 VGND.n33 VGND.t8 75.714
R162 VGND.n0 VGND.t2 54.285
R163 VGND.n1 VGND.t11 54.285
R164 VGND.n12 VGND.t1 41.428
R165 VGND.n12 VGND.t10 38.571
R166 VGND.n33 VGND.t9 38.571
R167 VGND.n47 VGND.t5 38.571
R168 VGND.n47 VGND.t3 38.571
R169 VGND.n0 VGND.t6 25.934
R170 VGND.n1 VGND.t0 25.934
R171 VGND.n35 VGND.n34 15.435
R172 VGND.n14 VGND.n13 4.894
R173 VGND.n5 VGND.n4 4.65
R174 VGND.n7 VGND.n6 4.65
R175 VGND.n9 VGND.n8 4.65
R176 VGND.n11 VGND.n10 4.65
R177 VGND.n15 VGND.n14 4.65
R178 VGND.n17 VGND.n16 4.65
R179 VGND.n19 VGND.n18 4.65
R180 VGND.n21 VGND.n20 4.65
R181 VGND.n23 VGND.n22 4.65
R182 VGND.n26 VGND.n25 4.65
R183 VGND.n28 VGND.n27 4.65
R184 VGND.n30 VGND.n29 4.65
R185 VGND.n32 VGND.n31 4.65
R186 VGND.n36 VGND.n35 4.65
R187 VGND.n38 VGND.n37 4.65
R188 VGND.n40 VGND.n39 4.65
R189 VGND.n42 VGND.n41 4.65
R190 VGND.n44 VGND.n43 4.65
R191 VGND.n46 VGND.n45 4.65
R192 VGND.n25 VGND.n24 4.517
R193 VGND.n3 VGND.n2 3.969
R194 VGND.n49 VGND.n48 3.932
R195 VGND.n5 VGND.n3 0.146
R196 VGND.n49 VGND.n46 0.137
R197 VGND VGND.n49 0.121
R198 VGND.n7 VGND.n5 0.119
R199 VGND.n9 VGND.n7 0.119
R200 VGND.n11 VGND.n9 0.119
R201 VGND.n15 VGND.n11 0.119
R202 VGND.n17 VGND.n15 0.119
R203 VGND.n19 VGND.n17 0.119
R204 VGND.n21 VGND.n19 0.119
R205 VGND.n23 VGND.n21 0.119
R206 VGND.n26 VGND.n23 0.119
R207 VGND.n28 VGND.n26 0.119
R208 VGND.n30 VGND.n28 0.119
R209 VGND.n32 VGND.n30 0.119
R210 VGND.n36 VGND.n32 0.119
R211 VGND.n38 VGND.n36 0.119
R212 VGND.n40 VGND.n38 0.119
R213 VGND.n42 VGND.n40 0.119
R214 VGND.n44 VGND.n42 0.119
R215 VGND.n46 VGND.n44 0.119
R216 a_1663_329.t0 a_1663_329.t1 49.25
R217 CLK.n0 CLK.t0 269.919
R218 CLK.n0 CLK.t1 234.573
R219 CLK.n1 CLK.n0 76
R220 CLK CLK.n1 7.571
R221 CLK.n1 CLK 4.687
R222 a_27_47.n0 a_27_47.t7 534.467
R223 a_27_47.n3 a_27_47.t6 263.171
R224 a_27_47.t0 a_27_47.n5 239.261
R225 a_27_47.n1 a_27_47.t2 238.257
R226 a_27_47.n1 a_27_47.t5 231.324
R227 a_27_47.n3 a_27_47.t3 227.825
R228 a_27_47.n4 a_27_47.t1 190.021
R229 a_27_47.n0 a_27_47.t4 137.933
R230 a_27_47.n4 a_27_47.n3 76
R231 a_27_47.n5 a_27_47.n4 35.339
R232 a_27_47.n2 a_27_47.n0 12.947
R233 a_27_47.n5 a_27_47.n2 6.189
R234 a_27_47.n2 a_27_47.n1 4.65
R235 D.n0 D.t0 331.508
R236 D.n0 D.t1 209.401
R237 D.n1 D.n0 76
R238 D.n1 D 8.585
R239 D D.n1 2.029
R240 a_381_47.n1 a_381_47.n0 573.431
R241 a_381_47.n1 a_381_47.t2 84.428
R242 a_381_47.n0 a_381_47.t3 63.333
R243 a_381_47.t0 a_381_47.n1 63.321
R244 a_381_47.n0 a_381_47.t1 29.726
R245 a_1341_413.t0 a_1341_413.t1 206.38
R246 a_474_413.n3 a_474_413.n2 413.812
R247 a_474_413.n1 a_474_413.t4 216.899
R248 a_474_413.n1 a_474_413.t5 210.473
R249 a_474_413.n2 a_474_413.n0 195.144
R250 a_474_413.n2 a_474_413.n1 142.333
R251 a_474_413.n0 a_474_413.t0 63.333
R252 a_474_413.n0 a_474_413.t3 63.333
R253 a_474_413.n3 a_474_413.t2 63.321
R254 a_474_413.t1 a_474_413.n3 63.321
R255 a_1545_47.n0 a_1545_47.t1 274.441
R256 a_1545_47.n0 a_1545_47.t2 64.285
R257 a_1545_47.t0 a_1545_47.n0 49.151
R258 a_2136_47.n0 a_2136_47.t2 239.038
R259 a_2136_47.t0 a_2136_47.n1 237.868
R260 a_2136_47.n0 a_2136_47.t3 166.738
R261 a_2136_47.n1 a_2136_47.t1 150.778
R262 a_2136_47.n1 a_2136_47.n0 99.078
R263 a_193_47.n1 a_193_47.t4 538.588
R264 a_193_47.t0 a_193_47.n3 278.596
R265 a_193_47.n0 a_193_47.t3 267.397
R266 a_193_47.n0 a_193_47.t5 207.297
R267 a_193_47.n3 a_193_47.t1 150.413
R268 a_193_47.n1 a_193_47.t2 135.791
R269 a_193_47.n2 a_193_47.n1 10.055
R270 a_193_47.n2 a_193_47.n0 7.532
R271 a_193_47.n3 a_193_47.n2 6.171
R272 a_582_47.t1 a_582_47.t0 93.516
R273 SET_B.n0 SET_B.t1 397.142
R274 SET_B.n3 SET_B.t0 394.428
R275 SET_B.n0 SET_B.t2 134.984
R276 SET_B.n3 SET_B.t3 134.495
R277 SET_B SET_B.n6 13.6
R278 SET_B.n5 SET_B.n3 13.011
R279 SET_B.n1 SET_B.n0 6.954
R280 SET_B.n6 SET_B.n5 6.318
R281 SET_B.n6 SET_B.n1 2.521
R282 SET_B.n2 SET_B 2.521
R283 SET_B.n6 SET_B.n2 0.775
R284 SET_B.n5 SET_B.n4 0.001
R285 a_1255_47.n3 a_1255_47.n2 399.793
R286 a_1255_47.n1 a_1255_47.t4 241.535
R287 a_1255_47.n1 a_1255_47.t5 196.547
R288 a_1255_47.n2 a_1255_47.n0 183.436
R289 a_1255_47.n2 a_1255_47.n1 159.918
R290 a_1255_47.n0 a_1255_47.t1 70
R291 a_1255_47.t0 a_1255_47.n3 63.321
R292 a_1255_47.n3 a_1255_47.t3 63.321
R293 a_1255_47.n0 a_1255_47.t2 61.666
R294 a_1160_47.n1 a_1160_47.n0 67.2
R295 a_1160_47.n0 a_1160_47.t0 66.666
R296 a_1160_47.n0 a_1160_47.t1 13.143
R297 a_1113_329.t0 a_1113_329.t1 236.868
R298 Q.n1 Q.t0 207.372
R299 Q.n0 Q.t1 117.423
R300 Q Q.n0 66.695
R301 Q.n1 Q 9.019
R302 Q Q.n1 7.458
R303 Q.n0 Q 6.646
R304 Q_N.n1 Q_N.t0 207.566
R305 Q_N.n0 Q_N.t1 117.423
R306 Q_N Q_N.n0 71.502
R307 Q_N.n1 Q_N 8.185
R308 Q_N Q_N.n1 6.859
R309 Q_N.n0 Q_N 5.614
R310 a_892_329.t0 a_892_329.t1 63.321
R311 a_558_413.t0 a_558_413.t1 211.071
C0 VPWR VGND 0.12fF
C1 VGND SET_B 0.36fF
C2 VPWR VPB 0.25fF
C3 VPWR Q 0.14fF
C4 VGND Q_N 0.12fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__dfrbp_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__dfrbp_1 Q Q_N RESET_B D CLK VGND VPWR VNB VPB
X0 Q.t0 a_1283_21.t3 VPWR.t8 VPB.t12 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_1217_47.t0 a_27_47.t2 a_1108_47.t2 VNB.t9 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X2 a_805_47.t1 a_761_289.t4 a_639_47.t1 VNB.t6 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3 VPWR.t7 a_1283_21.t4 a_1847_47.t0 VPB.t11 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X4 a_1108_47.t0 a_193_47.t2 a_761_289.t0 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X5 a_1283_21.t0 a_1108_47.t4 a_1462_47.t0 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 a_651_413.t0 a_27_47.t3 a_543_47.t3 VPB.t8 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7 VGND.t2 RESET_B.t0 a_805_47.t0 VNB.t13 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 VPWR.t2 CLK.t0 a_27_47.t0 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X9 Q_N.t0 a_1847_47.t2 VGND.t4 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 a_448_47.t1 D.t0 VPWR.t1 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11 VGND.t7 a_1283_21.t5 a_1847_47.t1 VNB.t12 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12 a_761_289.t1 a_543_47.t4 VGND.t0 VNB.t5 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X13 Q.t1 a_1283_21.t6 VGND.t8 VNB.t11 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14 a_193_47.t1 a_27_47.t4 VGND.t5 VNB.t8 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15 a_1108_47.t3 a_27_47.t5 a_761_289.t3 VPB.t9 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16 a_543_47.t2 a_27_47.t6 a_448_47.t3 VNB.t7 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X17 a_1462_47.t1 RESET_B.t1 VGND.t3 VNB.t14 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18 a_543_47.t0 a_193_47.t3 a_448_47.t2 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19 a_448_47.t0 D.t1 VGND.t1 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20 VPWR.t6 a_1283_21.t7 a_1270_413.t1 VPB.t10 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21 VPWR.t3 a_1108_47.t5 a_1283_21.t1 VPB.t5 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22 a_1270_413.t0 a_193_47.t4 a_1108_47.t1 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23 a_193_47.t0 a_27_47.t7 VPWR.t4 VPB.t6 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X24 a_1283_21.t2 RESET_B.t2 VPWR.t10 VPB.t14 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X25 VPWR.t9 a_761_289.t5 a_651_413.t2 VPB.t13 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X26 a_639_47.t0 a_193_47.t5 a_543_47.t1 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X27 Q_N.t1 a_1847_47.t3 VPWR.t0 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X28 VGND.t6 a_1283_21.t8 a_1217_47.t1 VNB.t10 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X29 a_651_413.t1 RESET_B.t3 VPWR.t11 VPB.t15 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X30 VGND.t9 CLK.t1 a_27_47.t1 VNB.t15 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X31 a_761_289.t2 a_543_47.t5 VPWR.t5 VPB.t7 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
R0 a_1283_21.n4 a_1283_21.n0 454.156
R1 a_1283_21.n5 a_1283_21.t7 389.181
R2 a_1283_21.n1 a_1283_21.t4 256.987
R3 a_1283_21.n3 a_1283_21.t3 212.079
R4 a_1283_21.n6 a_1283_21.n5 175.164
R5 a_1283_21.n5 a_1283_21.t8 174.888
R6 a_1283_21.n1 a_1283_21.t5 163.801
R7 a_1283_21.n2 a_1283_21.t6 139.779
R8 a_1283_21.t0 a_1283_21.n6 131.071
R9 a_1283_21.n2 a_1283_21.n1 129.263
R10 a_1283_21.n4 a_1283_21.n3 105.942
R11 a_1283_21.n0 a_1283_21.t1 63.321
R12 a_1283_21.n0 a_1283_21.t2 63.321
R13 a_1283_21.n6 a_1283_21.n4 24.698
R14 a_1283_21.n3 a_1283_21.n2 22.639
R15 VPWR.n19 VPWR.t5 514.01
R16 VPWR.n35 VPWR.t1 375.277
R17 VPWR.n11 VPWR.n10 311.956
R18 VPWR.n42 VPWR.n41 311.893
R19 VPWR.n24 VPWR.n23 309.178
R20 VPWR.n5 VPWR.n4 292.5
R21 VPWR.n3 VPWR.n2 292.5
R22 VPWR.n1 VPWR.n0 148.685
R23 VPWR.n10 VPWR.t6 119.607
R24 VPWR.n23 VPWR.t9 93.809
R25 VPWR.n4 VPWR.t3 68.011
R26 VPWR.n10 VPWR.t10 63.321
R27 VPWR.n23 VPWR.t11 63.321
R28 VPWR.n0 VPWR.t7 61.915
R29 VPWR.n41 VPWR.t4 41.554
R30 VPWR.n41 VPWR.t2 41.554
R31 VPWR.n0 VPWR.t0 30.238
R32 VPWR.n2 VPWR.t8 29.315
R33 VPWR.n6 VPWR.n3 5.003
R34 VPWR.n7 VPWR.n6 4.65
R35 VPWR.n9 VPWR.n8 4.65
R36 VPWR.n12 VPWR.n11 4.65
R37 VPWR.n14 VPWR.n13 4.65
R38 VPWR.n16 VPWR.n15 4.65
R39 VPWR.n18 VPWR.n17 4.65
R40 VPWR.n20 VPWR.n19 4.65
R41 VPWR.n22 VPWR.n21 4.65
R42 VPWR.n26 VPWR.n25 4.65
R43 VPWR.n28 VPWR.n27 4.65
R44 VPWR.n30 VPWR.n29 4.65
R45 VPWR.n32 VPWR.n31 4.65
R46 VPWR.n34 VPWR.n33 4.65
R47 VPWR.n36 VPWR.n35 4.65
R48 VPWR.n38 VPWR.n37 4.65
R49 VPWR.n40 VPWR.n39 4.65
R50 VPWR.n6 VPWR.n5 4.072
R51 VPWR.n43 VPWR.n42 3.932
R52 VPWR.n25 VPWR.n24 3.764
R53 VPWR.n7 VPWR.n1 0.143
R54 VPWR.n43 VPWR.n40 0.137
R55 VPWR VPWR.n43 0.123
R56 VPWR.n9 VPWR.n7 0.119
R57 VPWR.n12 VPWR.n9 0.119
R58 VPWR.n14 VPWR.n12 0.119
R59 VPWR.n16 VPWR.n14 0.119
R60 VPWR.n18 VPWR.n16 0.119
R61 VPWR.n20 VPWR.n18 0.119
R62 VPWR.n22 VPWR.n20 0.119
R63 VPWR.n26 VPWR.n22 0.119
R64 VPWR.n28 VPWR.n26 0.119
R65 VPWR.n30 VPWR.n28 0.119
R66 VPWR.n32 VPWR.n30 0.119
R67 VPWR.n34 VPWR.n32 0.119
R68 VPWR.n36 VPWR.n34 0.119
R69 VPWR.n38 VPWR.n36 0.119
R70 VPWR.n40 VPWR.n38 0.119
R71 Q Q.t0 149.239
R72 Q Q.t1 102.342
R73 VPB.t6 VPB.t3 790.186
R74 VPB.t12 VPB.t11 648.13
R75 VPB.t15 VPB.t7 583.021
R76 VPB.t5 VPB.t12 485.358
R77 VPB.t8 VPB.t13 414.33
R78 VPB.t10 VPB.t14 319.626
R79 VPB.t7 VPB.t9 292.99
R80 VPB.t0 VPB.t8 292.99
R81 VPB.t11 VPB.t2 287.071
R82 VPB.t13 VPB.t15 287.071
R83 VPB.t3 VPB.t0 272.274
R84 VPB.t9 VPB.t1 254.517
R85 VPB.t14 VPB.t5 248.598
R86 VPB.t1 VPB.t10 248.598
R87 VPB.t4 VPB.t6 248.598
R88 VPB VPB.t4 192.367
R89 a_27_47.n1 a_27_47.t3 530.008
R90 a_27_47.n0 a_27_47.t5 331.026
R91 a_27_47.t0 a_27_47.n9 271.418
R92 a_27_47.n4 a_27_47.t7 255.459
R93 a_27_47.n6 a_27_47.t4 224.611
R94 a_27_47.n0 a_27_47.t2 204.373
R95 a_27_47.n3 a_27_47.t1 186.535
R96 a_27_47.n1 a_27_47.t6 141.921
R97 a_27_47.n2 a_27_47.n1 90.158
R98 a_27_47.n2 a_27_47.n0 12.643
R99 a_27_47.n7 a_27_47.n6 8.764
R100 a_27_47.n5 a_27_47.n4 7.712
R101 a_27_47.n9 a_27_47.n8 3.339
R102 a_27_47.n6 a_27_47.n5 3.213
R103 a_27_47.n3 a_27_47.n2 3.151
R104 a_27_47.n8 a_27_47.n7 1.391
R105 a_27_47.n7 a_27_47.n3 1.094
R106 a_1108_47.n1 a_1108_47.t4 366.855
R107 a_1108_47.n3 a_1108_47.n2 344.452
R108 a_1108_47.n2 a_1108_47.n0 207.699
R109 a_1108_47.n1 a_1108_47.t5 174.055
R110 a_1108_47.n2 a_1108_47.n1 149.035
R111 a_1108_47.n0 a_1108_47.t0 70
R112 a_1108_47.n3 a_1108_47.t3 68.011
R113 a_1108_47.t1 a_1108_47.n3 63.321
R114 a_1108_47.n0 a_1108_47.t2 61.666
R115 a_1217_47.t1 a_1217_47.t0 94.726
R116 VNB.t8 VNB.t2 8250
R117 VNB VNB.t15 6470.59
R118 VNB.t4 VNB.t6 5370.59
R119 VNB.t3 VNB.t11 5321.88
R120 VNB.t10 VNB.t14 4820.59
R121 VNB.t11 VNB.t12 4545.05
R122 VNB.t13 VNB.t5 3550.91
R123 VNB.t0 VNB.t9 3526.47
R124 VNB.t9 VNB.t10 3105.88
R125 VNB.t7 VNB.t4 3105.88
R126 VNB.t2 VNB.t7 3073.53
R127 VNB.t14 VNB.t3 2944.12
R128 VNB.t15 VNB.t8 2717.65
R129 VNB.t5 VNB.t0 2377.92
R130 VNB.t12 VNB.t1 2345.05
R131 VNB.t6 VNB.t13 2329.41
R132 a_761_289.n3 a_761_289.n2 354.616
R133 a_761_289.n1 a_761_289.t4 350.253
R134 a_761_289.n1 a_761_289.t5 189.586
R135 a_761_289.n2 a_761_289.n1 170.117
R136 a_761_289.n2 a_761_289.n0 167.836
R137 a_761_289.n3 a_761_289.t3 89.119
R138 a_761_289.n0 a_761_289.t0 63.333
R139 a_761_289.t2 a_761_289.n3 41.041
R140 a_761_289.n0 a_761_289.t1 31.979
R141 a_639_47.t1 a_639_47.t0 198.571
R142 a_805_47.t0 a_805_47.t1 60
R143 a_1847_47.t0 a_1847_47.n1 240.007
R144 a_1847_47.n0 a_1847_47.t3 239.038
R145 a_1847_47.n0 a_1847_47.t2 166.738
R146 a_1847_47.n1 a_1847_47.t1 157.454
R147 a_1847_47.n1 a_1847_47.n0 99.66
R148 a_193_47.n0 a_193_47.t2 275.928
R149 a_193_47.n1 a_193_47.t5 258.716
R150 a_193_47.n1 a_193_47.t3 233.933
R151 a_193_47.n3 a_193_47.t1 232.798
R152 a_193_47.n0 a_193_47.t4 145.905
R153 a_193_47.t0 a_193_47.n3 123.515
R154 a_193_47.n2 a_193_47.n0 5.469
R155 a_193_47.n2 a_193_47.n1 4.65
R156 a_193_47.n3 a_193_47.n2 3.654
R157 a_1462_47.t0 a_1462_47.t1 87.142
R158 a_543_47.n3 a_543_47.n2 381.836
R159 a_543_47.n1 a_543_47.t5 332.579
R160 a_543_47.n2 a_543_47.n0 191.51
R161 a_543_47.n2 a_543_47.n1 177.646
R162 a_543_47.n1 a_543_47.t4 168.699
R163 a_543_47.n3 a_543_47.t3 96.154
R164 a_543_47.t0 a_543_47.n3 65.666
R165 a_543_47.n0 a_543_47.t2 65
R166 a_543_47.n0 a_543_47.t1 45
R167 a_651_413.n0 a_651_413.t1 742.814
R168 a_651_413.t0 a_651_413.n0 194.654
R169 a_651_413.n0 a_651_413.t2 63.321
R170 RESET_B.n1 RESET_B.t3 413.312
R171 RESET_B.n4 RESET_B.t2 344.005
R172 RESET_B.n3 RESET_B.t1 187.32
R173 RESET_B.n1 RESET_B.t0 126.126
R174 RESET_B.n2 RESET_B.n1 13.102
R175 RESET_B.n5 RESET_B.n4 9.3
R176 RESET_B.n4 RESET_B.n3 9.159
R177 RESET_B.n2 RESET_B.n0 4.734
R178 RESET_B.n0 RESET_B 4.533
R179 RESET_B.n5 RESET_B.n2 3.214
R180 RESET_B RESET_B.n7 3.113
R181 RESET_B.n7 RESET_B.n6 1.556
R182 RESET_B.n6 RESET_B.n5 1.383
R183 VGND.n35 VGND.t1 215.034
R184 VGND.n1 VGND.t8 154.317
R185 VGND.n2 VGND.n0 128.755
R186 VGND.n10 VGND.n9 116.752
R187 VGND.n20 VGND.n19 107.239
R188 VGND.n40 VGND.n39 107.239
R189 VGND.n9 VGND.t3 100
R190 VGND.n19 VGND.t2 72.857
R191 VGND.n9 VGND.t6 70
R192 VGND.n19 VGND.t0 60.579
R193 VGND.n0 VGND.t7 57.142
R194 VGND.n39 VGND.t5 38.571
R195 VGND.n39 VGND.t9 38.571
R196 VGND.n0 VGND.t4 25.428
R197 VGND.n2 VGND.n1 10.907
R198 VGND.n4 VGND.n3 4.65
R199 VGND.n6 VGND.n5 4.65
R200 VGND.n8 VGND.n7 4.65
R201 VGND.n12 VGND.n11 4.65
R202 VGND.n14 VGND.n13 4.65
R203 VGND.n16 VGND.n15 4.65
R204 VGND.n18 VGND.n17 4.65
R205 VGND.n22 VGND.n21 4.65
R206 VGND.n24 VGND.n23 4.65
R207 VGND.n26 VGND.n25 4.65
R208 VGND.n28 VGND.n27 4.65
R209 VGND.n30 VGND.n29 4.65
R210 VGND.n32 VGND.n31 4.65
R211 VGND.n34 VGND.n33 4.65
R212 VGND.n36 VGND.n35 4.65
R213 VGND.n38 VGND.n37 4.65
R214 VGND.n41 VGND.n40 3.932
R215 VGND.n11 VGND.n10 2.635
R216 VGND.n21 VGND.n20 1.882
R217 VGND.n4 VGND.n2 0.143
R218 VGND.n41 VGND.n38 0.137
R219 VGND VGND.n41 0.123
R220 VGND.n6 VGND.n4 0.119
R221 VGND.n8 VGND.n6 0.119
R222 VGND.n12 VGND.n8 0.119
R223 VGND.n14 VGND.n12 0.119
R224 VGND.n16 VGND.n14 0.119
R225 VGND.n18 VGND.n16 0.119
R226 VGND.n22 VGND.n18 0.119
R227 VGND.n24 VGND.n22 0.119
R228 VGND.n26 VGND.n24 0.119
R229 VGND.n28 VGND.n26 0.119
R230 VGND.n30 VGND.n28 0.119
R231 VGND.n32 VGND.n30 0.119
R232 VGND.n34 VGND.n32 0.119
R233 VGND.n36 VGND.n34 0.119
R234 VGND.n38 VGND.n36 0.119
R235 CLK.n0 CLK.t0 294.554
R236 CLK.n0 CLK.t1 211.008
R237 CLK.n1 CLK.n0 76
R238 CLK.n1 CLK 10.422
R239 CLK CLK.n1 2.011
R240 Q_N Q_N.t1 254.291
R241 Q_N Q_N.t0 144.6
R242 D.n0 D.t1 333.651
R243 D.n0 D.t0 297.233
R244 D D.n0 120.734
R245 a_448_47.n1 a_448_47.n0 541.024
R246 a_448_47.n0 a_448_47.t2 82.083
R247 a_448_47.n1 a_448_47.t3 63.333
R248 a_448_47.n0 a_448_47.t1 63.321
R249 a_448_47.n2 a_448_47.t0 26.393
R250 a_448_47.n3 a_448_47.n2 14.4
R251 a_448_47.n2 a_448_47.n1 3.333
R252 a_1270_413.t0 a_1270_413.t1 126.642
C0 VGND Q 0.12fF
C1 VPWR Q 0.11fF
C2 VPWR VGND 0.12fF
C3 RESET_B VGND 0.37fF
C4 D VPWR 0.11fF
C5 VPWR VPB 0.22fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__dfrbp_2.ext - technology: sky130A

.subckt sky130_fd_sc_hd__dfrbp_2 Q Q_N RESET_B D CLK VGND VPWR VNB VPB
X0 a_1217_47.t0 a_27_47.t2 a_1108_47.t0 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X1 a_805_47.t0 a_761_289.t4 a_639_47.t0 VNB.t9 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 a_1108_47.t2 a_193_47.t2 a_761_289.t3 VNB.t10 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X3 a_1283_21.t1 a_1108_47.t4 a_1462_47.t1 VNB.t17 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 Q_N.t1 a_1659_47.t2 VGND.t5 VNB.t15 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 a_651_413.t2 a_27_47.t3 a_543_47.t1 VPB.t13 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 VGND.t9 RESET_B.t0 a_805_47.t1 VNB.t5 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7 VPWR.t3 a_1283_21.t3 Q.t3 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 VPWR.t10 CLK.t0 a_27_47.t0 VPB.t9 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X9 a_448_47.t2 D.t0 VPWR.t11 VPB.t10 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10 VPWR.t4 a_1283_21.t4 a_1659_47.t0 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X11 a_761_289.t1 a_543_47.t4 VGND.t11 VNB.t7 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X12 VGND.t2 a_1283_21.t5 a_1659_47.t1 VNB.t8 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13 a_193_47.t0 a_27_47.t4 VGND.t8 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14 a_1108_47.t1 a_27_47.t5 a_761_289.t0 VPB.t12 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15 VPWR.t9 a_1659_47.t3 Q_N.t3 VPB.t8 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16 a_543_47.t0 a_27_47.t6 a_448_47.t0 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X17 a_1462_47.t0 RESET_B.t1 VGND.t10 VNB.t6 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18 VGND.t4 a_1659_47.t4 Q_N.t0 VNB.t16 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X19 a_543_47.t2 a_193_47.t3 a_448_47.t3 VPB.t16 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20 a_448_47.t1 D.t1 VGND.t7 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21 VPWR.t5 a_1283_21.t6 a_1270_413.t0 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22 VPWR.t13 a_1108_47.t5 a_1283_21.t2 VPB.t17 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23 a_1270_413.t1 a_193_47.t4 a_1108_47.t3 VPB.t15 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24 a_193_47.t1 a_27_47.t7 VPWR.t12 VPB.t11 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X25 a_1283_21.t0 RESET_B.t2 VPWR.t0 VPB.t14 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X26 Q.t1 a_1283_21.t7 VGND.t1 VNB.t12 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X27 VPWR.t6 a_761_289.t5 a_651_413.t1 VPB.t5 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X28 VGND.t0 a_1283_21.t8 Q.t0 VNB.t13 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X29 Q_N.t2 a_1659_47.t5 VPWR.t8 VPB.t7 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X30 Q.t2 a_1283_21.t9 VPWR.t2 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X31 a_639_47.t1 a_193_47.t5 a_543_47.t3 VNB.t11 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X32 VGND.t3 a_1283_21.t10 a_1217_47.t1 VNB.t14 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X33 a_651_413.t0 RESET_B.t3 VPWR.t1 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X34 VGND.t6 CLK.t1 a_27_47.t1 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X35 a_761_289.t2 a_543_47.t5 VPWR.t7 VPB.t6 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
R0 a_27_47.n1 a_27_47.t3 530.008
R1 a_27_47.n0 a_27_47.t5 331.026
R2 a_27_47.t0 a_27_47.n9 271.418
R3 a_27_47.n4 a_27_47.t7 255.459
R4 a_27_47.n6 a_27_47.t4 224.611
R5 a_27_47.n0 a_27_47.t2 204.373
R6 a_27_47.n3 a_27_47.t1 186.535
R7 a_27_47.n1 a_27_47.t6 141.921
R8 a_27_47.n2 a_27_47.n1 90.158
R9 a_27_47.n2 a_27_47.n0 12.643
R10 a_27_47.n7 a_27_47.n6 8.764
R11 a_27_47.n5 a_27_47.n4 7.712
R12 a_27_47.n9 a_27_47.n8 3.339
R13 a_27_47.n6 a_27_47.n5 3.213
R14 a_27_47.n3 a_27_47.n2 3.151
R15 a_27_47.n8 a_27_47.n7 1.391
R16 a_27_47.n7 a_27_47.n3 1.094
R17 a_1108_47.n1 a_1108_47.t4 366.855
R18 a_1108_47.n3 a_1108_47.n2 344.452
R19 a_1108_47.n2 a_1108_47.n0 207.699
R20 a_1108_47.n1 a_1108_47.t5 174.055
R21 a_1108_47.n2 a_1108_47.n1 149.035
R22 a_1108_47.n0 a_1108_47.t2 70
R23 a_1108_47.t1 a_1108_47.n3 68.011
R24 a_1108_47.n3 a_1108_47.t3 63.321
R25 a_1108_47.n0 a_1108_47.t0 61.666
R26 a_1217_47.t1 a_1217_47.t0 94.726
R27 VNB.t3 VNB.t1 8250
R28 VNB VNB.t0 6470.59
R29 VNB.t17 VNB.t8 6082.35
R30 VNB.t11 VNB.t9 5370.59
R31 VNB.t14 VNB.t6 4820.59
R32 VNB.t5 VNB.t7 3550.91
R33 VNB.t10 VNB.t4 3526.47
R34 VNB.t4 VNB.t14 3105.88
R35 VNB.t2 VNB.t11 3105.88
R36 VNB.t1 VNB.t2 3073.53
R37 VNB.t6 VNB.t17 2944.12
R38 VNB.t0 VNB.t3 2717.65
R39 VNB.t7 VNB.t10 2377.92
R40 VNB.t9 VNB.t5 2329.41
R41 VNB.t8 VNB.t12 2303.7
R42 VNB.t12 VNB.t13 2224.18
R43 VNB.t15 VNB.t16 2030.77
R44 VNB.t13 VNB.t15 2030.77
R45 a_761_289.n3 a_761_289.n2 354.616
R46 a_761_289.n1 a_761_289.t4 350.253
R47 a_761_289.n1 a_761_289.t5 189.586
R48 a_761_289.n2 a_761_289.n1 170.117
R49 a_761_289.n2 a_761_289.n0 167.836
R50 a_761_289.n3 a_761_289.t0 89.119
R51 a_761_289.n0 a_761_289.t3 63.333
R52 a_761_289.t2 a_761_289.n3 41.041
R53 a_761_289.n0 a_761_289.t1 31.979
R54 a_639_47.t0 a_639_47.t1 198.571
R55 a_805_47.t0 a_805_47.t1 60
R56 a_193_47.n0 a_193_47.t2 275.928
R57 a_193_47.n1 a_193_47.t5 258.716
R58 a_193_47.n1 a_193_47.t3 233.933
R59 a_193_47.n3 a_193_47.t0 232.798
R60 a_193_47.n0 a_193_47.t4 145.905
R61 a_193_47.t1 a_193_47.n3 123.515
R62 a_193_47.n2 a_193_47.n0 5.469
R63 a_193_47.n2 a_193_47.n1 4.65
R64 a_193_47.n3 a_193_47.n2 3.654
R65 a_1462_47.t0 a_1462_47.t1 87.142
R66 a_1283_21.n6 a_1283_21.n5 403.181
R67 a_1283_21.n3 a_1283_21.t6 389.181
R68 a_1283_21.n2 a_1283_21.t4 257.066
R69 a_1283_21.n0 a_1283_21.t3 212.079
R70 a_1283_21.n1 a_1283_21.t9 212.079
R71 a_1283_21.n4 a_1283_21.n3 178.364
R72 a_1283_21.n2 a_1283_21.t5 176.733
R73 a_1283_21.n3 a_1283_21.t10 174.888
R74 a_1283_21.n0 a_1283_21.t8 139.779
R75 a_1283_21.n1 a_1283_21.t7 139.779
R76 a_1283_21.n4 a_1283_21.t1 131.071
R77 a_1283_21.n5 a_1283_21.n2 113.818
R78 a_1283_21.n2 a_1283_21.n1 70.839
R79 a_1283_21.n1 a_1283_21.n0 67.187
R80 a_1283_21.n6 a_1283_21.t2 63.321
R81 a_1283_21.t0 a_1283_21.n6 63.321
R82 a_1283_21.n5 a_1283_21.n4 55.017
R83 a_1659_47.t0 a_1659_47.n2 239.157
R84 a_1659_47.n2 a_1659_47.t1 238.53
R85 a_1659_47.n1 a_1659_47.t5 212.079
R86 a_1659_47.n0 a_1659_47.t3 212.079
R87 a_1659_47.n2 a_1659_47.n1 187.917
R88 a_1659_47.n1 a_1659_47.t2 139.779
R89 a_1659_47.n0 a_1659_47.t4 139.779
R90 a_1659_47.n1 a_1659_47.n0 61.345
R91 VGND.n42 VGND.t7 215.034
R92 VGND.n1 VGND.n0 128.641
R93 VGND.n2 VGND.t4 119.488
R94 VGND.n17 VGND.n16 116.752
R95 VGND.n6 VGND.n5 113.197
R96 VGND.n27 VGND.n26 107.239
R97 VGND.n47 VGND.n46 107.239
R98 VGND.n16 VGND.t10 100
R99 VGND.n26 VGND.t9 72.857
R100 VGND.n16 VGND.t3 70
R101 VGND.n26 VGND.t11 60.579
R102 VGND.n5 VGND.t2 57.142
R103 VGND.n46 VGND.t8 38.571
R104 VGND.n46 VGND.t6 38.571
R105 VGND.n5 VGND.t1 25.428
R106 VGND.n0 VGND.t5 24.923
R107 VGND.n0 VGND.t0 24.923
R108 VGND.n2 VGND.n1 11.878
R109 VGND.n4 VGND.n3 4.65
R110 VGND.n7 VGND.n6 4.65
R111 VGND.n9 VGND.n8 4.65
R112 VGND.n11 VGND.n10 4.65
R113 VGND.n13 VGND.n12 4.65
R114 VGND.n15 VGND.n14 4.65
R115 VGND.n19 VGND.n18 4.65
R116 VGND.n21 VGND.n20 4.65
R117 VGND.n23 VGND.n22 4.65
R118 VGND.n25 VGND.n24 4.65
R119 VGND.n29 VGND.n28 4.65
R120 VGND.n31 VGND.n30 4.65
R121 VGND.n33 VGND.n32 4.65
R122 VGND.n35 VGND.n34 4.65
R123 VGND.n37 VGND.n36 4.65
R124 VGND.n39 VGND.n38 4.65
R125 VGND.n41 VGND.n40 4.65
R126 VGND.n43 VGND.n42 4.65
R127 VGND.n45 VGND.n44 4.65
R128 VGND.n48 VGND.n47 3.932
R129 VGND.n18 VGND.n17 2.635
R130 VGND.n28 VGND.n27 1.882
R131 VGND.n4 VGND.n2 0.301
R132 VGND.n48 VGND.n45 0.137
R133 VGND VGND.n48 0.123
R134 VGND.n7 VGND.n4 0.119
R135 VGND.n9 VGND.n7 0.119
R136 VGND.n11 VGND.n9 0.119
R137 VGND.n13 VGND.n11 0.119
R138 VGND.n15 VGND.n13 0.119
R139 VGND.n19 VGND.n15 0.119
R140 VGND.n21 VGND.n19 0.119
R141 VGND.n23 VGND.n21 0.119
R142 VGND.n25 VGND.n23 0.119
R143 VGND.n29 VGND.n25 0.119
R144 VGND.n31 VGND.n29 0.119
R145 VGND.n33 VGND.n31 0.119
R146 VGND.n35 VGND.n33 0.119
R147 VGND.n37 VGND.n35 0.119
R148 VGND.n39 VGND.n37 0.119
R149 VGND.n41 VGND.n39 0.119
R150 VGND.n43 VGND.n41 0.119
R151 VGND.n45 VGND.n43 0.119
R152 Q_N Q_N.n0 138.494
R153 Q_N Q_N.n1 73.268
R154 Q_N.n0 Q_N.t3 26.595
R155 Q_N.n0 Q_N.t2 26.595
R156 Q_N.n1 Q_N.t0 24.923
R157 Q_N.n1 Q_N.t1 24.923
R158 a_543_47.n3 a_543_47.n2 381.836
R159 a_543_47.n1 a_543_47.t5 332.579
R160 a_543_47.n2 a_543_47.n0 191.51
R161 a_543_47.n2 a_543_47.n1 177.646
R162 a_543_47.n1 a_543_47.t4 168.699
R163 a_543_47.t1 a_543_47.n3 96.154
R164 a_543_47.n3 a_543_47.t2 65.666
R165 a_543_47.n0 a_543_47.t0 65
R166 a_543_47.n0 a_543_47.t3 45
R167 a_651_413.t0 a_651_413.n0 742.814
R168 a_651_413.n0 a_651_413.t2 194.654
R169 a_651_413.n0 a_651_413.t1 63.321
R170 VPB.t11 VPB.t10 790.186
R171 VPB.t4 VPB.t6 583.021
R172 VPB.t17 VPB.t2 577.102
R173 VPB.t13 VPB.t5 414.33
R174 VPB.t1 VPB.t14 319.626
R175 VPB.t6 VPB.t12 292.99
R176 VPB.t16 VPB.t13 292.99
R177 VPB.t2 VPB.t0 287.071
R178 VPB.t5 VPB.t4 287.071
R179 VPB.t0 VPB.t3 272.274
R180 VPB.t10 VPB.t16 272.274
R181 VPB.t12 VPB.t15 254.517
R182 VPB.t7 VPB.t8 248.598
R183 VPB.t3 VPB.t7 248.598
R184 VPB.t14 VPB.t17 248.598
R185 VPB.t15 VPB.t1 248.598
R186 VPB.t9 VPB.t11 248.598
R187 VPB VPB.t9 192.367
R188 RESET_B.n1 RESET_B.t3 413.312
R189 RESET_B.n4 RESET_B.t2 344.005
R190 RESET_B.n3 RESET_B.t1 187.32
R191 RESET_B.n1 RESET_B.t0 126.126
R192 RESET_B.n2 RESET_B.n1 13.102
R193 RESET_B.n5 RESET_B.n4 9.3
R194 RESET_B.n4 RESET_B.n3 9.159
R195 RESET_B.n2 RESET_B.n0 4.734
R196 RESET_B.n0 RESET_B 4.533
R197 RESET_B.n5 RESET_B.n2 3.214
R198 RESET_B RESET_B.n7 3.113
R199 RESET_B.n7 RESET_B.n6 1.556
R200 RESET_B.n6 RESET_B.n5 1.383
R201 Q Q.n0 313.323
R202 Q Q.n1 109.12
R203 Q.n0 Q.t3 34.475
R204 Q.n1 Q.t0 32.307
R205 Q.n0 Q.t2 26.595
R206 Q.n1 Q.t1 24.923
R207 VPWR.n23 VPWR.t7 514.01
R208 VPWR.n39 VPWR.t11 375.277
R209 VPWR.n10 VPWR.t13 374.609
R210 VPWR.n15 VPWR.n14 311.956
R211 VPWR.n46 VPWR.n45 311.893
R212 VPWR.n28 VPWR.n27 309.178
R213 VPWR.n6 VPWR.n5 308.688
R214 VPWR.n1 VPWR.n0 307.239
R215 VPWR.n2 VPWR.t9 179.026
R216 VPWR.n14 VPWR.t5 119.607
R217 VPWR.n27 VPWR.t6 93.809
R218 VPWR.n14 VPWR.t0 63.321
R219 VPWR.n27 VPWR.t1 63.321
R220 VPWR.n5 VPWR.t4 61.562
R221 VPWR.n45 VPWR.t12 41.554
R222 VPWR.n45 VPWR.t10 41.554
R223 VPWR.n5 VPWR.t2 31.012
R224 VPWR.n0 VPWR.t8 26.595
R225 VPWR.n0 VPWR.t3 26.595
R226 VPWR.n4 VPWR.n3 4.65
R227 VPWR.n7 VPWR.n6 4.65
R228 VPWR.n9 VPWR.n8 4.65
R229 VPWR.n11 VPWR.n10 4.65
R230 VPWR.n13 VPWR.n12 4.65
R231 VPWR.n16 VPWR.n15 4.65
R232 VPWR.n18 VPWR.n17 4.65
R233 VPWR.n20 VPWR.n19 4.65
R234 VPWR.n22 VPWR.n21 4.65
R235 VPWR.n24 VPWR.n23 4.65
R236 VPWR.n26 VPWR.n25 4.65
R237 VPWR.n30 VPWR.n29 4.65
R238 VPWR.n32 VPWR.n31 4.65
R239 VPWR.n34 VPWR.n33 4.65
R240 VPWR.n36 VPWR.n35 4.65
R241 VPWR.n38 VPWR.n37 4.65
R242 VPWR.n40 VPWR.n39 4.65
R243 VPWR.n42 VPWR.n41 4.65
R244 VPWR.n44 VPWR.n43 4.65
R245 VPWR.n47 VPWR.n46 3.932
R246 VPWR.n2 VPWR.n1 3.895
R247 VPWR.n29 VPWR.n28 3.764
R248 VPWR.n4 VPWR.n2 0.321
R249 VPWR.n47 VPWR.n44 0.137
R250 VPWR VPWR.n47 0.123
R251 VPWR.n7 VPWR.n4 0.119
R252 VPWR.n9 VPWR.n7 0.119
R253 VPWR.n11 VPWR.n9 0.119
R254 VPWR.n13 VPWR.n11 0.119
R255 VPWR.n16 VPWR.n13 0.119
R256 VPWR.n18 VPWR.n16 0.119
R257 VPWR.n20 VPWR.n18 0.119
R258 VPWR.n22 VPWR.n20 0.119
R259 VPWR.n24 VPWR.n22 0.119
R260 VPWR.n26 VPWR.n24 0.119
R261 VPWR.n30 VPWR.n26 0.119
R262 VPWR.n32 VPWR.n30 0.119
R263 VPWR.n34 VPWR.n32 0.119
R264 VPWR.n36 VPWR.n34 0.119
R265 VPWR.n38 VPWR.n36 0.119
R266 VPWR.n40 VPWR.n38 0.119
R267 VPWR.n42 VPWR.n40 0.119
R268 VPWR.n44 VPWR.n42 0.119
R269 CLK.n0 CLK.t0 294.554
R270 CLK.n0 CLK.t1 211.008
R271 CLK.n1 CLK.n0 76
R272 CLK.n1 CLK 10.422
R273 CLK CLK.n1 2.011
R274 D.n0 D.t1 333.651
R275 D.n0 D.t0 297.233
R276 D D.n0 120.734
R277 a_448_47.n1 a_448_47.n0 541.024
R278 a_448_47.n0 a_448_47.t3 82.083
R279 a_448_47.n1 a_448_47.t0 63.333
R280 a_448_47.n0 a_448_47.t2 63.321
R281 a_448_47.n2 a_448_47.t1 26.393
R282 a_448_47.n3 a_448_47.n2 14.4
R283 a_448_47.n2 a_448_47.n1 3.333
R284 a_1270_413.t0 a_1270_413.t1 126.642
C0 VGND RESET_B 0.37fF
C1 VPWR D 0.11fF
C2 VPWR VPB 0.23fF
C3 VGND Q_N 0.24fF
C4 VPWR Q_N 0.24fF
C5 VGND Q 0.15fF
C6 VPWR VGND 0.14fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__dfrtn_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__dfrtn_1 CLK_N Q RESET_B D VGND VPWR VNB VPB
X0 a_1217_47.t0 a_193_47.t2 a_1108_47.t1 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X1 a_805_47.t0 a_761_289.t4 a_639_47.t0 VNB.t7 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 a_1108_47.t2 a_27_47.t2 a_761_289.t3 VNB.t8 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X3 a_1283_21.t0 a_1108_47.t4 a_1462_47.t0 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 a_651_413.t0 a_193_47.t3 a_543_47.t1 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 VGND.t5 RESET_B.t0 a_805_47.t1 VNB.t12 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 Q.t1 a_1283_21.t3 VPWR.t1 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 VPWR.t2 CLK_N.t0 a_27_47.t0 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X8 a_448_47.t1 D.t0 VPWR.t9 VPB.t13 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9 a_761_289.t0 a_543_47.t4 VGND.t6 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X10 a_193_47.t0 a_27_47.t3 VGND.t3 VNB.t9 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11 a_1108_47.t0 a_193_47.t4 a_761_289.t2 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12 a_543_47.t0 a_193_47.t5 a_448_47.t2 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X13 a_1462_47.t1 RESET_B.t1 VGND.t4 VNB.t13 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14 a_543_47.t3 a_27_47.t4 a_448_47.t3 VPB.t7 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15 a_448_47.t0 D.t1 VGND.t7 VNB.t11 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16 VPWR.t0 a_1283_21.t4 a_1270_413.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17 VPWR.t4 a_1108_47.t5 a_1283_21.t1 VPB.t8 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18 a_1270_413.t1 a_27_47.t5 a_1108_47.t3 VPB.t6 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19 a_193_47.t1 a_27_47.t6 VPWR.t3 VPB.t5 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X20 a_1283_21.t2 RESET_B.t2 VPWR.t5 VPB.t10 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21 VPWR.t7 a_761_289.t5 a_651_413.t1 VPB.t9 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22 Q.t0 a_1283_21.t5 VGND.t0 VNB.t5 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X23 a_639_47.t1 a_27_47.t7 a_543_47.t2 VNB.t10 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X24 VGND.t1 a_1283_21.t6 a_1217_47.t1 VNB.t6 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X25 a_651_413.t2 RESET_B.t3 VPWR.t6 VPB.t11 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X26 VGND.t2 CLK_N.t1 a_27_47.t1 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X27 a_761_289.t1 a_543_47.t5 VPWR.t8 VPB.t12 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
R0 a_193_47.n1 a_193_47.t3 530.008
R1 a_193_47.n0 a_193_47.t4 331.026
R2 a_193_47.t1 a_193_47.n3 274.937
R3 a_193_47.n0 a_193_47.t2 204.373
R4 a_193_47.n3 a_193_47.t0 182.271
R5 a_193_47.n1 a_193_47.t5 141.921
R6 a_193_47.n2 a_193_47.n1 90.158
R7 a_193_47.n2 a_193_47.n0 12.643
R8 a_193_47.n3 a_193_47.n2 5.823
R9 a_1108_47.n1 a_1108_47.t4 366.855
R10 a_1108_47.n3 a_1108_47.n2 344.452
R11 a_1108_47.n2 a_1108_47.n0 207.699
R12 a_1108_47.n1 a_1108_47.t5 174.055
R13 a_1108_47.n2 a_1108_47.n1 149.035
R14 a_1108_47.n0 a_1108_47.t2 70
R15 a_1108_47.t0 a_1108_47.n3 68.011
R16 a_1108_47.n3 a_1108_47.t3 63.321
R17 a_1108_47.n0 a_1108_47.t1 61.666
R18 a_1217_47.t1 a_1217_47.t0 94.726
R19 VNB.t9 VNB.t11 8250
R20 VNB VNB.t1 6470.59
R21 VNB.t4 VNB.t5 5985.29
R22 VNB.t10 VNB.t7 5370.59
R23 VNB.t6 VNB.t13 4820.59
R24 VNB.t12 VNB.t0 3550.91
R25 VNB.t8 VNB.t3 3526.47
R26 VNB.t3 VNB.t6 3105.88
R27 VNB.t2 VNB.t10 3105.88
R28 VNB.t11 VNB.t2 3073.53
R29 VNB.t13 VNB.t4 2944.12
R30 VNB.t1 VNB.t9 2717.65
R31 VNB.t0 VNB.t8 2377.92
R32 VNB.t7 VNB.t12 2329.41
R33 a_761_289.n3 a_761_289.n2 354.616
R34 a_761_289.n1 a_761_289.t4 350.253
R35 a_761_289.n1 a_761_289.t5 189.586
R36 a_761_289.n2 a_761_289.n1 170.117
R37 a_761_289.n2 a_761_289.n0 167.836
R38 a_761_289.n3 a_761_289.t2 89.119
R39 a_761_289.n0 a_761_289.t3 63.333
R40 a_761_289.t1 a_761_289.n3 41.041
R41 a_761_289.n0 a_761_289.t0 31.979
R42 a_639_47.t0 a_639_47.t1 198.571
R43 a_805_47.t0 a_805_47.t1 60
R44 a_27_47.n0 a_27_47.t2 275.928
R45 a_27_47.n3 a_27_47.t6 263.171
R46 a_27_47.n1 a_27_47.t7 258.716
R47 a_27_47.t0 a_27_47.n5 239.418
R48 a_27_47.n1 a_27_47.t4 233.933
R49 a_27_47.n3 a_27_47.t3 227.825
R50 a_27_47.n4 a_27_47.t1 190.224
R51 a_27_47.n0 a_27_47.t5 145.905
R52 a_27_47.n4 a_27_47.n3 76
R53 a_27_47.n5 a_27_47.n4 35.339
R54 a_27_47.n5 a_27_47.n2 6.556
R55 a_27_47.n2 a_27_47.n0 5.469
R56 a_27_47.n2 a_27_47.n1 4.65
R57 a_1462_47.t0 a_1462_47.t1 87.142
R58 a_1283_21.n2 a_1283_21.n0 515.369
R59 a_1283_21.n3 a_1283_21.t4 389.181
R60 a_1283_21.n1 a_1283_21.t3 239.038
R61 a_1283_21.n4 a_1283_21.n3 175.164
R62 a_1283_21.n3 a_1283_21.t6 174.888
R63 a_1283_21.n1 a_1283_21.t5 166.738
R64 a_1283_21.t0 a_1283_21.n4 131.071
R65 a_1283_21.n2 a_1283_21.n1 88.16
R66 a_1283_21.n0 a_1283_21.t1 63.321
R67 a_1283_21.n0 a_1283_21.t2 63.321
R68 a_1283_21.n4 a_1283_21.n2 37.718
R69 a_543_47.n3 a_543_47.n2 381.836
R70 a_543_47.n1 a_543_47.t5 332.579
R71 a_543_47.n2 a_543_47.n0 191.51
R72 a_543_47.n2 a_543_47.n1 177.646
R73 a_543_47.n1 a_543_47.t4 168.699
R74 a_543_47.t1 a_543_47.n3 96.154
R75 a_543_47.n3 a_543_47.t3 65.666
R76 a_543_47.n0 a_543_47.t0 65
R77 a_543_47.n0 a_543_47.t2 45
R78 a_651_413.n0 a_651_413.t2 742.814
R79 a_651_413.t0 a_651_413.n0 194.654
R80 a_651_413.n0 a_651_413.t1 63.321
R81 VPB.t5 VPB.t13 790.186
R82 VPB.t8 VPB.t1 636.292
R83 VPB.t11 VPB.t12 583.021
R84 VPB.t4 VPB.t9 414.33
R85 VPB.t0 VPB.t10 319.626
R86 VPB.t12 VPB.t3 292.99
R87 VPB.t7 VPB.t4 292.99
R88 VPB.t9 VPB.t11 287.071
R89 VPB.t13 VPB.t7 272.274
R90 VPB.t3 VPB.t6 254.517
R91 VPB.t10 VPB.t8 248.598
R92 VPB.t6 VPB.t0 248.598
R93 VPB.t2 VPB.t5 248.598
R94 VPB VPB.t2 192.367
R95 RESET_B.n1 RESET_B.t3 413.312
R96 RESET_B.n4 RESET_B.t2 344.005
R97 RESET_B.n3 RESET_B.t1 187.32
R98 RESET_B.n1 RESET_B.t0 126.126
R99 RESET_B.n2 RESET_B.n1 13.102
R100 RESET_B.n5 RESET_B.n4 9.3
R101 RESET_B.n4 RESET_B.n3 9.159
R102 RESET_B.n2 RESET_B.n0 4.734
R103 RESET_B.n0 RESET_B 4.533
R104 RESET_B.n5 RESET_B.n2 3.214
R105 RESET_B RESET_B.n7 3.113
R106 RESET_B.n7 RESET_B.n6 1.556
R107 RESET_B.n6 RESET_B.n5 1.383
R108 VGND.n27 VGND.t7 215.034
R109 VGND.n0 VGND.t0 138.166
R110 VGND.n2 VGND.n1 116.752
R111 VGND.n12 VGND.n11 107.239
R112 VGND.n32 VGND.n31 107.239
R113 VGND.n1 VGND.t4 100
R114 VGND.n11 VGND.t5 72.857
R115 VGND.n1 VGND.t1 70
R116 VGND.n11 VGND.t6 60.579
R117 VGND.n31 VGND.t3 38.571
R118 VGND.n31 VGND.t2 38.571
R119 VGND.n4 VGND.n3 4.65
R120 VGND.n6 VGND.n5 4.65
R121 VGND.n8 VGND.n7 4.65
R122 VGND.n10 VGND.n9 4.65
R123 VGND.n14 VGND.n13 4.65
R124 VGND.n16 VGND.n15 4.65
R125 VGND.n18 VGND.n17 4.65
R126 VGND.n20 VGND.n19 4.65
R127 VGND.n22 VGND.n21 4.65
R128 VGND.n24 VGND.n23 4.65
R129 VGND.n26 VGND.n25 4.65
R130 VGND.n28 VGND.n27 4.65
R131 VGND.n30 VGND.n29 4.65
R132 VGND.n33 VGND.n32 3.932
R133 VGND.n3 VGND.n2 2.635
R134 VGND.n13 VGND.n12 1.882
R135 VGND.n4 VGND.n0 0.14
R136 VGND.n33 VGND.n30 0.137
R137 VGND VGND.n33 0.123
R138 VGND.n6 VGND.n4 0.119
R139 VGND.n8 VGND.n6 0.119
R140 VGND.n10 VGND.n8 0.119
R141 VGND.n14 VGND.n10 0.119
R142 VGND.n16 VGND.n14 0.119
R143 VGND.n18 VGND.n16 0.119
R144 VGND.n20 VGND.n18 0.119
R145 VGND.n22 VGND.n20 0.119
R146 VGND.n24 VGND.n22 0.119
R147 VGND.n26 VGND.n24 0.119
R148 VGND.n28 VGND.n26 0.119
R149 VGND.n30 VGND.n28 0.119
R150 VPWR.n13 VPWR.t8 514.01
R151 VPWR.n29 VPWR.t9 375.277
R152 VPWR.n0 VPWR.t4 375.25
R153 VPWR.n5 VPWR.n4 311.956
R154 VPWR.n36 VPWR.n35 311.893
R155 VPWR.n18 VPWR.n17 309.178
R156 VPWR.n1 VPWR.t1 200.298
R157 VPWR.n4 VPWR.t0 119.607
R158 VPWR.n17 VPWR.t7 93.809
R159 VPWR.n4 VPWR.t5 63.321
R160 VPWR.n17 VPWR.t6 63.321
R161 VPWR.n35 VPWR.t3 41.554
R162 VPWR.n35 VPWR.t2 41.554
R163 VPWR.n3 VPWR.n2 4.65
R164 VPWR.n6 VPWR.n5 4.65
R165 VPWR.n8 VPWR.n7 4.65
R166 VPWR.n10 VPWR.n9 4.65
R167 VPWR.n12 VPWR.n11 4.65
R168 VPWR.n14 VPWR.n13 4.65
R169 VPWR.n16 VPWR.n15 4.65
R170 VPWR.n20 VPWR.n19 4.65
R171 VPWR.n22 VPWR.n21 4.65
R172 VPWR.n24 VPWR.n23 4.65
R173 VPWR.n26 VPWR.n25 4.65
R174 VPWR.n28 VPWR.n27 4.65
R175 VPWR.n30 VPWR.n29 4.65
R176 VPWR.n32 VPWR.n31 4.65
R177 VPWR.n34 VPWR.n33 4.65
R178 VPWR.n1 VPWR.n0 4.195
R179 VPWR.n37 VPWR.n36 3.932
R180 VPWR.n19 VPWR.n18 3.764
R181 VPWR.n3 VPWR.n1 0.683
R182 VPWR.n37 VPWR.n34 0.137
R183 VPWR VPWR.n37 0.123
R184 VPWR.n6 VPWR.n3 0.119
R185 VPWR.n8 VPWR.n6 0.119
R186 VPWR.n10 VPWR.n8 0.119
R187 VPWR.n12 VPWR.n10 0.119
R188 VPWR.n14 VPWR.n12 0.119
R189 VPWR.n16 VPWR.n14 0.119
R190 VPWR.n20 VPWR.n16 0.119
R191 VPWR.n22 VPWR.n20 0.119
R192 VPWR.n24 VPWR.n22 0.119
R193 VPWR.n26 VPWR.n24 0.119
R194 VPWR.n28 VPWR.n26 0.119
R195 VPWR.n30 VPWR.n28 0.119
R196 VPWR.n32 VPWR.n30 0.119
R197 VPWR.n34 VPWR.n32 0.119
R198 Q.n1 Q.t1 207.309
R199 Q.n0 Q.t0 117.423
R200 Q Q.n0 47.901
R201 Q.n0 Q 10.29
R202 Q.n1 Q 9.192
R203 Q Q.n1 7.602
R204 CLK_N.n0 CLK_N.t0 294.554
R205 CLK_N.n0 CLK_N.t1 211.008
R206 CLK_N CLK_N.n0 77.87
R207 D.n0 D.t1 333.651
R208 D.n0 D.t0 297.233
R209 D D.n0 120.734
R210 a_448_47.n1 a_448_47.n0 541.024
R211 a_448_47.n0 a_448_47.t3 82.083
R212 a_448_47.n1 a_448_47.t2 63.333
R213 a_448_47.n0 a_448_47.t1 63.321
R214 a_448_47.n2 a_448_47.t0 26.393
R215 a_448_47.n3 a_448_47.n2 14.4
R216 a_448_47.n2 a_448_47.n1 3.333
R217 a_1270_413.t0 a_1270_413.t1 126.642
C0 VPWR Q 0.13fF
C1 RESET_B VGND 0.37fF
C2 VPWR VPB 0.19fF
C3 D VPWR 0.11fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__dfrtp_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__dfrtp_1 Q RESET_B D CLK VGND VPWR VNB VPB
X0 a_1217_47.t0 a_27_47.t2 a_1108_47.t0 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X1 a_805_47.t0 a_761_289.t4 a_639_47.t0 VNB.t11 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 a_1108_47.t2 a_193_47.t2 a_761_289.t1 VNB.t9 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X3 a_1283_21.t0 a_1108_47.t4 a_1462_47.t0 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 a_651_413.t1 a_27_47.t3 a_543_47.t2 VPB.t10 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 VGND.t5 RESET_B.t0 a_805_47.t1 VNB.t7 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 Q.t0 a_1283_21.t3 VPWR.t4 VPB.t6 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 VPWR.t7 CLK.t0 a_27_47.t1 VPB.t11 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X8 a_448_47.t1 D.t0 VPWR.t1 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9 a_761_289.t2 a_543_47.t4 VGND.t1 VNB.t12 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X10 a_193_47.t0 a_27_47.t4 VGND.t4 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11 a_1108_47.t1 a_27_47.t5 a_761_289.t0 VPB.t9 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12 a_543_47.t3 a_27_47.t6 a_448_47.t3 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X13 a_1462_47.t1 RESET_B.t1 VGND.t6 VNB.t8 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14 a_543_47.t1 a_193_47.t3 a_448_47.t0 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15 a_448_47.t2 D.t1 VGND.t7 VNB.t13 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16 VPWR.t3 a_1283_21.t4 a_1270_413.t1 VPB.t5 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17 VPWR.t5 a_1108_47.t5 a_1283_21.t1 VPB.t7 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18 a_1270_413.t0 a_193_47.t4 a_1108_47.t3 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19 a_193_47.t1 a_27_47.t7 VPWR.t6 VPB.t8 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X20 a_1283_21.t2 RESET_B.t2 VPWR.t8 VPB.t12 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21 VPWR.t0 a_761_289.t5 a_651_413.t0 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22 Q.t1 a_1283_21.t5 VGND.t3 VNB.t5 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X23 a_639_47.t1 a_193_47.t5 a_543_47.t0 VNB.t10 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X24 VGND.t2 a_1283_21.t6 a_1217_47.t1 VNB.t6 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X25 a_651_413.t2 RESET_B.t3 VPWR.t9 VPB.t13 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X26 VGND.t0 CLK.t1 a_27_47.t0 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X27 a_761_289.t3 a_543_47.t5 VPWR.t2 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
R0 a_27_47.n1 a_27_47.t3 530.008
R1 a_27_47.n0 a_27_47.t5 331.026
R2 a_27_47.t1 a_27_47.n9 271.418
R3 a_27_47.n4 a_27_47.t7 255.459
R4 a_27_47.n6 a_27_47.t4 224.611
R5 a_27_47.n0 a_27_47.t2 204.373
R6 a_27_47.n3 a_27_47.t0 186.535
R7 a_27_47.n1 a_27_47.t6 141.921
R8 a_27_47.n2 a_27_47.n1 90.158
R9 a_27_47.n2 a_27_47.n0 12.643
R10 a_27_47.n7 a_27_47.n6 8.764
R11 a_27_47.n5 a_27_47.n4 7.712
R12 a_27_47.n9 a_27_47.n8 3.339
R13 a_27_47.n6 a_27_47.n5 3.213
R14 a_27_47.n3 a_27_47.n2 3.151
R15 a_27_47.n8 a_27_47.n7 1.391
R16 a_27_47.n7 a_27_47.n3 1.094
R17 a_1108_47.n1 a_1108_47.t4 366.855
R18 a_1108_47.n3 a_1108_47.n2 344.452
R19 a_1108_47.n2 a_1108_47.n0 207.699
R20 a_1108_47.n1 a_1108_47.t5 174.055
R21 a_1108_47.n2 a_1108_47.n1 149.035
R22 a_1108_47.n0 a_1108_47.t2 70
R23 a_1108_47.t1 a_1108_47.n3 68.011
R24 a_1108_47.n3 a_1108_47.t3 63.321
R25 a_1108_47.n0 a_1108_47.t0 61.666
R26 a_1217_47.t1 a_1217_47.t0 94.726
R27 VNB.t3 VNB.t13 8250
R28 VNB VNB.t0 6470.59
R29 VNB.t1 VNB.t5 5985.29
R30 VNB.t10 VNB.t11 5370.59
R31 VNB.t6 VNB.t8 4820.59
R32 VNB.t7 VNB.t12 3550.91
R33 VNB.t9 VNB.t4 3526.47
R34 VNB.t4 VNB.t6 3105.88
R35 VNB.t2 VNB.t10 3105.88
R36 VNB.t13 VNB.t2 3073.53
R37 VNB.t8 VNB.t1 2944.12
R38 VNB.t0 VNB.t3 2717.65
R39 VNB.t12 VNB.t9 2377.92
R40 VNB.t11 VNB.t7 2329.41
R41 a_761_289.n3 a_761_289.n2 354.616
R42 a_761_289.n1 a_761_289.t4 350.253
R43 a_761_289.n1 a_761_289.t5 189.586
R44 a_761_289.n2 a_761_289.n1 170.117
R45 a_761_289.n2 a_761_289.n0 167.836
R46 a_761_289.n3 a_761_289.t0 89.119
R47 a_761_289.n0 a_761_289.t1 63.333
R48 a_761_289.t3 a_761_289.n3 41.041
R49 a_761_289.n0 a_761_289.t2 31.979
R50 a_639_47.t0 a_639_47.t1 198.571
R51 a_805_47.t0 a_805_47.t1 60
R52 a_193_47.n0 a_193_47.t2 275.928
R53 a_193_47.n1 a_193_47.t5 258.716
R54 a_193_47.n1 a_193_47.t3 233.933
R55 a_193_47.n3 a_193_47.t0 232.798
R56 a_193_47.n0 a_193_47.t4 145.905
R57 a_193_47.t1 a_193_47.n3 123.515
R58 a_193_47.n2 a_193_47.n0 5.469
R59 a_193_47.n2 a_193_47.n1 4.65
R60 a_193_47.n3 a_193_47.n2 3.654
R61 a_1462_47.t0 a_1462_47.t1 87.142
R62 a_1283_21.n2 a_1283_21.n0 515.369
R63 a_1283_21.n3 a_1283_21.t4 389.181
R64 a_1283_21.n1 a_1283_21.t3 239.038
R65 a_1283_21.n4 a_1283_21.n3 175.164
R66 a_1283_21.n3 a_1283_21.t6 174.888
R67 a_1283_21.n1 a_1283_21.t5 166.738
R68 a_1283_21.t0 a_1283_21.n4 131.071
R69 a_1283_21.n2 a_1283_21.n1 88.16
R70 a_1283_21.n0 a_1283_21.t1 63.321
R71 a_1283_21.n0 a_1283_21.t2 63.321
R72 a_1283_21.n4 a_1283_21.n2 37.718
R73 a_543_47.n3 a_543_47.n2 381.836
R74 a_543_47.n1 a_543_47.t5 332.579
R75 a_543_47.n2 a_543_47.n0 191.51
R76 a_543_47.n2 a_543_47.n1 177.646
R77 a_543_47.n1 a_543_47.t4 168.699
R78 a_543_47.n3 a_543_47.t2 96.154
R79 a_543_47.t1 a_543_47.n3 65.666
R80 a_543_47.n0 a_543_47.t3 65
R81 a_543_47.n0 a_543_47.t0 45
R82 a_651_413.n0 a_651_413.t2 742.814
R83 a_651_413.n0 a_651_413.t1 194.654
R84 a_651_413.t0 a_651_413.n0 63.321
R85 VPB.t8 VPB.t3 790.186
R86 VPB.t7 VPB.t6 636.292
R87 VPB.t13 VPB.t4 583.021
R88 VPB.t10 VPB.t2 414.33
R89 VPB.t5 VPB.t12 319.626
R90 VPB.t4 VPB.t9 292.99
R91 VPB.t1 VPB.t10 292.99
R92 VPB.t2 VPB.t13 287.071
R93 VPB.t3 VPB.t1 272.274
R94 VPB.t9 VPB.t0 254.517
R95 VPB.t12 VPB.t7 248.598
R96 VPB.t0 VPB.t5 248.598
R97 VPB.t11 VPB.t8 248.598
R98 VPB VPB.t11 192.367
R99 RESET_B.n1 RESET_B.t3 413.312
R100 RESET_B.n4 RESET_B.t2 344.005
R101 RESET_B.n3 RESET_B.t1 187.32
R102 RESET_B.n1 RESET_B.t0 126.126
R103 RESET_B.n2 RESET_B.n1 13.102
R104 RESET_B.n5 RESET_B.n4 9.3
R105 RESET_B.n4 RESET_B.n3 9.159
R106 RESET_B.n2 RESET_B.n0 4.734
R107 RESET_B.n0 RESET_B 4.533
R108 RESET_B.n5 RESET_B.n2 3.214
R109 RESET_B RESET_B.n7 3.113
R110 RESET_B.n7 RESET_B.n6 1.556
R111 RESET_B.n6 RESET_B.n5 1.383
R112 VGND.n27 VGND.t7 215.034
R113 VGND.n0 VGND.t3 138.166
R114 VGND.n2 VGND.n1 116.752
R115 VGND.n12 VGND.n11 107.239
R116 VGND.n32 VGND.n31 107.239
R117 VGND.n1 VGND.t6 100
R118 VGND.n11 VGND.t5 72.857
R119 VGND.n1 VGND.t2 70
R120 VGND.n11 VGND.t1 60.579
R121 VGND.n31 VGND.t4 38.571
R122 VGND.n31 VGND.t0 38.571
R123 VGND.n4 VGND.n3 4.65
R124 VGND.n6 VGND.n5 4.65
R125 VGND.n8 VGND.n7 4.65
R126 VGND.n10 VGND.n9 4.65
R127 VGND.n14 VGND.n13 4.65
R128 VGND.n16 VGND.n15 4.65
R129 VGND.n18 VGND.n17 4.65
R130 VGND.n20 VGND.n19 4.65
R131 VGND.n22 VGND.n21 4.65
R132 VGND.n24 VGND.n23 4.65
R133 VGND.n26 VGND.n25 4.65
R134 VGND.n28 VGND.n27 4.65
R135 VGND.n30 VGND.n29 4.65
R136 VGND.n33 VGND.n32 3.932
R137 VGND.n3 VGND.n2 2.635
R138 VGND.n13 VGND.n12 1.882
R139 VGND.n4 VGND.n0 0.14
R140 VGND.n33 VGND.n30 0.137
R141 VGND VGND.n33 0.123
R142 VGND.n6 VGND.n4 0.119
R143 VGND.n8 VGND.n6 0.119
R144 VGND.n10 VGND.n8 0.119
R145 VGND.n14 VGND.n10 0.119
R146 VGND.n16 VGND.n14 0.119
R147 VGND.n18 VGND.n16 0.119
R148 VGND.n20 VGND.n18 0.119
R149 VGND.n22 VGND.n20 0.119
R150 VGND.n24 VGND.n22 0.119
R151 VGND.n26 VGND.n24 0.119
R152 VGND.n28 VGND.n26 0.119
R153 VGND.n30 VGND.n28 0.119
R154 VPWR.n13 VPWR.t2 514.01
R155 VPWR.n29 VPWR.t1 375.277
R156 VPWR.n0 VPWR.t5 375.25
R157 VPWR.n5 VPWR.n4 311.956
R158 VPWR.n36 VPWR.n35 311.893
R159 VPWR.n18 VPWR.n17 309.178
R160 VPWR.n1 VPWR.t4 200.298
R161 VPWR.n4 VPWR.t3 119.607
R162 VPWR.n17 VPWR.t0 93.809
R163 VPWR.n4 VPWR.t8 63.321
R164 VPWR.n17 VPWR.t9 63.321
R165 VPWR.n35 VPWR.t6 41.554
R166 VPWR.n35 VPWR.t7 41.554
R167 VPWR.n3 VPWR.n2 4.65
R168 VPWR.n6 VPWR.n5 4.65
R169 VPWR.n8 VPWR.n7 4.65
R170 VPWR.n10 VPWR.n9 4.65
R171 VPWR.n12 VPWR.n11 4.65
R172 VPWR.n14 VPWR.n13 4.65
R173 VPWR.n16 VPWR.n15 4.65
R174 VPWR.n20 VPWR.n19 4.65
R175 VPWR.n22 VPWR.n21 4.65
R176 VPWR.n24 VPWR.n23 4.65
R177 VPWR.n26 VPWR.n25 4.65
R178 VPWR.n28 VPWR.n27 4.65
R179 VPWR.n30 VPWR.n29 4.65
R180 VPWR.n32 VPWR.n31 4.65
R181 VPWR.n34 VPWR.n33 4.65
R182 VPWR.n1 VPWR.n0 4.195
R183 VPWR.n37 VPWR.n36 3.932
R184 VPWR.n19 VPWR.n18 3.764
R185 VPWR.n3 VPWR.n1 0.683
R186 VPWR.n37 VPWR.n34 0.137
R187 VPWR VPWR.n37 0.123
R188 VPWR.n6 VPWR.n3 0.119
R189 VPWR.n8 VPWR.n6 0.119
R190 VPWR.n10 VPWR.n8 0.119
R191 VPWR.n12 VPWR.n10 0.119
R192 VPWR.n14 VPWR.n12 0.119
R193 VPWR.n16 VPWR.n14 0.119
R194 VPWR.n20 VPWR.n16 0.119
R195 VPWR.n22 VPWR.n20 0.119
R196 VPWR.n24 VPWR.n22 0.119
R197 VPWR.n26 VPWR.n24 0.119
R198 VPWR.n28 VPWR.n26 0.119
R199 VPWR.n30 VPWR.n28 0.119
R200 VPWR.n32 VPWR.n30 0.119
R201 VPWR.n34 VPWR.n32 0.119
R202 Q.n1 Q.t0 207.309
R203 Q.n0 Q.t1 117.423
R204 Q Q.n0 47.901
R205 Q.n0 Q 10.29
R206 Q.n1 Q 9.192
R207 Q Q.n1 7.602
R208 CLK.n0 CLK.t0 294.554
R209 CLK.n0 CLK.t1 211.008
R210 CLK.n1 CLK.n0 76
R211 CLK.n1 CLK 10.422
R212 CLK CLK.n1 2.011
R213 D.n0 D.t1 333.651
R214 D.n0 D.t0 297.233
R215 D D.n0 120.734
R216 a_448_47.n1 a_448_47.n0 541.024
R217 a_448_47.t0 a_448_47.n1 82.083
R218 a_448_47.n0 a_448_47.t3 63.333
R219 a_448_47.n1 a_448_47.t1 63.321
R220 a_448_47.n0 a_448_47.t2 29.726
R221 a_1270_413.t0 a_1270_413.t1 126.642
C0 D VPWR 0.11fF
C1 VPB VPWR 0.19fF
C2 VPWR Q 0.13fF
C3 RESET_B VGND 0.37fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__dfrtp_2.ext - technology: sky130A

.subckt sky130_fd_sc_hd__dfrtp_2 Q RESET_B D CLK VGND VPWR VNB VPB
X0 a_1217_47.t0 a_27_47.t2 a_1108_47.t0 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X1 a_805_47.t0 a_761_289.t4 a_639_47.t1 VNB.t8 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 VGND.t1 a_1283_21.t3 Q.t1 VNB.t6 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 a_1108_47.t2 a_193_47.t2 a_761_289.t3 VNB.t11 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X4 a_1283_21.t0 a_1108_47.t4 a_1462_47.t0 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 a_651_413.t0 a_27_47.t3 a_543_47.t2 VPB.t8 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 VPWR.t1 a_1283_21.t4 Q.t3 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 VGND.t7 RESET_B.t0 a_805_47.t1 VNB.t13 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 Q.t2 a_1283_21.t5 VPWR.t0 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 VPWR.t3 CLK.t0 a_27_47.t0 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X10 a_448_47.t2 D.t0 VPWR.t10 VPB.t14 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11 a_761_289.t1 a_543_47.t4 VGND.t6 VNB.t9 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X12 a_193_47.t1 a_27_47.t4 VGND.t4 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13 a_1108_47.t1 a_27_47.t5 a_761_289.t0 VPB.t7 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14 a_543_47.t3 a_27_47.t6 a_448_47.t1 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X15 a_1462_47.t1 RESET_B.t1 VGND.t8 VNB.t14 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16 a_543_47.t0 a_193_47.t3 a_448_47.t0 VPB.t5 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17 a_448_47.t3 D.t1 VGND.t5 VNB.t5 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18 VPWR.t2 a_1283_21.t6 a_1270_413.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19 VPWR.t5 a_1108_47.t5 a_1283_21.t1 VPB.t9 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20 a_1270_413.t1 a_193_47.t4 a_1108_47.t3 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21 a_193_47.t0 a_27_47.t7 VPWR.t4 VPB.t6 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X22 a_1283_21.t2 RESET_B.t2 VPWR.t8 VPB.t12 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23 VPWR.t7 a_761_289.t5 a_651_413.t1 VPB.t11 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24 Q.t0 a_1283_21.t7 VGND.t0 VNB.t7 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X25 a_639_47.t0 a_193_47.t5 a_543_47.t1 VNB.t12 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X26 VGND.t2 a_1283_21.t8 a_1217_47.t1 VNB.t10 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X27 a_651_413.t2 RESET_B.t3 VPWR.t9 VPB.t13 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X28 VGND.t3 CLK.t1 a_27_47.t1 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X29 a_761_289.t2 a_543_47.t5 VPWR.t6 VPB.t10 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
R0 a_27_47.n1 a_27_47.t3 530.008
R1 a_27_47.n0 a_27_47.t5 331.026
R2 a_27_47.t0 a_27_47.n9 271.418
R3 a_27_47.n4 a_27_47.t7 255.459
R4 a_27_47.n6 a_27_47.t4 224.611
R5 a_27_47.n0 a_27_47.t2 204.373
R6 a_27_47.n3 a_27_47.t1 186.535
R7 a_27_47.n1 a_27_47.t6 141.921
R8 a_27_47.n2 a_27_47.n1 90.158
R9 a_27_47.n2 a_27_47.n0 12.643
R10 a_27_47.n7 a_27_47.n6 8.764
R11 a_27_47.n5 a_27_47.n4 7.712
R12 a_27_47.n9 a_27_47.n8 3.339
R13 a_27_47.n6 a_27_47.n5 3.213
R14 a_27_47.n3 a_27_47.n2 3.151
R15 a_27_47.n8 a_27_47.n7 1.391
R16 a_27_47.n7 a_27_47.n3 1.094
R17 a_1108_47.n1 a_1108_47.t4 366.855
R18 a_1108_47.n3 a_1108_47.n2 344.452
R19 a_1108_47.n2 a_1108_47.n0 207.699
R20 a_1108_47.n1 a_1108_47.t5 174.055
R21 a_1108_47.n2 a_1108_47.n1 149.035
R22 a_1108_47.n0 a_1108_47.t2 70
R23 a_1108_47.t1 a_1108_47.n3 68.011
R24 a_1108_47.n3 a_1108_47.t3 63.321
R25 a_1108_47.n0 a_1108_47.t0 61.666
R26 a_1217_47.t1 a_1217_47.t0 94.726
R27 VNB.t2 VNB.t5 8250
R28 VNB VNB.t0 6470.59
R29 VNB.t4 VNB.t7 5985.29
R30 VNB.t12 VNB.t8 5370.59
R31 VNB.t10 VNB.t14 4820.59
R32 VNB.t13 VNB.t9 3550.91
R33 VNB.t11 VNB.t3 3526.47
R34 VNB.t3 VNB.t10 3105.88
R35 VNB.t1 VNB.t12 3105.88
R36 VNB.t5 VNB.t1 3073.53
R37 VNB.t14 VNB.t4 2944.12
R38 VNB.t0 VNB.t2 2717.65
R39 VNB.t9 VNB.t11 2377.92
R40 VNB.t8 VNB.t13 2329.41
R41 VNB.t7 VNB.t6 2030.77
R42 a_761_289.n3 a_761_289.n2 354.616
R43 a_761_289.n1 a_761_289.t4 350.253
R44 a_761_289.n1 a_761_289.t5 189.586
R45 a_761_289.n2 a_761_289.n1 170.117
R46 a_761_289.n2 a_761_289.n0 167.836
R47 a_761_289.n3 a_761_289.t0 89.119
R48 a_761_289.n0 a_761_289.t3 63.333
R49 a_761_289.t2 a_761_289.n3 41.041
R50 a_761_289.n0 a_761_289.t1 31.979
R51 a_639_47.t1 a_639_47.t0 198.571
R52 a_805_47.t0 a_805_47.t1 60
R53 a_1283_21.n3 a_1283_21.n0 515.369
R54 a_1283_21.n4 a_1283_21.t6 389.181
R55 a_1283_21.n1 a_1283_21.t4 212.079
R56 a_1283_21.n2 a_1283_21.t5 212.079
R57 a_1283_21.n5 a_1283_21.n4 175.164
R58 a_1283_21.n4 a_1283_21.t8 174.888
R59 a_1283_21.n1 a_1283_21.t3 139.779
R60 a_1283_21.n2 a_1283_21.t7 139.779
R61 a_1283_21.t0 a_1283_21.n5 131.071
R62 a_1283_21.n3 a_1283_21.n2 100.575
R63 a_1283_21.n0 a_1283_21.t1 63.321
R64 a_1283_21.n0 a_1283_21.t2 63.321
R65 a_1283_21.n2 a_1283_21.n1 61.345
R66 a_1283_21.n5 a_1283_21.n3 37.718
R67 Q.n3 Q.n2 142.894
R68 Q.n1 Q.n0 92.5
R69 Q Q.n1 49.033
R70 Q.n2 Q.t3 26.595
R71 Q.n2 Q.t2 26.595
R72 Q.n0 Q.t1 24.923
R73 Q.n0 Q.t0 24.923
R74 Q.n1 Q 10.496
R75 Q.n3 Q 9.375
R76 Q Q.n3 7.629
R77 VGND.n34 VGND.t5 215.034
R78 VGND.n1 VGND.t1 149.626
R79 VGND.n0 VGND.t0 134.381
R80 VGND.n9 VGND.n8 116.752
R81 VGND.n19 VGND.n18 107.239
R82 VGND.n39 VGND.n38 107.239
R83 VGND.n8 VGND.t8 100
R84 VGND.n18 VGND.t7 72.857
R85 VGND.n8 VGND.t2 70
R86 VGND.n18 VGND.t6 60.579
R87 VGND.n38 VGND.t4 38.571
R88 VGND.n38 VGND.t3 38.571
R89 VGND.n3 VGND.n2 4.65
R90 VGND.n5 VGND.n4 4.65
R91 VGND.n7 VGND.n6 4.65
R92 VGND.n11 VGND.n10 4.65
R93 VGND.n13 VGND.n12 4.65
R94 VGND.n15 VGND.n14 4.65
R95 VGND.n17 VGND.n16 4.65
R96 VGND.n21 VGND.n20 4.65
R97 VGND.n23 VGND.n22 4.65
R98 VGND.n25 VGND.n24 4.65
R99 VGND.n27 VGND.n26 4.65
R100 VGND.n29 VGND.n28 4.65
R101 VGND.n31 VGND.n30 4.65
R102 VGND.n33 VGND.n32 4.65
R103 VGND.n35 VGND.n34 4.65
R104 VGND.n37 VGND.n36 4.65
R105 VGND.n40 VGND.n39 3.932
R106 VGND.n1 VGND.n0 3.811
R107 VGND.n10 VGND.n9 2.635
R108 VGND.n20 VGND.n19 1.882
R109 VGND.n3 VGND.n1 0.243
R110 VGND.n40 VGND.n37 0.137
R111 VGND VGND.n40 0.123
R112 VGND.n5 VGND.n3 0.119
R113 VGND.n7 VGND.n5 0.119
R114 VGND.n11 VGND.n7 0.119
R115 VGND.n13 VGND.n11 0.119
R116 VGND.n15 VGND.n13 0.119
R117 VGND.n17 VGND.n15 0.119
R118 VGND.n21 VGND.n17 0.119
R119 VGND.n23 VGND.n21 0.119
R120 VGND.n25 VGND.n23 0.119
R121 VGND.n27 VGND.n25 0.119
R122 VGND.n29 VGND.n27 0.119
R123 VGND.n31 VGND.n29 0.119
R124 VGND.n33 VGND.n31 0.119
R125 VGND.n35 VGND.n33 0.119
R126 VGND.n37 VGND.n35 0.119
R127 a_193_47.n0 a_193_47.t2 275.928
R128 a_193_47.n1 a_193_47.t5 258.716
R129 a_193_47.n1 a_193_47.t3 233.933
R130 a_193_47.n3 a_193_47.t1 232.798
R131 a_193_47.n0 a_193_47.t4 145.905
R132 a_193_47.t0 a_193_47.n3 123.515
R133 a_193_47.n2 a_193_47.n0 5.469
R134 a_193_47.n2 a_193_47.n1 4.65
R135 a_193_47.n3 a_193_47.n2 3.654
R136 a_1462_47.t0 a_1462_47.t1 87.142
R137 a_543_47.n3 a_543_47.n2 381.836
R138 a_543_47.n1 a_543_47.t5 332.579
R139 a_543_47.n2 a_543_47.n0 191.51
R140 a_543_47.n2 a_543_47.n1 177.646
R141 a_543_47.n1 a_543_47.t4 168.699
R142 a_543_47.n3 a_543_47.t2 96.154
R143 a_543_47.t0 a_543_47.n3 65.666
R144 a_543_47.n0 a_543_47.t3 65
R145 a_543_47.n0 a_543_47.t1 45
R146 a_651_413.n0 a_651_413.t2 742.814
R147 a_651_413.t0 a_651_413.n0 194.654
R148 a_651_413.n0 a_651_413.t1 63.321
R149 VPB.t6 VPB.t14 790.186
R150 VPB.t9 VPB.t1 636.292
R151 VPB.t13 VPB.t10 583.021
R152 VPB.t8 VPB.t11 414.33
R153 VPB.t0 VPB.t12 319.626
R154 VPB.t10 VPB.t7 292.99
R155 VPB.t5 VPB.t8 292.99
R156 VPB.t11 VPB.t13 287.071
R157 VPB.t14 VPB.t5 272.274
R158 VPB.t7 VPB.t4 254.517
R159 VPB.t1 VPB.t2 248.598
R160 VPB.t12 VPB.t9 248.598
R161 VPB.t4 VPB.t0 248.598
R162 VPB.t3 VPB.t6 248.598
R163 VPB VPB.t3 192.367
R164 VPWR.n16 VPWR.t6 514.01
R165 VPWR.n32 VPWR.t10 375.277
R166 VPWR.n2 VPWR.t5 375.25
R167 VPWR.n8 VPWR.n7 311.956
R168 VPWR.n39 VPWR.n38 311.893
R169 VPWR.n21 VPWR.n20 309.178
R170 VPWR.n0 VPWR.t0 197.285
R171 VPWR.n1 VPWR.t1 156.759
R172 VPWR.n7 VPWR.t2 119.607
R173 VPWR.n20 VPWR.t7 93.809
R174 VPWR.n7 VPWR.t8 63.321
R175 VPWR.n20 VPWR.t9 63.321
R176 VPWR.n38 VPWR.t4 41.554
R177 VPWR.n38 VPWR.t3 41.554
R178 VPWR.n4 VPWR.n3 4.65
R179 VPWR.n6 VPWR.n5 4.65
R180 VPWR.n9 VPWR.n8 4.65
R181 VPWR.n11 VPWR.n10 4.65
R182 VPWR.n13 VPWR.n12 4.65
R183 VPWR.n15 VPWR.n14 4.65
R184 VPWR.n17 VPWR.n16 4.65
R185 VPWR.n19 VPWR.n18 4.65
R186 VPWR.n23 VPWR.n22 4.65
R187 VPWR.n25 VPWR.n24 4.65
R188 VPWR.n27 VPWR.n26 4.65
R189 VPWR.n29 VPWR.n28 4.65
R190 VPWR.n31 VPWR.n30 4.65
R191 VPWR.n33 VPWR.n32 4.65
R192 VPWR.n35 VPWR.n34 4.65
R193 VPWR.n37 VPWR.n36 4.65
R194 VPWR.n40 VPWR.n39 3.932
R195 VPWR.n1 VPWR.n0 3.811
R196 VPWR.n22 VPWR.n21 3.764
R197 VPWR.n3 VPWR.n2 0.752
R198 VPWR.n4 VPWR.n1 0.243
R199 VPWR.n40 VPWR.n37 0.137
R200 VPWR VPWR.n40 0.123
R201 VPWR.n6 VPWR.n4 0.119
R202 VPWR.n9 VPWR.n6 0.119
R203 VPWR.n11 VPWR.n9 0.119
R204 VPWR.n13 VPWR.n11 0.119
R205 VPWR.n15 VPWR.n13 0.119
R206 VPWR.n17 VPWR.n15 0.119
R207 VPWR.n19 VPWR.n17 0.119
R208 VPWR.n23 VPWR.n19 0.119
R209 VPWR.n25 VPWR.n23 0.119
R210 VPWR.n27 VPWR.n25 0.119
R211 VPWR.n29 VPWR.n27 0.119
R212 VPWR.n31 VPWR.n29 0.119
R213 VPWR.n33 VPWR.n31 0.119
R214 VPWR.n35 VPWR.n33 0.119
R215 VPWR.n37 VPWR.n35 0.119
R216 RESET_B.n1 RESET_B.t3 413.312
R217 RESET_B.n4 RESET_B.t2 344.005
R218 RESET_B.n3 RESET_B.t1 187.32
R219 RESET_B.n1 RESET_B.t0 126.126
R220 RESET_B.n2 RESET_B.n1 13.102
R221 RESET_B.n5 RESET_B.n4 9.3
R222 RESET_B.n4 RESET_B.n3 9.159
R223 RESET_B.n2 RESET_B.n0 4.734
R224 RESET_B.n0 RESET_B 4.533
R225 RESET_B.n5 RESET_B.n2 3.214
R226 RESET_B RESET_B.n7 3.113
R227 RESET_B.n7 RESET_B.n6 1.556
R228 RESET_B.n6 RESET_B.n5 1.383
R229 CLK.n0 CLK.t0 294.554
R230 CLK.n0 CLK.t1 211.008
R231 CLK.n1 CLK.n0 76
R232 CLK.n1 CLK 10.422
R233 CLK CLK.n1 2.011
R234 D.n0 D.t1 333.651
R235 D.n0 D.t0 297.233
R236 D D.n0 120.734
R237 a_448_47.n1 a_448_47.n0 541.024
R238 a_448_47.t0 a_448_47.n1 82.083
R239 a_448_47.n0 a_448_47.t1 63.333
R240 a_448_47.n1 a_448_47.t2 63.321
R241 a_448_47.n0 a_448_47.t3 29.726
R242 a_1270_413.t0 a_1270_413.t1 126.642
C0 VGND Q 0.15fF
C1 VPWR Q 0.27fF
C2 VPWR VGND 0.11fF
C3 RESET_B VGND 0.37fF
C4 D VPWR 0.11fF
C5 VPB VPWR 0.20fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__dfrtp_4.ext - technology: sky130A

.subckt sky130_fd_sc_hd__dfrtp_4 Q RESET_B D CLK VGND VPWR VNB VPB
X0 a_1217_47.t0 a_27_47.t2 a_1108_47.t1 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X1 a_805_47.t0 a_761_289.t4 a_639_47.t1 VNB.t16 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 a_1108_47.t2 a_193_47.t2 a_761_289.t1 VNB.t11 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X3 a_1283_21.t0 a_1108_47.t4 a_1462_47.t0 VNB.t10 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 a_651_413.t0 a_27_47.t3 a_543_47.t1 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 VGND.t8 RESET_B.t0 a_805_47.t1 VNB.t13 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 VPWR.t5 a_1283_21.t3 Q.t7 VPB.t7 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 VPWR.t12 CLK.t0 a_27_47.t0 VPB.t15 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X8 a_448_47.t2 D.t0 VPWR.t7 VPB.t11 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9 Q.t6 a_1283_21.t4 VPWR.t4 VPB.t6 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 VPWR.t3 a_1283_21.t5 Q.t5 VPB.t5 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 a_761_289.t2 a_543_47.t4 VGND.t6 VNB.t12 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X12 Q.t3 a_1283_21.t6 VGND.t5 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 a_193_47.t0 a_27_47.t4 VGND.t0 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14 a_1108_47.t0 a_27_47.t5 a_761_289.t0 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15 a_543_47.t0 a_27_47.t6 a_448_47.t0 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X16 a_1462_47.t1 RESET_B.t1 VGND.t9 VNB.t14 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17 a_543_47.t3 a_193_47.t3 a_448_47.t3 VPB.t10 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18 a_448_47.t1 D.t1 VGND.t7 VNB.t8 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19 VPWR.t1 a_1283_21.t7 a_1270_413.t0 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20 VPWR.t8 a_1108_47.t5 a_1283_21.t1 VPB.t12 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21 Q.t4 a_1283_21.t8 VPWR.t2 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X22 a_1270_413.t1 a_193_47.t4 a_1108_47.t3 VPB.t9 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23 a_193_47.t1 a_27_47.t7 VPWR.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X24 a_1283_21.t2 RESET_B.t2 VPWR.t9 VPB.t14 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X25 VGND.t4 a_1283_21.t9 Q.t2 VNB.t5 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X26 VGND.t3 a_1283_21.t10 Q.t1 VNB.t6 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X27 VPWR.t11 a_761_289.t5 a_651_413.t1 VPB.t13 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X28 a_639_47.t0 a_193_47.t5 a_543_47.t2 VNB.t9 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X29 VGND.t1 a_1283_21.t11 a_1217_47.t1 VNB.t7 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X30 a_651_413.t2 RESET_B.t3 VPWR.t10 VPB.t16 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X31 VGND.t10 CLK.t1 a_27_47.t1 VNB.t15 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X32 a_761_289.t3 a_543_47.t5 VPWR.t6 VPB.t8 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X33 Q.t0 a_1283_21.t12 VGND.t2 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
R0 a_27_47.n1 a_27_47.t3 530.008
R1 a_27_47.n0 a_27_47.t5 331.026
R2 a_27_47.t0 a_27_47.n9 271.418
R3 a_27_47.n4 a_27_47.t7 255.459
R4 a_27_47.n6 a_27_47.t4 224.611
R5 a_27_47.n0 a_27_47.t2 204.373
R6 a_27_47.n3 a_27_47.t1 186.535
R7 a_27_47.n1 a_27_47.t6 141.921
R8 a_27_47.n2 a_27_47.n1 90.158
R9 a_27_47.n2 a_27_47.n0 12.643
R10 a_27_47.n7 a_27_47.n6 8.764
R11 a_27_47.n5 a_27_47.n4 7.712
R12 a_27_47.n9 a_27_47.n8 3.339
R13 a_27_47.n6 a_27_47.n5 3.213
R14 a_27_47.n3 a_27_47.n2 3.151
R15 a_27_47.n8 a_27_47.n7 1.391
R16 a_27_47.n7 a_27_47.n3 1.094
R17 a_1108_47.n1 a_1108_47.t4 366.855
R18 a_1108_47.n3 a_1108_47.n2 344.452
R19 a_1108_47.n2 a_1108_47.n0 207.699
R20 a_1108_47.n1 a_1108_47.t5 174.055
R21 a_1108_47.n2 a_1108_47.n1 149.035
R22 a_1108_47.n0 a_1108_47.t2 70
R23 a_1108_47.t0 a_1108_47.n3 68.011
R24 a_1108_47.n3 a_1108_47.t3 63.321
R25 a_1108_47.n0 a_1108_47.t1 61.666
R26 a_1217_47.t1 a_1217_47.t0 94.726
R27 VNB.t1 VNB.t8 8250
R28 VNB VNB.t15 6470.59
R29 VNB.t9 VNB.t16 5370.59
R30 VNB.t10 VNB.t4 5321.88
R31 VNB.t7 VNB.t14 4820.59
R32 VNB.t13 VNB.t12 3550.91
R33 VNB.t11 VNB.t2 3526.47
R34 VNB.t2 VNB.t7 3105.88
R35 VNB.t0 VNB.t9 3105.88
R36 VNB.t8 VNB.t0 3073.53
R37 VNB.t14 VNB.t10 2944.12
R38 VNB.t15 VNB.t1 2717.65
R39 VNB.t12 VNB.t11 2377.92
R40 VNB.t16 VNB.t13 2329.41
R41 VNB.t3 VNB.t6 2030.77
R42 VNB.t5 VNB.t3 2030.77
R43 VNB.t4 VNB.t5 2030.77
R44 a_761_289.n3 a_761_289.n2 354.616
R45 a_761_289.n1 a_761_289.t4 350.253
R46 a_761_289.n1 a_761_289.t5 189.586
R47 a_761_289.n2 a_761_289.n1 170.117
R48 a_761_289.n2 a_761_289.n0 167.836
R49 a_761_289.n3 a_761_289.t0 89.119
R50 a_761_289.n0 a_761_289.t1 63.333
R51 a_761_289.t3 a_761_289.n3 41.041
R52 a_761_289.n0 a_761_289.t2 31.979
R53 a_639_47.t1 a_639_47.t0 198.571
R54 a_805_47.t0 a_805_47.t1 60
R55 a_193_47.n0 a_193_47.t2 275.928
R56 a_193_47.n1 a_193_47.t5 258.716
R57 a_193_47.n1 a_193_47.t3 233.933
R58 a_193_47.n3 a_193_47.t0 232.798
R59 a_193_47.n0 a_193_47.t4 145.905
R60 a_193_47.t1 a_193_47.n3 123.515
R61 a_193_47.n2 a_193_47.n0 5.469
R62 a_193_47.n2 a_193_47.n1 4.65
R63 a_193_47.n3 a_193_47.n2 3.654
R64 a_1462_47.t0 a_1462_47.t1 87.142
R65 a_1283_21.n12 a_1283_21.n11 400.294
R66 a_1283_21.n13 a_1283_21.t7 389.181
R67 a_1283_21.n0 a_1283_21.t3 212.079
R68 a_1283_21.n2 a_1283_21.t4 212.079
R69 a_1283_21.n5 a_1283_21.t5 212.079
R70 a_1283_21.n8 a_1283_21.t8 212.079
R71 a_1283_21.n14 a_1283_21.n13 175.164
R72 a_1283_21.n13 a_1283_21.t11 174.888
R73 a_1283_21.n0 a_1283_21.t10 139.779
R74 a_1283_21.n2 a_1283_21.t12 139.779
R75 a_1283_21.n5 a_1283_21.t9 139.779
R76 a_1283_21.n8 a_1283_21.t6 139.779
R77 a_1283_21.t0 a_1283_21.n14 131.071
R78 a_1283_21.n4 a_1283_21.n1 96.723
R79 a_1283_21.n10 a_1283_21.n9 76
R80 a_1283_21.n4 a_1283_21.n3 76
R81 a_1283_21.n7 a_1283_21.n6 76
R82 a_1283_21.n11 a_1283_21.t1 63.321
R83 a_1283_21.n11 a_1283_21.t2 63.321
R84 a_1283_21.n1 a_1283_21.n0 30.672
R85 a_1283_21.n12 a_1283_21.n10 30.476
R86 a_1283_21.n14 a_1283_21.n12 28.338
R87 a_1283_21.n7 a_1283_21.n4 20.723
R88 a_1283_21.n10 a_1283_21.n7 20.723
R89 a_1283_21.n3 a_1283_21.n2 18.987
R90 a_1283_21.n6 a_1283_21.n5 7.303
R91 a_1283_21.n9 a_1283_21.n8 4.381
R92 a_543_47.n3 a_543_47.n2 381.836
R93 a_543_47.n1 a_543_47.t5 332.579
R94 a_543_47.n2 a_543_47.n0 191.51
R95 a_543_47.n2 a_543_47.n1 177.646
R96 a_543_47.n1 a_543_47.t4 168.699
R97 a_543_47.t1 a_543_47.n3 96.154
R98 a_543_47.n3 a_543_47.t3 65.666
R99 a_543_47.n0 a_543_47.t0 65
R100 a_543_47.n0 a_543_47.t2 45
R101 a_651_413.n0 a_651_413.t2 742.814
R102 a_651_413.t0 a_651_413.n0 194.654
R103 a_651_413.n0 a_651_413.t1 63.321
R104 VPB.t0 VPB.t11 790.186
R105 VPB.t16 VPB.t8 583.021
R106 VPB.t12 VPB.t3 577.102
R107 VPB.t2 VPB.t13 414.33
R108 VPB.t4 VPB.t14 319.626
R109 VPB.t8 VPB.t1 292.99
R110 VPB.t10 VPB.t2 292.99
R111 VPB.t13 VPB.t16 287.071
R112 VPB.t11 VPB.t10 272.274
R113 VPB.t1 VPB.t9 254.517
R114 VPB.t6 VPB.t7 248.598
R115 VPB.t5 VPB.t6 248.598
R116 VPB.t3 VPB.t5 248.598
R117 VPB.t14 VPB.t12 248.598
R118 VPB.t9 VPB.t4 248.598
R119 VPB.t15 VPB.t0 248.598
R120 VPB VPB.t15 192.367
R121 RESET_B.n1 RESET_B.t3 413.312
R122 RESET_B.n4 RESET_B.t2 344.005
R123 RESET_B.n3 RESET_B.t1 187.32
R124 RESET_B.n1 RESET_B.t0 126.126
R125 RESET_B.n2 RESET_B.n1 13.102
R126 RESET_B.n5 RESET_B.n4 9.3
R127 RESET_B.n4 RESET_B.n3 9.159
R128 RESET_B.n2 RESET_B.n0 4.734
R129 RESET_B.n0 RESET_B 4.533
R130 RESET_B.n5 RESET_B.n2 3.214
R131 RESET_B RESET_B.n7 3.113
R132 RESET_B.n7 RESET_B.n6 1.556
R133 RESET_B.n6 RESET_B.n5 1.383
R134 VGND.n40 VGND.t7 215.034
R135 VGND.n2 VGND.t3 198.965
R136 VGND.n15 VGND.n14 116.752
R137 VGND.n1 VGND.n0 115.464
R138 VGND.n5 VGND.t5 114.4
R139 VGND.n25 VGND.n24 107.239
R140 VGND.n45 VGND.n44 107.239
R141 VGND.n14 VGND.t9 100
R142 VGND.n24 VGND.t8 72.857
R143 VGND.n14 VGND.t1 70
R144 VGND.n24 VGND.t6 60.579
R145 VGND.n44 VGND.t0 38.571
R146 VGND.n44 VGND.t10 38.571
R147 VGND.n0 VGND.t2 24.923
R148 VGND.n0 VGND.t4 24.923
R149 VGND.n2 VGND.n1 16.676
R150 VGND.n6 VGND.n5 6.776
R151 VGND.n4 VGND.n3 4.65
R152 VGND.n7 VGND.n6 4.65
R153 VGND.n9 VGND.n8 4.65
R154 VGND.n11 VGND.n10 4.65
R155 VGND.n13 VGND.n12 4.65
R156 VGND.n17 VGND.n16 4.65
R157 VGND.n19 VGND.n18 4.65
R158 VGND.n21 VGND.n20 4.65
R159 VGND.n23 VGND.n22 4.65
R160 VGND.n27 VGND.n26 4.65
R161 VGND.n29 VGND.n28 4.65
R162 VGND.n31 VGND.n30 4.65
R163 VGND.n33 VGND.n32 4.65
R164 VGND.n35 VGND.n34 4.65
R165 VGND.n37 VGND.n36 4.65
R166 VGND.n39 VGND.n38 4.65
R167 VGND.n41 VGND.n40 4.65
R168 VGND.n43 VGND.n42 4.65
R169 VGND.n46 VGND.n45 3.932
R170 VGND.n16 VGND.n15 2.635
R171 VGND.n26 VGND.n25 1.882
R172 VGND.n4 VGND.n2 0.398
R173 VGND.n46 VGND.n43 0.137
R174 VGND VGND.n46 0.123
R175 VGND.n7 VGND.n4 0.119
R176 VGND.n9 VGND.n7 0.119
R177 VGND.n11 VGND.n9 0.119
R178 VGND.n13 VGND.n11 0.119
R179 VGND.n17 VGND.n13 0.119
R180 VGND.n19 VGND.n17 0.119
R181 VGND.n21 VGND.n19 0.119
R182 VGND.n23 VGND.n21 0.119
R183 VGND.n27 VGND.n23 0.119
R184 VGND.n29 VGND.n27 0.119
R185 VGND.n31 VGND.n29 0.119
R186 VGND.n33 VGND.n31 0.119
R187 VGND.n35 VGND.n33 0.119
R188 VGND.n37 VGND.n35 0.119
R189 VGND.n39 VGND.n37 0.119
R190 VGND.n41 VGND.n39 0.119
R191 VGND.n43 VGND.n41 0.119
R192 Q.n2 Q.n0 150.4
R193 Q.n2 Q.n1 110.76
R194 Q.n5 Q.n3 91.218
R195 Q.n5 Q.n4 52.818
R196 Q.n0 Q.t5 26.595
R197 Q.n0 Q.t4 26.595
R198 Q.n1 Q.t7 26.595
R199 Q.n1 Q.t6 26.595
R200 Q.n3 Q.t2 24.923
R201 Q.n3 Q.t3 24.923
R202 Q.n4 Q.t1 24.923
R203 Q.n4 Q.t0 24.923
R204 Q Q.n2 19.906
R205 Q.n6 Q.n5 13.929
R206 Q Q.n6 8.897
R207 Q.n6  1.717
R208 VPWR.n22 VPWR.t6 514.01
R209 VPWR.n38 VPWR.t7 375.277
R210 VPWR.n8 VPWR.t8 375.25
R211 VPWR.n14 VPWR.n13 311.956
R212 VPWR.n45 VPWR.n44 311.893
R213 VPWR.n27 VPWR.n26 309.178
R214 VPWR.n2 VPWR.t5 214.845
R215 VPWR.n5 VPWR.t2 201.189
R216 VPWR.n1 VPWR.n0 177.606
R217 VPWR.n13 VPWR.t1 119.607
R218 VPWR.n26 VPWR.t11 93.809
R219 VPWR.n13 VPWR.t9 63.321
R220 VPWR.n26 VPWR.t10 63.321
R221 VPWR.n44 VPWR.t0 41.554
R222 VPWR.n44 VPWR.t12 41.554
R223 VPWR.n0 VPWR.t4 26.595
R224 VPWR.n0 VPWR.t3 26.595
R225 VPWR.n2 VPWR.n1 16.676
R226 VPWR.n6 VPWR.n5 6.776
R227 VPWR.n4 VPWR.n3 4.65
R228 VPWR.n7 VPWR.n6 4.65
R229 VPWR.n10 VPWR.n9 4.65
R230 VPWR.n12 VPWR.n11 4.65
R231 VPWR.n15 VPWR.n14 4.65
R232 VPWR.n17 VPWR.n16 4.65
R233 VPWR.n19 VPWR.n18 4.65
R234 VPWR.n21 VPWR.n20 4.65
R235 VPWR.n23 VPWR.n22 4.65
R236 VPWR.n25 VPWR.n24 4.65
R237 VPWR.n29 VPWR.n28 4.65
R238 VPWR.n31 VPWR.n30 4.65
R239 VPWR.n33 VPWR.n32 4.65
R240 VPWR.n35 VPWR.n34 4.65
R241 VPWR.n37 VPWR.n36 4.65
R242 VPWR.n39 VPWR.n38 4.65
R243 VPWR.n41 VPWR.n40 4.65
R244 VPWR.n43 VPWR.n42 4.65
R245 VPWR.n46 VPWR.n45 3.932
R246 VPWR.n28 VPWR.n27 3.764
R247 VPWR.n9 VPWR.n8 0.752
R248 VPWR.n4 VPWR.n2 0.398
R249 VPWR.n46 VPWR.n43 0.137
R250 VPWR VPWR.n46 0.123
R251 VPWR.n7 VPWR.n4 0.119
R252 VPWR.n10 VPWR.n7 0.119
R253 VPWR.n12 VPWR.n10 0.119
R254 VPWR.n15 VPWR.n12 0.119
R255 VPWR.n17 VPWR.n15 0.119
R256 VPWR.n19 VPWR.n17 0.119
R257 VPWR.n21 VPWR.n19 0.119
R258 VPWR.n23 VPWR.n21 0.119
R259 VPWR.n25 VPWR.n23 0.119
R260 VPWR.n29 VPWR.n25 0.119
R261 VPWR.n31 VPWR.n29 0.119
R262 VPWR.n33 VPWR.n31 0.119
R263 VPWR.n35 VPWR.n33 0.119
R264 VPWR.n37 VPWR.n35 0.119
R265 VPWR.n39 VPWR.n37 0.119
R266 VPWR.n41 VPWR.n39 0.119
R267 VPWR.n43 VPWR.n41 0.119
R268 CLK.n0 CLK.t0 294.554
R269 CLK.n0 CLK.t1 211.008
R270 CLK.n1 CLK.n0 76
R271 CLK.n1 CLK 10.422
R272 CLK CLK.n1 2.011
R273 D.n0 D.t1 333.651
R274 D.n0 D.t0 297.233
R275 D D.n0 120.734
R276 a_448_47.n1 a_448_47.n0 541.024
R277 a_448_47.n0 a_448_47.t3 82.083
R278 a_448_47.n1 a_448_47.t0 63.333
R279 a_448_47.n0 a_448_47.t2 63.321
R280 a_448_47.n2 a_448_47.t1 26.393
R281 a_448_47.n3 a_448_47.n2 14.4
R282 a_448_47.n2 a_448_47.n1 3.333
R283 a_1270_413.t0 a_1270_413.t1 126.642
C0 VPWR VPB 0.22fF
C1 VPWR VGND 0.12fF
C2 RESET_B VGND 0.37fF
C3 D VPWR 0.11fF
C4 Q VGND 0.49fF
C5 Q VPWR 0.60fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__dfsbp_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__dfsbp_1 Q Q_N D VPWR SET_B CLK VGND VNB VPB
X0 a_1178_261.t1 a_1028_413.t5 VPWR.t1 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X1 VGND.t8 a_652_21.t3 a_586_47.t0 VNB.t10 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 a_1178_261.t0 a_1028_413.t6 VGND.t2 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=540000u l=150000u
X3 a_956_413.t0 a_476_47.t4 VPWR.t10 VPB.t12 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 a_1136_413.t0 a_193_47.t2 a_1028_413.t3 VPB.t14 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 VPWR.t11 a_476_47.t5 a_652_21.t1 VPB.t13 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 a_586_47.t1 a_193_47.t3 a_476_47.t2 VNB.t14 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X7 VPWR.t0 CLK.t0 a_27_47.t1 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X8 a_476_47.t0 a_27_47.t2 a_381_47.t3 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X9 a_1056_47.t0 a_476_47.t6 VGND.t9 VNB.t12 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10 Q.t0 a_1786_47.t2 VGND.t10 VNB.t16 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 a_381_47.t1 D.t0 VPWR.t7 VPB.t8 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X12 a_652_21.t0 SET_B.t0 VPWR.t8 VPB.t9 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13 a_1224_47.t1 a_27_47.t3 a_1028_413.t0 VNB.t5 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14 VGND.t3 a_1028_413.t7 a_1786_47.t0 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15 a_562_413.t1 a_27_47.t4 a_476_47.t1 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16 VPWR.t3 a_1028_413.t8 a_1786_47.t1 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X17 a_1028_413.t4 a_193_47.t4 a_1056_47.t1 VNB.t15 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18 a_476_47.t3 a_193_47.t5 a_381_47.t0 VPB.t15 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19 a_1296_47.t0 a_1178_261.t2 a_1224_47.t0 VNB.t11 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20 Q_N.t0 a_1028_413.t9 VGND.t1 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X21 a_193_47.t0 a_27_47.t5 VGND.t4 VNB.t6 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22 VPWR.t6 a_652_21.t4 a_562_413.t0 VPB.t7 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23 VGND.t6 SET_B.t1 a_1296_47.t1 VNB.t8 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24 a_1028_413.t1 a_27_47.t6 a_956_413.t1 VPB.t5 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X25 VPWR.t5 a_1178_261.t3 a_1136_413.t1 VPB.t11 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X26 a_193_47.t1 a_27_47.t7 VPWR.t4 VPB.t6 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X27 Q_N.t1 a_1028_413.t10 VPWR.t2 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X28 a_796_47.t1 SET_B.t2 VGND.t7 VNB.t9 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X29 a_381_47.t2 D.t1 VGND.t5 VNB.t7 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X30 Q.t1 a_1786_47.t3 VPWR.t12 VPB.t16 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X31 a_652_21.t2 a_476_47.t7 a_796_47.t0 VNB.t13 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X32 VPWR.t9 SET_B.t3 a_1028_413.t2 VPB.t10 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X33 VGND.t0 CLK.t1 a_27_47.t0 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
R0 a_1028_413.n5 a_1028_413.t2 432.15
R1 a_1028_413.n5 a_1028_413.n4 319.003
R2 a_1028_413.n3 a_1028_413.t5 258.673
R3 a_1028_413.n0 a_1028_413.t8 257.18
R4 a_1028_413.n1 a_1028_413.t10 221.719
R5 a_1028_413.n2 a_1028_413.t6 210.473
R6 a_1028_413.n7 a_1028_413.n6 194.899
R7 a_1028_413.n0 a_1028_413.t7 163.994
R8 a_1028_413.n2 a_1028_413.n1 154.418
R9 a_1028_413.n1 a_1028_413.t9 149.419
R10 a_1028_413.n1 a_1028_413.n0 144.6
R11 a_1028_413.n6 a_1028_413.n3 141.253
R12 a_1028_413.n4 a_1028_413.t3 119.607
R13 a_1028_413.n6 a_1028_413.n5 93.364
R14 a_1028_413.n4 a_1028_413.t1 63.321
R15 a_1028_413.t0 a_1028_413.n7 47.142
R16 a_1028_413.n7 a_1028_413.t4 47.142
R17 a_1028_413.n3 a_1028_413.n2 32.133
R18 VPWR.n34 VPWR.t7 429.335
R19 VPWR.n10 VPWR.t5 355.821
R20 VPWR.n6 VPWR.n5 312.281
R21 VPWR.n39 VPWR.n38 311.893
R22 VPWR.n20 VPWR.n19 307.239
R23 VPWR.n25 VPWR.n24 292.5
R24 VPWR.n2 VPWR.n0 183.421
R25 VPWR.n1 VPWR.t2 163.592
R26 VPWR.n24 VPWR.t8 91.464
R27 VPWR.n5 VPWR.t9 91.464
R28 VPWR.n24 VPWR.t6 86.773
R29 VPWR.n19 VPWR.t10 63.321
R30 VPWR.n19 VPWR.t11 63.321
R31 VPWR.n0 VPWR.t3 58.484
R32 VPWR.n38 VPWR.t4 41.554
R33 VPWR.n38 VPWR.t0 41.554
R34 VPWR.n5 VPWR.t1 32.833
R35 VPWR.n0 VPWR.t12 31.605
R36 VPWR.n4 VPWR.n3 4.65
R37 VPWR.n7 VPWR.n6 4.65
R38 VPWR.n9 VPWR.n8 4.65
R39 VPWR.n12 VPWR.n11 4.65
R40 VPWR.n14 VPWR.n13 4.65
R41 VPWR.n16 VPWR.n15 4.65
R42 VPWR.n18 VPWR.n17 4.65
R43 VPWR.n21 VPWR.n20 4.65
R44 VPWR.n23 VPWR.n22 4.65
R45 VPWR.n27 VPWR.n26 4.65
R46 VPWR.n29 VPWR.n28 4.65
R47 VPWR.n31 VPWR.n30 4.65
R48 VPWR.n33 VPWR.n32 4.65
R49 VPWR.n35 VPWR.n34 4.65
R50 VPWR.n37 VPWR.n36 4.65
R51 VPWR.n2 VPWR.n1 3.956
R52 VPWR.n40 VPWR.n39 3.932
R53 VPWR.n26 VPWR.n25 3.374
R54 VPWR.n11 VPWR.n10 0.814
R55 VPWR.n4 VPWR.n2 0.144
R56 VPWR.n40 VPWR.n37 0.137
R57 VPWR.n7 VPWR.n4 0.119
R58 VPWR.n9 VPWR.n7 0.119
R59 VPWR.n12 VPWR.n9 0.119
R60 VPWR.n14 VPWR.n12 0.119
R61 VPWR.n16 VPWR.n14 0.119
R62 VPWR.n18 VPWR.n16 0.119
R63 VPWR.n21 VPWR.n18 0.119
R64 VPWR.n23 VPWR.n21 0.119
R65 VPWR.n27 VPWR.n23 0.119
R66 VPWR.n29 VPWR.n27 0.119
R67 VPWR.n31 VPWR.n29 0.119
R68 VPWR.n33 VPWR.n31 0.119
R69 VPWR.n35 VPWR.n33 0.119
R70 VPWR.n37 VPWR.n35 0.119
R71 VPWR VPWR.n40 0.101
R72 a_1178_261.n0 a_1178_261.t2 372.273
R73 a_1178_261.t1 a_1178_261.n1 224.916
R74 a_1178_261.n1 a_1178_261.t0 198.825
R75 a_1178_261.n1 a_1178_261.n0 188.267
R76 a_1178_261.n0 a_1178_261.t3 167.991
R77 VPB.t1 VPB.t2 556.386
R78 VPB.t3 VPB.t1 556.386
R79 VPB.t11 VPB.t10 556.386
R80 VPB.t6 VPB.t8 556.386
R81 VPB.t4 VPB.t7 355.14
R82 VPB.t5 VPB.t14 319.626
R83 VPB.t7 VPB.t9 313.707
R84 VPB.t8 VPB.t15 287.071
R85 VPB.t10 VPB.t3 284.112
R86 VPB.t2 VPB.t16 281.152
R87 VPB.t13 VPB.t12 248.598
R88 VPB.t9 VPB.t13 248.598
R89 VPB.t15 VPB.t4 248.598
R90 VPB.t0 VPB.t6 248.598
R91 VPB.t14 VPB.t11 213.084
R92 VPB.t12 VPB.t5 213.084
R93 VPB VPB.t0 142.056
R94 a_652_21.n0 a_652_21.t3 387.959
R95 a_652_21.n2 a_652_21.n1 301.911
R96 a_652_21.n1 a_652_21.t2 241.655
R97 a_652_21.n0 a_652_21.t4 143.746
R98 a_652_21.n1 a_652_21.n0 111.072
R99 a_652_21.n2 a_652_21.t1 63.321
R100 a_652_21.t0 a_652_21.n2 63.321
R101 a_586_47.t0 a_586_47.t1 93.516
R102 VGND.n33 VGND.t5 188.008
R103 VGND.n17 VGND.t9 145.376
R104 VGND.n2 VGND.n0 123.539
R105 VGND.n1 VGND.t1 119.208
R106 VGND.n38 VGND.n37 107.239
R107 VGND.n6 VGND.n5 92.5
R108 VGND.n22 VGND.n21 92.5
R109 VGND.n21 VGND.t8 81.428
R110 VGND.n5 VGND.t6 67.142
R111 VGND.n5 VGND.t2 55.301
R112 VGND.n0 VGND.t3 54.285
R113 VGND.n21 VGND.t7 38.571
R114 VGND.n37 VGND.t4 38.571
R115 VGND.n37 VGND.t0 38.571
R116 VGND.n0 VGND.t10 25.934
R117 VGND.n4 VGND.n3 4.65
R118 VGND.n8 VGND.n7 4.65
R119 VGND.n10 VGND.n9 4.65
R120 VGND.n12 VGND.n11 4.65
R121 VGND.n14 VGND.n13 4.65
R122 VGND.n16 VGND.n15 4.65
R123 VGND.n18 VGND.n17 4.65
R124 VGND.n20 VGND.n19 4.65
R125 VGND.n24 VGND.n23 4.65
R126 VGND.n26 VGND.n25 4.65
R127 VGND.n28 VGND.n27 4.65
R128 VGND.n30 VGND.n29 4.65
R129 VGND.n32 VGND.n31 4.65
R130 VGND.n34 VGND.n33 4.65
R131 VGND.n36 VGND.n35 4.65
R132 VGND.n23 VGND.n22 4.511
R133 VGND.n2 VGND.n1 3.956
R134 VGND.n39 VGND.n38 3.932
R135 VGND.n7 VGND.n6 1.083
R136 VGND.n4 VGND.n2 0.144
R137 VGND.n39 VGND.n36 0.137
R138 VGND.n8 VGND.n4 0.119
R139 VGND.n10 VGND.n8 0.119
R140 VGND.n12 VGND.n10 0.119
R141 VGND.n14 VGND.n12 0.119
R142 VGND.n16 VGND.n14 0.119
R143 VGND.n18 VGND.n16 0.119
R144 VGND.n20 VGND.n18 0.119
R145 VGND.n24 VGND.n20 0.119
R146 VGND.n26 VGND.n24 0.119
R147 VGND.n28 VGND.n26 0.119
R148 VGND.n30 VGND.n28 0.119
R149 VGND.n32 VGND.n30 0.119
R150 VGND.n34 VGND.n32 0.119
R151 VGND.n36 VGND.n34 0.119
R152 VGND VGND.n39 0.101
R153 VNB.t13 VNB.t12 6082.35
R154 VNB.t6 VNB.t7 5346.86
R155 VNB.t3 VNB.t1 4860.85
R156 VNB.t1 VNB.t2 4545.05
R157 VNB VNB.t0 4270.59
R158 VNB.t10 VNB.t9 3688.24
R159 VNB.t8 VNB.t3 3570.15
R160 VNB.t4 VNB.t14 3558.82
R161 VNB.t15 VNB.t5 3105.88
R162 VNB.t14 VNB.t10 3105.88
R163 VNB.t0 VNB.t6 2717.65
R164 VNB.t11 VNB.t8 2329.41
R165 VNB.t5 VNB.t11 2329.41
R166 VNB.t12 VNB.t15 2329.41
R167 VNB.t9 VNB.t13 2329.41
R168 VNB.t2 VNB.t16 2296.7
R169 VNB.t7 VNB.t4 2280.14
R170 a_476_47.n4 a_476_47.n3 415.031
R171 a_476_47.n1 a_476_47.t6 344.897
R172 a_476_47.n2 a_476_47.t4 289.491
R173 a_476_47.n2 a_476_47.t5 228.146
R174 a_476_47.n3 a_476_47.n0 196.424
R175 a_476_47.n3 a_476_47.n2 138.78
R176 a_476_47.n2 a_476_47.n1 105.747
R177 a_476_47.n1 a_476_47.t7 93.186
R178 a_476_47.n0 a_476_47.t0 70
R179 a_476_47.n0 a_476_47.t2 63.333
R180 a_476_47.t1 a_476_47.n4 63.321
R181 a_476_47.n4 a_476_47.t3 63.321
R182 a_956_413.t0 a_956_413.t1 98.5
R183 a_193_47.n1 a_193_47.t5 538.583
R184 a_193_47.n0 a_193_47.t2 368.674
R185 a_193_47.t1 a_193_47.n3 278.596
R186 a_193_47.n0 a_193_47.t4 260.944
R187 a_193_47.n3 a_193_47.t0 150.413
R188 a_193_47.n1 a_193_47.t3 135.794
R189 a_193_47.n2 a_193_47.n0 25.663
R190 a_193_47.n2 a_193_47.n1 10.05
R191 a_193_47.n3 a_193_47.n2 6.187
R192 a_1136_413.t0 a_1136_413.t1 98.5
R193 CLK.n0 CLK.t0 270.454
R194 CLK.n0 CLK.t1 235.108
R195 CLK.n1 CLK.n0 76
R196 CLK.n1 CLK 7.68
R197 CLK CLK.n1 4.754
R198 a_27_47.n0 a_27_47.t3 344.354
R199 a_27_47.n3 a_27_47.t7 263.171
R200 a_27_47.t1 a_27_47.n5 243.779
R201 a_27_47.n1 a_27_47.t2 235.952
R202 a_27_47.n1 a_27_47.t4 232.166
R203 a_27_47.n3 a_27_47.t5 227.825
R204 a_27_47.n4 a_27_47.t0 195.494
R205 a_27_47.n0 a_27_47.t6 158.045
R206 a_27_47.n4 a_27_47.n3 76
R207 a_27_47.n5 a_27_47.n4 35.339
R208 a_27_47.n2 a_27_47.n0 6.892
R209 a_27_47.n5 a_27_47.n2 6.154
R210 a_27_47.n2 a_27_47.n1 4.65
R211 a_381_47.n1 a_381_47.n0 405.201
R212 a_381_47.n1 a_381_47.t0 95.021
R213 a_381_47.n0 a_381_47.t3 63.333
R214 a_381_47.t1 a_381_47.n1 31.613
R215 a_381_47.n0 a_381_47.t2 26.77
R216 a_1056_47.t0 a_1056_47.t1 60
R217 a_1786_47.t1 a_1786_47.n1 240.007
R218 a_1786_47.n0 a_1786_47.t3 239.038
R219 a_1786_47.n0 a_1786_47.t2 166.738
R220 a_1786_47.n1 a_1786_47.t0 149.883
R221 a_1786_47.n1 a_1786_47.n0 99.272
R222 Q.n1 Q.t1 207.372
R223 Q.n0 Q.t0 117.423
R224 Q Q.n0 66.695
R225 Q.n1 Q 9.019
R226 Q Q.n1 7.458
R227 Q.n0 Q 6.646
R228 D.n0 D.t0 264.028
R229 D.n0 D.t1 174.054
R230 D.n1 D.n0 76
R231 D.n1 D 8.585
R232 D D.n1 2.029
R233 SET_B.n0 SET_B.t0 401.403
R234 SET_B.n1 SET_B.t3 386.89
R235 SET_B.n1 SET_B.t1 148.348
R236 SET_B.n0 SET_B.t2 141.967
R237 SET_B.n2 SET_B.n1 98.281
R238 SET_B.n2 SET_B.n0 6.974
R239 SET_B SET_B.n2 3.246
R240 a_1224_47.t0 a_1224_47.t1 60
R241 a_562_413.t0 a_562_413.t1 211.071
R242 a_1296_47.t0 a_1296_47.t1 60
R243 Q_N.n2 Q_N.n1 292.5
R244 Q_N.n3 Q_N.n2 147.104
R245 Q_N.n0 Q_N.t0 82.726
R246 Q_N.n2 Q_N.t1 26.595
R247 Q_N.n3 Q_N 10.71
R248 Q_N.n1 Q_N 8.339
R249 Q_N Q_N.n0 7.01
R250 Q_N.n0 Q_N 5.757
R251 Q_N.n1 Q_N 4.848
R252 Q_N Q_N.n3 2.439
R253 a_796_47.t0 a_796_47.t1 60
C0 VPB VPWR 0.22fF
C1 VGND Q_N 0.17fF
C2 VPWR Q_N 0.22fF
C3 VPWR VGND 0.15fF
C4 SET_B VGND 0.48fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__dfsbp_2.ext - technology: sky130A

.subckt sky130_fd_sc_hd__dfsbp_2 Q Q_N D VPWR SET_B CLK VGND VNB VPB
X0 a_1178_261.t1 a_1028_413.t5 VPWR.t7 VPB.t8 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X1 VPWR.t8 a_1028_413.t6 a_1870_47.t1 VPB.t7 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 VGND.t10 a_652_21.t3 a_586_47.t0 VNB.t14 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3 a_1178_261.t0 a_1028_413.t7 VGND.t8 VNB.t11 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=540000u l=150000u
X4 VGND.t5 a_1028_413.t8 a_1870_47.t0 VNB.t10 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 a_956_413.t0 a_476_47.t4 VPWR.t2 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 a_1136_413.t0 a_193_47.t2 a_1028_413.t4 VPB.t17 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7 VPWR.t3 a_476_47.t5 a_652_21.t0 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 a_586_47.t1 a_193_47.t3 a_476_47.t3 VNB.t17 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X9 VPWR.t9 CLK.t0 a_27_47.t1 VPB.t9 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X10 a_476_47.t1 a_27_47.t2 a_381_47.t3 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X11 a_1056_47.t1 a_476_47.t6 VGND.t2 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12 a_381_47.t1 D.t0 VPWR.t1 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X13 a_652_21.t2 SET_B.t0 VPWR.t13 VPB.t15 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14 a_1224_47.t0 a_27_47.t3 a_1028_413.t1 VNB.t12 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15 a_562_413.t0 a_27_47.t4 a_476_47.t2 VPB.t10 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16 VPWR.t11 a_1870_47.t2 Q.t3 VPB.t13 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17 a_1028_413.t0 a_193_47.t4 a_1056_47.t0 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18 VGND.t4 a_1870_47.t3 Q.t1 VNB.t7 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X19 a_476_47.t0 a_193_47.t5 a_381_47.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20 a_1296_47.t1 a_1178_261.t2 a_1224_47.t1 VNB.t18 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21 Q_N.t1 a_1028_413.t9 VGND.t7 VNB.t9 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X22 a_193_47.t0 a_27_47.t5 VGND.t9 VNB.t13 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23 VPWR.t4 a_652_21.t4 a_562_413.t1 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24 VGND.t11 SET_B.t1 a_1296_47.t0 VNB.t15 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X25 Q.t0 a_1870_47.t4 VGND.t3 VNB.t6 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X26 a_1028_413.t2 a_27_47.t6 a_956_413.t1 VPB.t11 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X27 VPWR.t0 a_1178_261.t3 a_1136_413.t1 VPB.t18 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X28 Q.t2 a_1870_47.t5 VPWR.t12 VPB.t14 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X29 VPWR.t6 a_1028_413.t10 Q_N.t3 VPB.t6 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X30 VGND.t6 a_1028_413.t11 Q_N.t0 VNB.t8 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X31 a_193_47.t1 a_27_47.t7 VPWR.t10 VPB.t12 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X32 Q_N.t2 a_1028_413.t12 VPWR.t5 VPB.t5 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X33 a_796_47.t0 SET_B.t2 VGND.t12 VNB.t16 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X34 a_381_47.t2 D.t1 VGND.t1 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X35 a_652_21.t1 a_476_47.t7 a_796_47.t1 VNB.t5 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X36 VPWR.t14 SET_B.t3 a_1028_413.t3 VPB.t16 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X37 VGND.t0 CLK.t1 a_27_47.t0 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
R0 a_1028_413.n6 a_1028_413.t3 432.15
R1 a_1028_413.n6 a_1028_413.n5 319.003
R2 a_1028_413.n4 a_1028_413.t5 258.673
R3 a_1028_413.n0 a_1028_413.t6 221.719
R4 a_1028_413.n1 a_1028_413.t10 221.719
R5 a_1028_413.n2 a_1028_413.t12 221.719
R6 a_1028_413.n3 a_1028_413.t7 210.473
R7 a_1028_413.n8 a_1028_413.n7 194.899
R8 a_1028_413.n1 a_1028_413.n0 167.807
R9 a_1028_413.n3 a_1028_413.n2 154.418
R10 a_1028_413.n0 a_1028_413.t8 149.419
R11 a_1028_413.n1 a_1028_413.t11 149.419
R12 a_1028_413.n2 a_1028_413.t9 149.419
R13 a_1028_413.n7 a_1028_413.n4 141.253
R14 a_1028_413.n5 a_1028_413.t4 119.607
R15 a_1028_413.n7 a_1028_413.n6 93.364
R16 a_1028_413.n2 a_1028_413.n1 74.977
R17 a_1028_413.n5 a_1028_413.t2 63.321
R18 a_1028_413.n8 a_1028_413.t1 47.142
R19 a_1028_413.t0 a_1028_413.n8 47.142
R20 a_1028_413.n4 a_1028_413.n3 32.133
R21 VPWR.n44 VPWR.t1 429.335
R22 VPWR.n20 VPWR.t0 355.821
R23 VPWR.n16 VPWR.n15 312.281
R24 VPWR.n49 VPWR.n48 311.893
R25 VPWR.n30 VPWR.n29 307.239
R26 VPWR.n35 VPWR.n34 292.5
R27 VPWR.n0 VPWR.t11 198.56
R28 VPWR.n11 VPWR.t5 163.592
R29 VPWR.n7 VPWR.t6 152.716
R30 VPWR.n2 VPWR.n1 132.865
R31 VPWR.n34 VPWR.t13 91.464
R32 VPWR.n15 VPWR.t14 91.464
R33 VPWR.n34 VPWR.t4 86.773
R34 VPWR.n29 VPWR.t2 63.321
R35 VPWR.n29 VPWR.t3 63.321
R36 VPWR.n48 VPWR.t10 41.554
R37 VPWR.n48 VPWR.t9 41.554
R38 VPWR.n15 VPWR.t7 32.833
R39 VPWR.n1 VPWR.t12 26.595
R40 VPWR.n1 VPWR.t8 26.595
R41 VPWR.n4 VPWR.n3 4.65
R42 VPWR.n6 VPWR.n5 4.65
R43 VPWR.n8 VPWR.n7 4.65
R44 VPWR.n10 VPWR.n9 4.65
R45 VPWR.n12 VPWR.n11 4.65
R46 VPWR.n14 VPWR.n13 4.65
R47 VPWR.n17 VPWR.n16 4.65
R48 VPWR.n19 VPWR.n18 4.65
R49 VPWR.n22 VPWR.n21 4.65
R50 VPWR.n24 VPWR.n23 4.65
R51 VPWR.n26 VPWR.n25 4.65
R52 VPWR.n28 VPWR.n27 4.65
R53 VPWR.n31 VPWR.n30 4.65
R54 VPWR.n33 VPWR.n32 4.65
R55 VPWR.n37 VPWR.n36 4.65
R56 VPWR.n39 VPWR.n38 4.65
R57 VPWR.n41 VPWR.n40 4.65
R58 VPWR.n43 VPWR.n42 4.65
R59 VPWR.n45 VPWR.n44 4.65
R60 VPWR.n47 VPWR.n46 4.65
R61 VPWR.n50 VPWR.n49 3.932
R62 VPWR.n36 VPWR.n35 3.374
R63 VPWR.n21 VPWR.n20 0.814
R64 VPWR.n4 VPWR.n0 0.813
R65 VPWR.n3 VPWR.n2 0.376
R66 VPWR.n50 VPWR.n47 0.137
R67 VPWR.n6 VPWR.n4 0.119
R68 VPWR.n8 VPWR.n6 0.119
R69 VPWR.n10 VPWR.n8 0.119
R70 VPWR.n12 VPWR.n10 0.119
R71 VPWR.n14 VPWR.n12 0.119
R72 VPWR.n17 VPWR.n14 0.119
R73 VPWR.n19 VPWR.n17 0.119
R74 VPWR.n22 VPWR.n19 0.119
R75 VPWR.n24 VPWR.n22 0.119
R76 VPWR.n26 VPWR.n24 0.119
R77 VPWR.n28 VPWR.n26 0.119
R78 VPWR.n31 VPWR.n28 0.119
R79 VPWR.n33 VPWR.n31 0.119
R80 VPWR.n37 VPWR.n33 0.119
R81 VPWR.n39 VPWR.n37 0.119
R82 VPWR.n41 VPWR.n39 0.119
R83 VPWR.n43 VPWR.n41 0.119
R84 VPWR.n45 VPWR.n43 0.119
R85 VPWR.n47 VPWR.n45 0.119
R86 VPWR VPWR.n50 0.101
R87 a_1178_261.n0 a_1178_261.t2 372.273
R88 a_1178_261.t1 a_1178_261.n1 224.916
R89 a_1178_261.n1 a_1178_261.t0 198.825
R90 a_1178_261.n1 a_1178_261.n0 188.267
R91 a_1178_261.n0 a_1178_261.t3 167.991
R92 VPB.t6 VPB.t7 556.386
R93 VPB.t8 VPB.t5 556.386
R94 VPB.t18 VPB.t16 556.386
R95 VPB.t12 VPB.t1 556.386
R96 VPB.t10 VPB.t4 355.14
R97 VPB.t11 VPB.t17 319.626
R98 VPB.t4 VPB.t15 313.707
R99 VPB.t1 VPB.t0 287.071
R100 VPB.t16 VPB.t8 284.112
R101 VPB.t14 VPB.t13 248.598
R102 VPB.t7 VPB.t14 248.598
R103 VPB.t5 VPB.t6 248.598
R104 VPB.t3 VPB.t2 248.598
R105 VPB.t15 VPB.t3 248.598
R106 VPB.t0 VPB.t10 248.598
R107 VPB.t9 VPB.t12 248.598
R108 VPB.t17 VPB.t18 213.084
R109 VPB.t2 VPB.t11 213.084
R110 VPB VPB.t9 142.056
R111 a_1870_47.n1 a_1870_47.t5 212.079
R112 a_1870_47.n0 a_1870_47.t2 212.079
R113 a_1870_47.t1 a_1870_47.n2 144.121
R114 a_1870_47.n2 a_1870_47.t0 143.806
R115 a_1870_47.n1 a_1870_47.t4 139.779
R116 a_1870_47.n0 a_1870_47.t3 139.779
R117 a_1870_47.n2 a_1870_47.n1 100.436
R118 a_1870_47.n1 a_1870_47.n0 61.345
R119 a_652_21.n0 a_652_21.t3 387.959
R120 a_652_21.n2 a_652_21.n1 301.911
R121 a_652_21.n1 a_652_21.t1 241.655
R122 a_652_21.n0 a_652_21.t4 143.746
R123 a_652_21.n1 a_652_21.n0 111.072
R124 a_652_21.t0 a_652_21.n2 63.321
R125 a_652_21.n2 a_652_21.t2 63.321
R126 a_586_47.t0 a_586_47.t1 93.516
R127 VGND.n2 VGND.t4 195.9
R128 VGND.n41 VGND.t1 188.008
R129 VGND.n25 VGND.t2 145.376
R130 VGND.n9 VGND.t7 119.208
R131 VGND.n5 VGND.t6 109.821
R132 VGND.n46 VGND.n45 107.239
R133 VGND.n14 VGND.n13 92.5
R134 VGND.n30 VGND.n29 92.5
R135 VGND.n29 VGND.t10 81.428
R136 VGND.n13 VGND.t11 67.142
R137 VGND.n1 VGND.n0 64.067
R138 VGND.n13 VGND.t8 55.301
R139 VGND.n29 VGND.t12 38.571
R140 VGND.n45 VGND.t9 38.571
R141 VGND.n45 VGND.t0 38.571
R142 VGND.n0 VGND.t3 24.923
R143 VGND.n0 VGND.t5 24.923
R144 VGND.n4 VGND.n3 4.65
R145 VGND.n6 VGND.n5 4.65
R146 VGND.n8 VGND.n7 4.65
R147 VGND.n10 VGND.n9 4.65
R148 VGND.n12 VGND.n11 4.65
R149 VGND.n16 VGND.n15 4.65
R150 VGND.n18 VGND.n17 4.65
R151 VGND.n20 VGND.n19 4.65
R152 VGND.n22 VGND.n21 4.65
R153 VGND.n24 VGND.n23 4.65
R154 VGND.n26 VGND.n25 4.65
R155 VGND.n28 VGND.n27 4.65
R156 VGND.n32 VGND.n31 4.65
R157 VGND.n34 VGND.n33 4.65
R158 VGND.n36 VGND.n35 4.65
R159 VGND.n38 VGND.n37 4.65
R160 VGND.n40 VGND.n39 4.65
R161 VGND.n42 VGND.n41 4.65
R162 VGND.n44 VGND.n43 4.65
R163 VGND.n31 VGND.n30 4.511
R164 VGND.n47 VGND.n46 3.932
R165 VGND.n2 VGND.n1 3.82
R166 VGND.n15 VGND.n14 1.083
R167 VGND.n4 VGND.n2 0.243
R168 VGND.n47 VGND.n44 0.137
R169 VGND.n6 VGND.n4 0.119
R170 VGND.n8 VGND.n6 0.119
R171 VGND.n10 VGND.n8 0.119
R172 VGND.n12 VGND.n10 0.119
R173 VGND.n16 VGND.n12 0.119
R174 VGND.n18 VGND.n16 0.119
R175 VGND.n20 VGND.n18 0.119
R176 VGND.n22 VGND.n20 0.119
R177 VGND.n24 VGND.n22 0.119
R178 VGND.n26 VGND.n24 0.119
R179 VGND.n28 VGND.n26 0.119
R180 VGND.n32 VGND.n28 0.119
R181 VGND.n34 VGND.n32 0.119
R182 VGND.n36 VGND.n34 0.119
R183 VGND.n38 VGND.n36 0.119
R184 VGND.n40 VGND.n38 0.119
R185 VGND.n42 VGND.n40 0.119
R186 VGND.n44 VGND.n42 0.119
R187 VGND VGND.n47 0.101
R188 VNB.t5 VNB.t4 6082.35
R189 VNB.t13 VNB.t3 5346.86
R190 VNB.t11 VNB.t9 4860.85
R191 VNB.t8 VNB.t10 4545.05
R192 VNB VNB.t0 4270.59
R193 VNB.t14 VNB.t16 3688.24
R194 VNB.t15 VNB.t11 3570.15
R195 VNB.t2 VNB.t17 3558.82
R196 VNB.t1 VNB.t12 3105.88
R197 VNB.t17 VNB.t14 3105.88
R198 VNB.t0 VNB.t13 2717.65
R199 VNB.t18 VNB.t15 2329.41
R200 VNB.t12 VNB.t18 2329.41
R201 VNB.t4 VNB.t1 2329.41
R202 VNB.t16 VNB.t5 2329.41
R203 VNB.t3 VNB.t2 2280.14
R204 VNB.t6 VNB.t7 2030.77
R205 VNB.t10 VNB.t6 2030.77
R206 VNB.t9 VNB.t8 2030.77
R207 a_476_47.n4 a_476_47.n3 415.031
R208 a_476_47.n1 a_476_47.t6 344.897
R209 a_476_47.n2 a_476_47.t4 289.491
R210 a_476_47.n2 a_476_47.t5 228.146
R211 a_476_47.n3 a_476_47.n0 196.424
R212 a_476_47.n3 a_476_47.n2 138.78
R213 a_476_47.n2 a_476_47.n1 105.747
R214 a_476_47.n1 a_476_47.t7 93.186
R215 a_476_47.n0 a_476_47.t1 70
R216 a_476_47.n0 a_476_47.t3 63.333
R217 a_476_47.n4 a_476_47.t2 63.321
R218 a_476_47.t0 a_476_47.n4 63.321
R219 a_956_413.t0 a_956_413.t1 98.5
R220 a_193_47.n1 a_193_47.t5 538.583
R221 a_193_47.n0 a_193_47.t2 368.674
R222 a_193_47.t1 a_193_47.n3 278.596
R223 a_193_47.n0 a_193_47.t4 260.944
R224 a_193_47.n3 a_193_47.t0 150.413
R225 a_193_47.n1 a_193_47.t3 135.794
R226 a_193_47.n2 a_193_47.n0 25.663
R227 a_193_47.n2 a_193_47.n1 10.05
R228 a_193_47.n3 a_193_47.n2 6.187
R229 a_1136_413.t0 a_1136_413.t1 98.5
R230 CLK.n0 CLK.t0 270.454
R231 CLK.n0 CLK.t1 235.108
R232 CLK.n1 CLK.n0 76
R233 CLK.n1 CLK 7.68
R234 CLK CLK.n1 4.754
R235 a_27_47.n0 a_27_47.t3 344.354
R236 a_27_47.n3 a_27_47.t7 263.171
R237 a_27_47.t1 a_27_47.n5 243.779
R238 a_27_47.n1 a_27_47.t2 235.952
R239 a_27_47.n1 a_27_47.t4 232.166
R240 a_27_47.n3 a_27_47.t5 227.825
R241 a_27_47.n4 a_27_47.t0 195.494
R242 a_27_47.n0 a_27_47.t6 158.045
R243 a_27_47.n4 a_27_47.n3 76
R244 a_27_47.n5 a_27_47.n4 35.339
R245 a_27_47.n2 a_27_47.n0 6.892
R246 a_27_47.n5 a_27_47.n2 6.154
R247 a_27_47.n2 a_27_47.n1 4.65
R248 a_381_47.n1 a_381_47.n0 405.201
R249 a_381_47.n1 a_381_47.t0 95.021
R250 a_381_47.n0 a_381_47.t3 63.333
R251 a_381_47.t1 a_381_47.n1 31.613
R252 a_381_47.n0 a_381_47.t2 26.77
R253 a_1056_47.t0 a_1056_47.t1 60
R254 D.n0 D.t0 264.028
R255 D.n0 D.t1 174.054
R256 D.n1 D.n0 76
R257 D.n1 D 8.585
R258 D D.n1 2.029
R259 SET_B.n0 SET_B.t0 401.403
R260 SET_B.n1 SET_B.t3 386.89
R261 SET_B.n1 SET_B.t1 148.348
R262 SET_B.n0 SET_B.t2 141.967
R263 SET_B.n2 SET_B.n1 98.281
R264 SET_B.n2 SET_B.n0 6.974
R265 SET_B SET_B.n2 3.246
R266 a_1224_47.t0 a_1224_47.t1 60
R267 a_562_413.t0 a_562_413.t1 211.071
R268 Q.n3 Q.n2 292.5
R269 Q.n4 Q.n3 147.104
R270 Q.n1 Q.n0 92.5
R271 Q Q.n1 48.16
R272 Q.n2 Q 33.088
R273 Q.n3 Q.t3 26.595
R274 Q.n3 Q.t2 26.595
R275 Q.n0 Q.t1 24.923
R276 Q.n0 Q.t0 24.923
R277 Q.n4 Q 10.71
R278 Q.n1 Q 6.912
R279 Q.n2 Q 4.654
R280 Q Q.n4 2.439
R281 a_1296_47.t0 a_1296_47.t1 60
R282 Q_N.n3 Q_N.n2 292.5
R283 Q_N.n4 Q_N.n3 147.104
R284 Q_N Q_N.n0 93.469
R285 Q_N.n1 Q_N.n0 92.5
R286 Q_N.n3 Q_N.t3 26.595
R287 Q_N.n3 Q_N.t2 26.595
R288 Q_N.n0 Q_N.t0 24.923
R289 Q_N.n0 Q_N.t1 24.923
R290 Q_N.n1 Q_N 12.218
R291 Q_N.n4 Q_N 10.71
R292 Q_N.n2 Q_N 8.339
R293 Q_N.n2 Q_N 4.848
R294 Q_N Q_N.n4 2.439
R295 Q_N Q_N.n1 0.969
R296 a_796_47.t0 a_796_47.t1 60
C0 VPWR VGND 0.17fF
C1 SET_B VGND 0.48fF
C2 VPB VPWR 0.23fF
C3 VGND Q 0.22fF
C4 VGND Q_N 0.28fF
C5 VPWR Q 0.38fF
C6 VPWR Q_N 0.39fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__dfstp_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__dfstp_1 D VPWR Q SET_B CLK VGND VNB VPB
X0 VGND.t4 a_652_21.t3 a_586_47.t0 VNB.t5 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1 a_956_413.t0 a_476_47.t4 VPWR.t4 VPB.t6 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 VPWR.t3 a_476_47.t5 a_652_21.t1 VPB.t5 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3 a_586_47.t1 a_193_47.t2 a_476_47.t0 VNB.t7 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X4 VPWR.t8 CLK.t0 a_27_47.t1 VPB.t12 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X5 a_476_47.t2 a_27_47.t2 a_381_47.t0 VNB.t10 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X6 a_1056_47.t0 a_476_47.t6 VGND.t8 VNB.t13 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7 a_381_47.t1 D.t0 VPWR.t5 VPB.t7 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X8 a_652_21.t0 SET_B.t0 VPWR.t1 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9 a_1224_47.t0 a_27_47.t3 a_1032_413.t0 VNB.t11 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10 a_562_413.t0 a_27_47.t4 a_476_47.t3 VPB.t9 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11 VGND.t2 a_1032_413.t5 a_1602_47.t0 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12 VPWR.t6 a_1182_261.t2 a_1140_413.t0 VPB.t8 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13 Q.t1 a_1602_47.t2 VPWR.t11 VPB.t15 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14 a_1032_413.t4 a_193_47.t3 a_1056_47.t1 VNB.t8 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15 a_476_47.t1 a_193_47.t4 a_381_47.t3 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16 a_1296_47.t1 a_1182_261.t3 a_1224_47.t1 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17 a_193_47.t0 a_27_47.t5 VGND.t7 VNB.t12 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18 VPWR.t2 a_652_21.t4 a_562_413.t1 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19 VPWR.t0 SET_B.t1 a_1032_413.t2 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20 a_1032_413.t1 a_27_47.t6 a_956_413.t1 VPB.t10 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21 a_1182_261.t1 a_1032_413.t6 VPWR.t9 VPB.t13 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X22 Q.t0 a_1602_47.t3 VGND.t5 VNB.t6 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X23 a_193_47.t1 a_27_47.t7 VPWR.t7 VPB.t11 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X24 a_1140_413.t1 a_193_47.t5 a_1032_413.t3 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X25 VPWR.t10 a_1032_413.t7 a_1602_47.t1 VPB.t14 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X26 a_796_47.t0 SET_B.t2 VGND.t0 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X27 a_381_47.t2 D.t1 VGND.t6 VNB.t9 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X28 a_1182_261.t0 a_1032_413.t8 VGND.t9 VNB.t15 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=540000u l=150000u
X29 a_652_21.t2 a_476_47.t7 a_796_47.t1 VNB.t14 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X30 VGND.t3 CLK.t1 a_27_47.t0 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X31 VGND.t1 SET_B.t3 a_1296_47.t0 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
R0 a_652_21.n0 a_652_21.t3 387.959
R1 a_652_21.n2 a_652_21.n1 301.911
R2 a_652_21.n1 a_652_21.t2 235.545
R3 a_652_21.n0 a_652_21.t4 143.746
R4 a_652_21.n1 a_652_21.n0 111.072
R5 a_652_21.n2 a_652_21.t1 63.321
R6 a_652_21.t0 a_652_21.n2 63.321
R7 a_586_47.t0 a_586_47.t1 93.516
R8 VGND.n28 VGND.t6 188.008
R9 VGND.n12 VGND.t8 146.271
R10 VGND.n3 VGND.n0 113.286
R11 VGND.n33 VGND.n32 107.239
R12 VGND.n2 VGND.n1 92.5
R13 VGND.n17 VGND.n16 92.5
R14 VGND.n16 VGND.t4 81.428
R15 VGND.n1 VGND.t1 67.142
R16 VGND.n1 VGND.t9 55.301
R17 VGND.n0 VGND.t2 54.285
R18 VGND.n16 VGND.t0 38.571
R19 VGND.n32 VGND.t7 38.571
R20 VGND.n32 VGND.t3 38.571
R21 VGND.n0 VGND.t5 25.934
R22 VGND.n5 VGND.n4 4.65
R23 VGND.n7 VGND.n6 4.65
R24 VGND.n9 VGND.n8 4.65
R25 VGND.n11 VGND.n10 4.65
R26 VGND.n13 VGND.n12 4.65
R27 VGND.n15 VGND.n14 4.65
R28 VGND.n19 VGND.n18 4.65
R29 VGND.n21 VGND.n20 4.65
R30 VGND.n23 VGND.n22 4.65
R31 VGND.n25 VGND.n24 4.65
R32 VGND.n27 VGND.n26 4.65
R33 VGND.n29 VGND.n28 4.65
R34 VGND.n31 VGND.n30 4.65
R35 VGND.n3 VGND.n2 4.623
R36 VGND.n18 VGND.n17 4.511
R37 VGND.n34 VGND.n33 3.932
R38 VGND.n5 VGND.n3 0.146
R39 VGND.n34 VGND.n31 0.137
R40 VGND VGND.n34 0.123
R41 VGND.n7 VGND.n5 0.119
R42 VGND.n9 VGND.n7 0.119
R43 VGND.n11 VGND.n9 0.119
R44 VGND.n13 VGND.n11 0.119
R45 VGND.n15 VGND.n13 0.119
R46 VGND.n19 VGND.n15 0.119
R47 VGND.n21 VGND.n19 0.119
R48 VGND.n23 VGND.n21 0.119
R49 VGND.n25 VGND.n23 0.119
R50 VGND.n27 VGND.n25 0.119
R51 VGND.n29 VGND.n27 0.119
R52 VGND.n31 VGND.n29 0.119
R53 VNB.t14 VNB.t13 6082.35
R54 VNB.t12 VNB.t9 5346.86
R55 VNB.t15 VNB.t2 5170
R56 VNB VNB.t4 4270.59
R57 VNB.t5 VNB.t0 3688.24
R58 VNB.t1 VNB.t15 3570.15
R59 VNB.t10 VNB.t7 3558.82
R60 VNB.t8 VNB.t11 3105.88
R61 VNB.t7 VNB.t5 3105.88
R62 VNB.t4 VNB.t12 2717.65
R63 VNB.t3 VNB.t1 2458.82
R64 VNB.t11 VNB.t3 2329.41
R65 VNB.t13 VNB.t8 2329.41
R66 VNB.t0 VNB.t14 2329.41
R67 VNB.t9 VNB.t10 2280.14
R68 VNB.t2 VNB.t6 342.561
R69 a_476_47.n4 a_476_47.n3 415.031
R70 a_476_47.n1 a_476_47.t6 344.897
R71 a_476_47.n2 a_476_47.t4 289.491
R72 a_476_47.n2 a_476_47.t5 228.146
R73 a_476_47.n3 a_476_47.n0 196.424
R74 a_476_47.n3 a_476_47.n2 138.78
R75 a_476_47.n2 a_476_47.n1 105.747
R76 a_476_47.n1 a_476_47.t7 93.186
R77 a_476_47.n0 a_476_47.t2 70
R78 a_476_47.n0 a_476_47.t0 63.333
R79 a_476_47.n4 a_476_47.t3 63.321
R80 a_476_47.t1 a_476_47.n4 63.321
R81 VPWR.n30 VPWR.t5 429.335
R82 VPWR.n6 VPWR.t6 355.821
R83 VPWR.n1 VPWR.n0 312.281
R84 VPWR.n35 VPWR.n34 311.893
R85 VPWR.n16 VPWR.n15 307.239
R86 VPWR.n21 VPWR.n20 292.5
R87 VPWR.n3 VPWR.n2 170.753
R88 VPWR.n20 VPWR.t1 91.464
R89 VPWR.n0 VPWR.t0 91.464
R90 VPWR.n20 VPWR.t2 86.773
R91 VPWR.n15 VPWR.t4 63.321
R92 VPWR.n15 VPWR.t3 63.321
R93 VPWR.n2 VPWR.t10 58.484
R94 VPWR.n34 VPWR.t7 41.554
R95 VPWR.n34 VPWR.t8 41.554
R96 VPWR.n0 VPWR.t9 32.833
R97 VPWR.n2 VPWR.t11 31.605
R98 VPWR.n5 VPWR.n4 4.65
R99 VPWR.n8 VPWR.n7 4.65
R100 VPWR.n10 VPWR.n9 4.65
R101 VPWR.n12 VPWR.n11 4.65
R102 VPWR.n14 VPWR.n13 4.65
R103 VPWR.n17 VPWR.n16 4.65
R104 VPWR.n19 VPWR.n18 4.65
R105 VPWR.n23 VPWR.n22 4.65
R106 VPWR.n25 VPWR.n24 4.65
R107 VPWR.n27 VPWR.n26 4.65
R108 VPWR.n29 VPWR.n28 4.65
R109 VPWR.n31 VPWR.n30 4.65
R110 VPWR.n33 VPWR.n32 4.65
R111 VPWR.n36 VPWR.n35 3.932
R112 VPWR.n3 VPWR.n1 3.795
R113 VPWR.n22 VPWR.n21 3.374
R114 VPWR.n7 VPWR.n6 0.349
R115 VPWR.n5 VPWR.n3 0.151
R116 VPWR.n36 VPWR.n33 0.137
R117 VPWR VPWR.n36 0.123
R118 VPWR.n8 VPWR.n5 0.119
R119 VPWR.n10 VPWR.n8 0.119
R120 VPWR.n12 VPWR.n10 0.119
R121 VPWR.n14 VPWR.n12 0.119
R122 VPWR.n17 VPWR.n14 0.119
R123 VPWR.n19 VPWR.n17 0.119
R124 VPWR.n23 VPWR.n19 0.119
R125 VPWR.n25 VPWR.n23 0.119
R126 VPWR.n27 VPWR.n25 0.119
R127 VPWR.n29 VPWR.n27 0.119
R128 VPWR.n31 VPWR.n29 0.119
R129 VPWR.n33 VPWR.n31 0.119
R130 a_956_413.t0 a_956_413.t1 107.88
R131 VPB.t13 VPB.t14 556.386
R132 VPB.t8 VPB.t1 556.386
R133 VPB.t11 VPB.t7 556.386
R134 VPB.t9 VPB.t3 355.14
R135 VPB.t10 VPB.t0 319.626
R136 VPB.t3 VPB.t2 313.707
R137 VPB.t7 VPB.t4 287.071
R138 VPB.t1 VPB.t13 284.112
R139 VPB.t14 VPB.t15 281.152
R140 VPB.t5 VPB.t6 248.598
R141 VPB.t2 VPB.t5 248.598
R142 VPB.t4 VPB.t9 248.598
R143 VPB.t12 VPB.t11 248.598
R144 VPB.t6 VPB.t10 224.922
R145 VPB.t0 VPB.t8 213.084
R146 VPB VPB.t12 142.056
R147 a_193_47.n1 a_193_47.t4 538.597
R148 a_193_47.n0 a_193_47.t5 379.019
R149 a_193_47.t1 a_193_47.n3 278.596
R150 a_193_47.n0 a_193_47.t3 261.35
R151 a_193_47.n3 a_193_47.t0 150.413
R152 a_193_47.n1 a_193_47.t2 135.786
R153 a_193_47.n2 a_193_47.n0 30.468
R154 a_193_47.n2 a_193_47.n1 10.203
R155 a_193_47.n3 a_193_47.n2 6.202
R156 CLK.n0 CLK.t0 270.454
R157 CLK.n0 CLK.t1 235.108
R158 CLK.n1 CLK.n0 76
R159 CLK.n1 CLK 7.68
R160 CLK CLK.n1 4.754
R161 a_27_47.n0 a_27_47.t3 345.62
R162 a_27_47.n3 a_27_47.t7 263.171
R163 a_27_47.t1 a_27_47.n5 243.779
R164 a_27_47.n1 a_27_47.t2 236.795
R165 a_27_47.n1 a_27_47.t4 231.324
R166 a_27_47.n3 a_27_47.t5 227.825
R167 a_27_47.n4 a_27_47.t0 195.494
R168 a_27_47.n0 a_27_47.t6 159.8
R169 a_27_47.n4 a_27_47.n3 76
R170 a_27_47.n5 a_27_47.n4 35.339
R171 a_27_47.n2 a_27_47.n0 7.19
R172 a_27_47.n5 a_27_47.n2 6.207
R173 a_27_47.n2 a_27_47.n1 4.65
R174 a_381_47.n1 a_381_47.n0 405.201
R175 a_381_47.n1 a_381_47.t3 95.021
R176 a_381_47.n0 a_381_47.t0 63.333
R177 a_381_47.t1 a_381_47.n1 31.613
R178 a_381_47.n0 a_381_47.t2 26.77
R179 a_1056_47.t0 a_1056_47.t1 60
R180 D.n0 D.t0 264.028
R181 D.n0 D.t1 174.054
R182 D.n1 D.n0 76
R183 D.n1 D 8.585
R184 D D.n1 2.029
R185 SET_B.n0 SET_B.t0 396.818
R186 SET_B.n1 SET_B.t1 386.89
R187 SET_B.n1 SET_B.t3 148.348
R188 SET_B.n0 SET_B.t2 134.069
R189 SET_B.n2 SET_B.n1 100.452
R190 SET_B.n2 SET_B.n0 7.921
R191 SET_B SET_B.n2 3.245
R192 a_1032_413.n3 a_1032_413.t2 433.656
R193 a_1032_413.n3 a_1032_413.n2 317.979
R194 a_1032_413.n0 a_1032_413.t7 237.786
R195 a_1032_413.n0 a_1032_413.t5 208.866
R196 a_1032_413.n1 a_1032_413.t6 205.653
R197 a_1032_413.n5 a_1032_413.n4 194.899
R198 a_1032_413.n1 a_1032_413.t8 189.586
R199 a_1032_413.n4 a_1032_413.n1 153.713
R200 a_1032_413.n1 a_1032_413.n0 137.296
R201 a_1032_413.n2 a_1032_413.t3 119.607
R202 a_1032_413.n4 a_1032_413.n3 93.364
R203 a_1032_413.n2 a_1032_413.t1 63.321
R204 a_1032_413.t0 a_1032_413.n5 47.142
R205 a_1032_413.n5 a_1032_413.t4 47.142
R206 a_1224_47.t0 a_1224_47.t1 60
R207 a_562_413.t0 a_562_413.t1 211.071
R208 a_1602_47.t1 a_1602_47.n1 247.33
R209 a_1602_47.n0 a_1602_47.t2 241.534
R210 a_1602_47.n0 a_1602_47.t3 169.234
R211 a_1602_47.n1 a_1602_47.t0 155.903
R212 a_1602_47.n1 a_1602_47.n0 98.884
R213 a_1182_261.n0 a_1182_261.t3 374.754
R214 a_1182_261.t1 a_1182_261.n1 224.916
R215 a_1182_261.n1 a_1182_261.t0 198.825
R216 a_1182_261.n1 a_1182_261.n0 189.773
R217 a_1182_261.n0 a_1182_261.t2 169.453
R218 a_1140_413.t0 a_1140_413.t1 98.5
R219 Q.n1 Q.t1 207.309
R220 Q.n0 Q.t0 117.423
R221 Q Q.n0 75.962
R222 Q.n0 Q 10.29
R223 Q.n1 Q 9.192
R224 Q Q.n1 7.602
R225 a_1296_47.t0 a_1296_47.t1 65.714
R226 a_796_47.t0 a_796_47.t1 60
C0 VPB VPWR 0.20fF
C1 VPWR VGND 0.11fF
C2 SET_B VGND 0.48fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__dfstp_2.ext - technology: sky130A

.subckt sky130_fd_sc_hd__dfstp_2 Q D VPWR SET_B CLK VGND VNB VPB
X0 VGND.t7 a_652_21.t3 a_586_47.t1 VNB.t12 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1 a_956_413.t1 a_476_47.t4 VPWR.t11 VPB.t16 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 a_1136_413.t0 a_193_47.t2 a_1028_413.t2 VPB.t8 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3 VPWR.t12 a_476_47.t5 a_652_21.t0 VPB.t15 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 a_586_47.t0 a_193_47.t3 a_476_47.t2 VNB.t9 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X5 a_1228_47.t0 a_27_47.t2 a_1028_413.t0 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 VPWR.t10 CLK.t0 a_27_47.t0 VPB.t14 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X7 a_476_47.t0 a_27_47.t3 a_381_47.t3 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X8 a_1056_47.t1 a_476_47.t6 VGND.t2 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9 a_381_47.t1 D.t0 VPWR.t3 VPB.t5 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X10 a_652_21.t1 SET_B.t0 VPWR.t8 VPB.t12 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11 VPWR.t4 a_1602_47.t2 Q.t1 VPB.t6 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 a_562_413.t0 a_27_47.t4 a_476_47.t1 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13 VGND.t0 a_1028_413.t5 a_1602_47.t1 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14 VGND.t5 a_1602_47.t3 Q.t3 VNB.t7 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X15 Q.t0 a_1602_47.t4 VPWR.t5 VPB.t7 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16 a_1028_413.t3 a_193_47.t4 a_1056_47.t0 VNB.t10 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17 a_476_47.t3 a_193_47.t5 a_381_47.t0 VPB.t9 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18 a_193_47.t0 a_27_47.t5 VGND.t3 VNB.t5 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19 VPWR.t0 a_1028_413.t6 a_1602_47.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X20 VPWR.t7 a_652_21.t4 a_562_413.t1 VPB.t11 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21 Q.t2 a_1602_47.t5 VGND.t6 VNB.t8 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X22 a_1028_413.t1 a_27_47.t6 a_956_413.t0 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23 VPWR.t6 a_1178_261.t2 a_1136_413.t1 VPB.t10 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24 a_193_47.t1 a_27_47.t7 VPWR.t2 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X25 a_1178_261.t0 a_1028_413.t7 VPWR.t1 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X26 a_796_47.t0 SET_B.t1 VGND.t8 VNB.t13 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X27 a_1300_47.t1 a_1178_261.t3 a_1228_47.t1 VNB.t11 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X28 a_381_47.t2 D.t1 VGND.t4 VNB.t6 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X29 a_1178_261.t1 a_1028_413.t8 VGND.t1 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=540000u l=150000u
X30 a_652_21.t2 a_476_47.t7 a_796_47.t1 VNB.t15 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X31 VPWR.t9 SET_B.t2 a_1028_413.t4 VPB.t13 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X32 VGND.t10 CLK.t1 a_27_47.t1 VNB.t16 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X33 VGND.t9 SET_B.t3 a_1300_47.t0 VNB.t14 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
R0 a_652_21.n0 a_652_21.t3 387.959
R1 a_652_21.n2 a_652_21.n1 301.911
R2 a_652_21.n1 a_652_21.t2 241.655
R3 a_652_21.n0 a_652_21.t4 143.746
R4 a_652_21.n1 a_652_21.n0 111.072
R5 a_652_21.t0 a_652_21.n2 63.321
R6 a_652_21.n2 a_652_21.t1 63.321
R7 a_586_47.t1 a_586_47.t0 93.516
R8 VGND.n2 VGND.t5 197.675
R9 VGND.n35 VGND.t4 188.008
R10 VGND.n19 VGND.t2 146.271
R11 VGND.n40 VGND.n39 107.239
R12 VGND.n8 VGND.n7 92.5
R13 VGND.n24 VGND.n23 92.5
R14 VGND.n23 VGND.t7 81.428
R15 VGND.n7 VGND.t9 67.142
R16 VGND.n1 VGND.n0 64.067
R17 VGND.n7 VGND.t1 55.301
R18 VGND.n23 VGND.t8 38.571
R19 VGND.n39 VGND.t3 38.571
R20 VGND.n39 VGND.t10 38.571
R21 VGND.n0 VGND.t6 24.923
R22 VGND.n0 VGND.t0 24.923
R23 VGND.n4 VGND.n3 4.65
R24 VGND.n6 VGND.n5 4.65
R25 VGND.n10 VGND.n9 4.65
R26 VGND.n12 VGND.n11 4.65
R27 VGND.n14 VGND.n13 4.65
R28 VGND.n16 VGND.n15 4.65
R29 VGND.n18 VGND.n17 4.65
R30 VGND.n20 VGND.n19 4.65
R31 VGND.n22 VGND.n21 4.65
R32 VGND.n26 VGND.n25 4.65
R33 VGND.n28 VGND.n27 4.65
R34 VGND.n30 VGND.n29 4.65
R35 VGND.n32 VGND.n31 4.65
R36 VGND.n34 VGND.n33 4.65
R37 VGND.n36 VGND.n35 4.65
R38 VGND.n38 VGND.n37 4.65
R39 VGND.n25 VGND.n24 4.511
R40 VGND.n41 VGND.n40 3.932
R41 VGND.n2 VGND.n1 3.74
R42 VGND.n9 VGND.n8 0.689
R43 VGND.n4 VGND.n2 0.247
R44 VGND.n41 VGND.n38 0.137
R45 VGND VGND.n41 0.123
R46 VGND.n6 VGND.n4 0.119
R47 VGND.n10 VGND.n6 0.119
R48 VGND.n12 VGND.n10 0.119
R49 VGND.n14 VGND.n12 0.119
R50 VGND.n16 VGND.n14 0.119
R51 VGND.n18 VGND.n16 0.119
R52 VGND.n20 VGND.n18 0.119
R53 VGND.n22 VGND.n20 0.119
R54 VGND.n26 VGND.n22 0.119
R55 VGND.n28 VGND.n26 0.119
R56 VGND.n30 VGND.n28 0.119
R57 VGND.n32 VGND.n30 0.119
R58 VGND.n34 VGND.n32 0.119
R59 VGND.n36 VGND.n34 0.119
R60 VGND.n38 VGND.n36 0.119
R61 VNB.t15 VNB.t2 6082.35
R62 VNB.t5 VNB.t6 5346.86
R63 VNB.t1 VNB.t0 4860.85
R64 VNB VNB.t16 4270.59
R65 VNB.t12 VNB.t13 3688.24
R66 VNB.t14 VNB.t1 3570.15
R67 VNB.t4 VNB.t9 3558.82
R68 VNB.t10 VNB.t3 3235.29
R69 VNB.t9 VNB.t12 3105.88
R70 VNB.t16 VNB.t5 2717.65
R71 VNB.t11 VNB.t14 2329.41
R72 VNB.t3 VNB.t11 2329.41
R73 VNB.t2 VNB.t10 2329.41
R74 VNB.t13 VNB.t15 2329.41
R75 VNB.t6 VNB.t4 2280.14
R76 VNB.t8 VNB.t7 2030.77
R77 VNB.t0 VNB.t8 2030.77
R78 a_476_47.n4 a_476_47.n3 415.031
R79 a_476_47.n1 a_476_47.t6 344.897
R80 a_476_47.n2 a_476_47.t4 289.491
R81 a_476_47.n2 a_476_47.t5 228.146
R82 a_476_47.n3 a_476_47.n0 196.424
R83 a_476_47.n3 a_476_47.n2 138.78
R84 a_476_47.n2 a_476_47.n1 105.747
R85 a_476_47.n1 a_476_47.t7 93.186
R86 a_476_47.n0 a_476_47.t0 70
R87 a_476_47.n0 a_476_47.t2 63.333
R88 a_476_47.t1 a_476_47.n4 63.321
R89 a_476_47.n4 a_476_47.t3 63.321
R90 VPWR.n38 VPWR.t3 429.335
R91 VPWR.n14 VPWR.t6 355.821
R92 VPWR.n10 VPWR.n9 312.281
R93 VPWR.n43 VPWR.n42 311.893
R94 VPWR.n24 VPWR.n23 307.239
R95 VPWR.n29 VPWR.n28 292.5
R96 VPWR.n0 VPWR.t4 199.193
R97 VPWR.n2 VPWR.n1 132.865
R98 VPWR.n28 VPWR.t8 91.464
R99 VPWR.n9 VPWR.t9 89.119
R100 VPWR.n28 VPWR.t7 86.773
R101 VPWR.n23 VPWR.t11 63.321
R102 VPWR.n23 VPWR.t12 63.321
R103 VPWR.n42 VPWR.t2 41.554
R104 VPWR.n42 VPWR.t10 41.554
R105 VPWR.n9 VPWR.t1 34.005
R106 VPWR.n1 VPWR.t5 26.595
R107 VPWR.n1 VPWR.t0 26.595
R108 VPWR.n4 VPWR.n3 4.65
R109 VPWR.n6 VPWR.n5 4.65
R110 VPWR.n8 VPWR.n7 4.65
R111 VPWR.n11 VPWR.n10 4.65
R112 VPWR.n13 VPWR.n12 4.65
R113 VPWR.n16 VPWR.n15 4.65
R114 VPWR.n18 VPWR.n17 4.65
R115 VPWR.n20 VPWR.n19 4.65
R116 VPWR.n22 VPWR.n21 4.65
R117 VPWR.n25 VPWR.n24 4.65
R118 VPWR.n27 VPWR.n26 4.65
R119 VPWR.n31 VPWR.n30 4.65
R120 VPWR.n33 VPWR.n32 4.65
R121 VPWR.n35 VPWR.n34 4.65
R122 VPWR.n37 VPWR.n36 4.65
R123 VPWR.n39 VPWR.n38 4.65
R124 VPWR.n41 VPWR.n40 4.65
R125 VPWR.n44 VPWR.n43 3.932
R126 VPWR.n3 VPWR.n2 3.388
R127 VPWR.n30 VPWR.n29 3.374
R128 VPWR.n15 VPWR.n14 0.814
R129 VPWR.n4 VPWR.n0 0.753
R130 VPWR.n44 VPWR.n41 0.137
R131 VPWR VPWR.n44 0.123
R132 VPWR.n6 VPWR.n4 0.119
R133 VPWR.n8 VPWR.n6 0.119
R134 VPWR.n11 VPWR.n8 0.119
R135 VPWR.n13 VPWR.n11 0.119
R136 VPWR.n16 VPWR.n13 0.119
R137 VPWR.n18 VPWR.n16 0.119
R138 VPWR.n20 VPWR.n18 0.119
R139 VPWR.n22 VPWR.n20 0.119
R140 VPWR.n25 VPWR.n22 0.119
R141 VPWR.n27 VPWR.n25 0.119
R142 VPWR.n31 VPWR.n27 0.119
R143 VPWR.n33 VPWR.n31 0.119
R144 VPWR.n35 VPWR.n33 0.119
R145 VPWR.n37 VPWR.n35 0.119
R146 VPWR.n39 VPWR.n37 0.119
R147 VPWR.n41 VPWR.n39 0.119
R148 a_956_413.t0 a_956_413.t1 98.5
R149 VPB.t1 VPB.t0 571.183
R150 VPB.t10 VPB.t13 556.386
R151 VPB.t4 VPB.t5 556.386
R152 VPB.t2 VPB.t11 355.14
R153 VPB.t3 VPB.t8 319.626
R154 VPB.t11 VPB.t12 313.707
R155 VPB.t5 VPB.t9 287.071
R156 VPB.t13 VPB.t1 281.152
R157 VPB.t7 VPB.t6 248.598
R158 VPB.t0 VPB.t7 248.598
R159 VPB.t15 VPB.t16 248.598
R160 VPB.t12 VPB.t15 248.598
R161 VPB.t9 VPB.t2 248.598
R162 VPB.t14 VPB.t4 248.598
R163 VPB.t8 VPB.t10 213.084
R164 VPB.t16 VPB.t3 213.084
R165 VPB VPB.t14 142.056
R166 a_193_47.n1 a_193_47.t5 538.583
R167 a_193_47.n0 a_193_47.t2 373.664
R168 a_193_47.t1 a_193_47.n3 277.278
R169 a_193_47.n0 a_193_47.t4 264.028
R170 a_193_47.n3 a_193_47.t0 150.131
R171 a_193_47.n1 a_193_47.t3 135.794
R172 a_193_47.n2 a_193_47.n0 27.501
R173 a_193_47.n2 a_193_47.n1 10.05
R174 a_193_47.n3 a_193_47.n2 6.187
R175 a_1028_413.n4 a_1028_413.t4 433.656
R176 a_1028_413.n2 a_1028_413.t7 399.218
R177 a_1028_413.n4 a_1028_413.n3 317.979
R178 a_1028_413.n6 a_1028_413.n5 194.899
R179 a_1028_413.n1 a_1028_413.t8 189.586
R180 a_1028_413.n0 a_1028_413.t6 184.766
R181 a_1028_413.n0 a_1028_413.t5 171.913
R182 a_1028_413.n1 a_1028_413.n0 143.834
R183 a_1028_413.n5 a_1028_413.n2 141.636
R184 a_1028_413.n3 a_1028_413.t2 119.607
R185 a_1028_413.n5 a_1028_413.n4 94.87
R186 a_1028_413.n3 a_1028_413.t1 63.321
R187 a_1028_413.t0 a_1028_413.n6 52.857
R188 a_1028_413.n6 a_1028_413.t3 47.142
R189 a_1028_413.n2 a_1028_413.n1 12.241
R190 a_1136_413.t0 a_1136_413.t1 98.5
R191 a_27_47.n0 a_27_47.t2 344.032
R192 a_27_47.n3 a_27_47.t7 262.942
R193 a_27_47.t0 a_27_47.n5 238.885
R194 a_27_47.n1 a_27_47.t3 235.952
R195 a_27_47.n1 a_27_47.t4 232.166
R196 a_27_47.n3 a_27_47.t5 227.596
R197 a_27_47.n4 a_27_47.t1 189.645
R198 a_27_47.n0 a_27_47.t6 158.045
R199 a_27_47.n4 a_27_47.n3 76
R200 a_27_47.n5 a_27_47.n4 35.339
R201 a_27_47.n2 a_27_47.n0 6.892
R202 a_27_47.n5 a_27_47.n2 6.189
R203 a_27_47.n2 a_27_47.n1 4.65
R204 a_1228_47.t0 a_1228_47.t1 60
R205 CLK.n0 CLK.t0 272.06
R206 CLK.n0 CLK.t1 236.714
R207 CLK.n1 CLK.n0 76
R208 CLK.n1 CLK 7.68
R209 CLK CLK.n1 4.754
R210 a_381_47.n1 a_381_47.n0 405.201
R211 a_381_47.n1 a_381_47.t0 95.021
R212 a_381_47.n0 a_381_47.t3 63.333
R213 a_381_47.t1 a_381_47.n1 31.613
R214 a_381_47.n0 a_381_47.t2 26.77
R215 a_1056_47.t0 a_1056_47.t1 60
R216 D.n0 D.t0 264.028
R217 D.n0 D.t1 174.054
R218 D.n1 D.n0 76
R219 D.n1 D 8.585
R220 D D.n1 2.029
R221 SET_B.n0 SET_B.t0 401.403
R222 SET_B.n1 SET_B.t2 372.146
R223 SET_B.n1 SET_B.t3 148.348
R224 SET_B.n0 SET_B.t1 141.967
R225 SET_B.n2 SET_B.n1 97.332
R226 SET_B.n2 SET_B.n0 6.974
R227 SET_B SET_B.n2 3.246
R228 a_1602_47.n1 a_1602_47.t4 212.079
R229 a_1602_47.n0 a_1602_47.t2 212.079
R230 a_1602_47.n2 a_1602_47.t1 155.491
R231 a_1602_47.t0 a_1602_47.n2 149.578
R232 a_1602_47.n1 a_1602_47.t5 139.779
R233 a_1602_47.n0 a_1602_47.t3 139.779
R234 a_1602_47.n2 a_1602_47.n1 98.884
R235 a_1602_47.n1 a_1602_47.n0 61.345
R236 Q.n6 Q.n5 292.5
R237 Q.n5 Q.n4 147.104
R238 Q.n2 Q.n0 93.852
R239 Q.n3 Q.n2 39.863
R240 Q.n7 Q.n6 33.745
R241 Q.n5 Q.t1 26.595
R242 Q.n5 Q.t0 26.595
R243 Q.n0 Q.t3 24.923
R244 Q.n0 Q.t2 24.923
R245 Q.n1 Q 13.552
R246 Q.n8 Q 12.8
R247 Q.n4 Q 10.71
R248 Q.n3 Q 9.244
R249 Q Q.n8 7.841
R250 Q.n7 Q 7.466
R251 Q.n1 Q 7.2
R252 Q.n2 Q.n1 6.698
R253 Q.n8 Q.n7 5.12
R254 Q.n6 Q 4.848
R255 Q.n9 Q 4.843
R256 Q Q.n9 2.998
R257 Q.n4 Q 2.439
R258 Q.n3 Q 1.969
R259 Q.n9 Q.n3 0.875
R260 a_562_413.t0 a_562_413.t1 211.071
R261 a_1178_261.n0 a_1178_261.t3 387.607
R262 a_1178_261.t0 a_1178_261.n1 223.706
R263 a_1178_261.n1 a_1178_261.t1 202.187
R264 a_1178_261.n1 a_1178_261.n0 189.773
R265 a_1178_261.n0 a_1178_261.t2 169.453
R266 a_796_47.t0 a_796_47.t1 60
R267 a_1300_47.t0 a_1300_47.t1 60
C0 VPB VPWR 0.20fF
C1 VGND Q 0.21fF
C2 VPWR Q 0.36fF
C3 VPWR VGND 0.11fF
C4 SET_B VGND 0.48fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__dfstp_4.ext - technology: sky130A

.subckt sky130_fd_sc_hd__dfstp_4 Q D VPWR SET_B CLK VGND VNB VPB
X0 a_1178_261.t0 a_1028_413.t5 VPWR.t15 VPB.t19 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X1 VGND.t10 a_652_21.t3 a_586_47.t1 VNB.t10 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 VPWR.t14 a_1028_413.t6 a_1598_47.t0 VPB.t18 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X3 a_1178_261.t1 a_1028_413.t7 VGND.t12 VNB.t15 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=540000u l=150000u
X4 VGND.t4 a_1598_47.t2 Q.t9 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 a_956_413.t0 a_476_47.t4 VPWR.t5 VPB.t7 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 a_1136_413.t1 a_193_47.t2 a_1028_413.t0 VPB.t5 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7 VPWR.t4 a_1598_47.t3 Q.t4 VPB.t6 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 VPWR.t6 a_476_47.t5 a_652_21.t0 VPB.t8 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9 a_586_47.t0 a_193_47.t3 a_476_47.t0 VNB.t5 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X10 VGND.t0 a_1598_47.t4 Q.t8 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 VPWR.t11 CLK.t0 a_27_47.t0 VPB.t14 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X12 Q.t7 a_1598_47.t5 VGND.t1 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 a_476_47.t2 a_27_47.t2 a_381_47.t3 VNB.t11 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X14 a_1056_47.t1 a_476_47.t6 VGND.t5 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15 a_381_47.t1 D.t0 VPWR.t7 VPB.t9 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X16 a_652_21.t2 SET_B.t0 VPWR.t8 VPB.t11 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17 a_1224_47.t1 a_27_47.t3 a_1028_413.t3 VNB.t12 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18 a_562_413.t1 a_27_47.t4 a_476_47.t3 VPB.t15 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19 a_1028_413.t1 a_193_47.t4 a_1056_47.t0 VNB.t6 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20 a_476_47.t1 a_193_47.t5 a_381_47.t0 VPB.t10 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21 Q.t3 a_1598_47.t6 VPWR.t0 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X22 a_1296_47.t0 a_1178_261.t2 a_1224_47.t0 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23 VGND.t13 a_1028_413.t8 a_1598_47.t1 VNB.t14 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24 a_193_47.t0 a_27_47.t5 VGND.t11 VNB.t13 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X25 VPWR.t10 a_652_21.t4 a_562_413.t0 VPB.t13 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X26 VPWR.t1 a_1598_47.t7 Q.t2 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X27 VGND.t7 SET_B.t1 a_1296_47.t1 VNB.t7 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X28 Q.t1 a_1598_47.t8 VPWR.t2 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X29 a_1028_413.t4 a_27_47.t6 a_956_413.t1 VPB.t16 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X30 VPWR.t12 a_1178_261.t3 a_1136_413.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X31 a_193_47.t1 a_27_47.t7 VPWR.t13 VPB.t17 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X32 Q.t0 a_1598_47.t9 VPWR.t3 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X33 a_796_47.t1 SET_B.t2 VGND.t8 VNB.t8 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X34 a_381_47.t2 D.t1 VGND.t6 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X35 Q.t6 a_1598_47.t10 VGND.t2 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X36 Q.t5 a_1598_47.t11 VGND.t3 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X37 a_652_21.t1 a_476_47.t7 a_796_47.t0 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X38 VPWR.t9 SET_B.t3 a_1028_413.t2 VPB.t12 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X39 VGND.t9 CLK.t1 a_27_47.t1 VNB.t9 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
R0 a_1028_413.n4 a_1028_413.t2 433.656
R1 a_1028_413.n5 a_1028_413.n4 317.979
R2 a_1028_413.n1 a_1028_413.t6 237.786
R3 a_1028_413.n1 a_1028_413.t8 208.866
R4 a_1028_413.n2 a_1028_413.t5 205.653
R5 a_1028_413.n3 a_1028_413.n0 194.899
R6 a_1028_413.n2 a_1028_413.t7 189.586
R7 a_1028_413.n3 a_1028_413.n2 152.207
R8 a_1028_413.n2 a_1028_413.n1 137.296
R9 a_1028_413.t0 a_1028_413.n5 119.607
R10 a_1028_413.n4 a_1028_413.n3 94.87
R11 a_1028_413.n5 a_1028_413.t4 63.321
R12 a_1028_413.n0 a_1028_413.t3 47.142
R13 a_1028_413.n0 a_1028_413.t1 47.142
R14 VPWR.n42 VPWR.t7 429.335
R15 VPWR.n18 VPWR.t12 355.821
R16 VPWR.n1 VPWR.n0 320.609
R17 VPWR.n14 VPWR.n13 312.281
R18 VPWR.n47 VPWR.n46 311.893
R19 VPWR.n28 VPWR.n27 307.239
R20 VPWR.n33 VPWR.n32 292.5
R21 VPWR.n7 VPWR.n6 167.037
R22 VPWR.n3 VPWR.n2 166.889
R23 VPWR.n32 VPWR.t8 91.464
R24 VPWR.n13 VPWR.t9 91.464
R25 VPWR.n32 VPWR.t10 86.773
R26 VPWR.n27 VPWR.t5 63.321
R27 VPWR.n27 VPWR.t6 63.321
R28 VPWR.n6 VPWR.t14 58.484
R29 VPWR.n46 VPWR.t13 41.554
R30 VPWR.n46 VPWR.t11 41.554
R31 VPWR.n13 VPWR.t15 32.833
R32 VPWR.n6 VPWR.t2 31.605
R33 VPWR.n2 VPWR.t3 26.595
R34 VPWR.n2 VPWR.t4 26.595
R35 VPWR.n0 VPWR.t0 26.595
R36 VPWR.n0 VPWR.t1 26.595
R37 VPWR.n5 VPWR.n4 4.65
R38 VPWR.n8 VPWR.n7 4.65
R39 VPWR.n10 VPWR.n9 4.65
R40 VPWR.n12 VPWR.n11 4.65
R41 VPWR.n15 VPWR.n14 4.65
R42 VPWR.n17 VPWR.n16 4.65
R43 VPWR.n20 VPWR.n19 4.65
R44 VPWR.n22 VPWR.n21 4.65
R45 VPWR.n24 VPWR.n23 4.65
R46 VPWR.n26 VPWR.n25 4.65
R47 VPWR.n29 VPWR.n28 4.65
R48 VPWR.n31 VPWR.n30 4.65
R49 VPWR.n35 VPWR.n34 4.65
R50 VPWR.n37 VPWR.n36 4.65
R51 VPWR.n39 VPWR.n38 4.65
R52 VPWR.n41 VPWR.n40 4.65
R53 VPWR.n43 VPWR.n42 4.65
R54 VPWR.n45 VPWR.n44 4.65
R55 VPWR.n48 VPWR.n47 3.932
R56 VPWR.n3 VPWR.n1 3.812
R57 VPWR.n34 VPWR.n33 3.374
R58 VPWR.n19 VPWR.n18 0.814
R59 VPWR.n5 VPWR.n3 0.255
R60 VPWR.n48 VPWR.n45 0.137
R61 VPWR VPWR.n48 0.123
R62 VPWR.n8 VPWR.n5 0.119
R63 VPWR.n10 VPWR.n8 0.119
R64 VPWR.n12 VPWR.n10 0.119
R65 VPWR.n15 VPWR.n12 0.119
R66 VPWR.n17 VPWR.n15 0.119
R67 VPWR.n20 VPWR.n17 0.119
R68 VPWR.n22 VPWR.n20 0.119
R69 VPWR.n24 VPWR.n22 0.119
R70 VPWR.n26 VPWR.n24 0.119
R71 VPWR.n29 VPWR.n26 0.119
R72 VPWR.n31 VPWR.n29 0.119
R73 VPWR.n35 VPWR.n31 0.119
R74 VPWR.n37 VPWR.n35 0.119
R75 VPWR.n39 VPWR.n37 0.119
R76 VPWR.n41 VPWR.n39 0.119
R77 VPWR.n43 VPWR.n41 0.119
R78 VPWR.n45 VPWR.n43 0.119
R79 a_1178_261.n0 a_1178_261.t2 381.181
R80 a_1178_261.t0 a_1178_261.n1 224.916
R81 a_1178_261.n1 a_1178_261.t1 193.368
R82 a_1178_261.n1 a_1178_261.n0 189.773
R83 a_1178_261.n0 a_1178_261.t3 169.453
R84 VPB.t19 VPB.t18 556.386
R85 VPB.t0 VPB.t12 556.386
R86 VPB.t17 VPB.t9 556.386
R87 VPB.t15 VPB.t13 355.14
R88 VPB.t16 VPB.t5 319.626
R89 VPB.t13 VPB.t11 313.707
R90 VPB.t9 VPB.t10 287.071
R91 VPB.t12 VPB.t19 284.112
R92 VPB.t18 VPB.t3 281.152
R93 VPB.t6 VPB.t4 248.598
R94 VPB.t1 VPB.t6 248.598
R95 VPB.t2 VPB.t1 248.598
R96 VPB.t3 VPB.t2 248.598
R97 VPB.t8 VPB.t7 248.598
R98 VPB.t11 VPB.t8 248.598
R99 VPB.t10 VPB.t15 248.598
R100 VPB.t14 VPB.t17 248.598
R101 VPB.t5 VPB.t0 213.084
R102 VPB.t7 VPB.t16 213.084
R103 VPB VPB.t14 142.056
R104 a_652_21.n0 a_652_21.t3 387.959
R105 a_652_21.n2 a_652_21.n1 301.911
R106 a_652_21.n1 a_652_21.t1 241.655
R107 a_652_21.n0 a_652_21.t4 143.746
R108 a_652_21.n1 a_652_21.n0 111.072
R109 a_652_21.t0 a_652_21.n2 63.321
R110 a_652_21.n2 a_652_21.t2 63.321
R111 a_586_47.t1 a_586_47.t0 93.516
R112 VGND.n41 VGND.t6 188.008
R113 VGND.n25 VGND.t5 145.376
R114 VGND.n2 VGND.n1 111.574
R115 VGND.n3 VGND.n0 110.69
R116 VGND.n7 VGND.n6 109.566
R117 VGND.n46 VGND.n45 107.239
R118 VGND.n14 VGND.n13 92.5
R119 VGND.n30 VGND.n29 92.5
R120 VGND.n29 VGND.t10 81.428
R121 VGND.n13 VGND.t7 67.142
R122 VGND.n13 VGND.t12 55.301
R123 VGND.n6 VGND.t13 54.285
R124 VGND.n29 VGND.t8 38.571
R125 VGND.n45 VGND.t11 38.571
R126 VGND.n45 VGND.t9 38.571
R127 VGND.n6 VGND.t2 25.934
R128 VGND.n0 VGND.t1 24.923
R129 VGND.n0 VGND.t0 24.923
R130 VGND.n1 VGND.t3 24.923
R131 VGND.n1 VGND.t4 24.923
R132 VGND.n5 VGND.n4 4.65
R133 VGND.n8 VGND.n7 4.65
R134 VGND.n10 VGND.n9 4.65
R135 VGND.n12 VGND.n11 4.65
R136 VGND.n16 VGND.n15 4.65
R137 VGND.n18 VGND.n17 4.65
R138 VGND.n20 VGND.n19 4.65
R139 VGND.n22 VGND.n21 4.65
R140 VGND.n24 VGND.n23 4.65
R141 VGND.n26 VGND.n25 4.65
R142 VGND.n28 VGND.n27 4.65
R143 VGND.n32 VGND.n31 4.65
R144 VGND.n34 VGND.n33 4.65
R145 VGND.n36 VGND.n35 4.65
R146 VGND.n38 VGND.n37 4.65
R147 VGND.n40 VGND.n39 4.65
R148 VGND.n42 VGND.n41 4.65
R149 VGND.n44 VGND.n43 4.65
R150 VGND.n31 VGND.n30 4.511
R151 VGND.n47 VGND.n46 3.932
R152 VGND.n3 VGND.n2 3.812
R153 VGND.n15 VGND.n14 1.083
R154 VGND.n5 VGND.n3 0.255
R155 VGND.n47 VGND.n44 0.137
R156 VGND VGND.n47 0.123
R157 VGND.n8 VGND.n5 0.119
R158 VGND.n10 VGND.n8 0.119
R159 VGND.n12 VGND.n10 0.119
R160 VGND.n16 VGND.n12 0.119
R161 VGND.n18 VGND.n16 0.119
R162 VGND.n20 VGND.n18 0.119
R163 VGND.n22 VGND.n20 0.119
R164 VGND.n24 VGND.n22 0.119
R165 VGND.n26 VGND.n24 0.119
R166 VGND.n28 VGND.n26 0.119
R167 VGND.n32 VGND.n28 0.119
R168 VGND.n34 VGND.n32 0.119
R169 VGND.n36 VGND.n34 0.119
R170 VGND.n38 VGND.n36 0.119
R171 VGND.n40 VGND.n38 0.119
R172 VGND.n42 VGND.n40 0.119
R173 VGND.n44 VGND.n42 0.119
R174 VNB.t3 VNB.t2 6082.35
R175 VNB.t13 VNB.t4 5346.86
R176 VNB.t15 VNB.t14 5170
R177 VNB VNB.t9 4270.59
R178 VNB.t10 VNB.t8 3688.24
R179 VNB.t7 VNB.t15 3570.15
R180 VNB.t11 VNB.t5 3558.82
R181 VNB.t6 VNB.t12 3105.88
R182 VNB.t5 VNB.t10 3105.88
R183 VNB.t9 VNB.t13 2717.65
R184 VNB.t0 VNB.t7 2329.41
R185 VNB.t12 VNB.t0 2329.41
R186 VNB.t2 VNB.t6 2329.41
R187 VNB.t8 VNB.t3 2329.41
R188 VNB.t4 VNB.t11 2280.14
R189 VNB.t14 VNB.t1 145.876
R190 a_1598_47.t0 a_1598_47.n14 255.522
R191 a_1598_47.n0 a_1598_47.t9 221.719
R192 a_1598_47.n2 a_1598_47.t3 221.719
R193 a_1598_47.n5 a_1598_47.t6 221.719
R194 a_1598_47.n8 a_1598_47.t7 221.719
R195 a_1598_47.n11 a_1598_47.t8 221.719
R196 a_1598_47.n14 a_1598_47.t1 164.607
R197 a_1598_47.n0 a_1598_47.t5 149.419
R198 a_1598_47.n2 a_1598_47.t4 149.419
R199 a_1598_47.n5 a_1598_47.t11 149.419
R200 a_1598_47.n8 a_1598_47.t2 149.419
R201 a_1598_47.n11 a_1598_47.t10 149.419
R202 a_1598_47.n4 a_1598_47.n1 95.781
R203 a_1598_47.n13 a_1598_47.n12 76
R204 a_1598_47.n4 a_1598_47.n3 76
R205 a_1598_47.n7 a_1598_47.n6 76
R206 a_1598_47.n10 a_1598_47.n9 76
R207 a_1598_47.n1 a_1598_47.n0 41.059
R208 a_1598_47.n14 a_1598_47.n13 35.49
R209 a_1598_47.n3 a_1598_47.n2 26.777
R210 a_1598_47.n7 a_1598_47.n4 19.781
R211 a_1598_47.n10 a_1598_47.n7 19.781
R212 a_1598_47.n13 a_1598_47.n10 19.781
R213 a_1598_47.n12 a_1598_47.n11 16.066
R214 a_1598_47.n6 a_1598_47.n5 12.496
R215 a_1598_47.n9 a_1598_47.n8 1.785
R216 Q.n10 Q.t0 208.199
R217 Q.n9 Q.n6 165.935
R218 Q.n8 Q.n7 142.828
R219 Q.n4 Q.t7 117.423
R220 Q.n3 Q.n0 98.9
R221 Q.n2 Q.n1 92.5
R222 Q.n9 Q 63.216
R223 Q.n3 Q.n2 60.081
R224 Q.n11 Q.n9 56.847
R225 Q.n5 Q.n3 56.847
R226 Q.n7 Q.t2 26.595
R227 Q.n7 Q.t1 26.595
R228 Q.n6 Q.t4 26.595
R229 Q.n6 Q.t3 26.595
R230 Q.n1 Q.t9 24.923
R231 Q.n1 Q.t6 24.923
R232 Q.n0 Q.t8 24.923
R233 Q.n0 Q.t5 24.923
R234 Q.n13 Q 12.243
R235 Q.n2 Q 10.71
R236 Q Q.n8 9.561
R237 Q.n11 Q 8.411
R238 Q.n8 Q 7.781
R239 Q.n4 Q 7.497
R240 Q Q.n10 6.727
R241 Q Q.n13 6.678
R242 Q.n10 Q 5.563
R243 Q Q.n4 4.937
R244 Q.n12 Q.n11 3.108
R245 Q.n13 Q.n5 3.108
R246 Q Q.n12 1.391
R247 Q.n5 Q 1.28
R248 Q.n12 Q 0.914
R249 a_476_47.n4 a_476_47.n3 415.031
R250 a_476_47.n1 a_476_47.t6 344.897
R251 a_476_47.n2 a_476_47.t4 289.491
R252 a_476_47.n2 a_476_47.t5 228.146
R253 a_476_47.n3 a_476_47.n0 196.424
R254 a_476_47.n3 a_476_47.n2 138.78
R255 a_476_47.n2 a_476_47.n1 105.747
R256 a_476_47.n1 a_476_47.t7 93.186
R257 a_476_47.n0 a_476_47.t2 70
R258 a_476_47.n0 a_476_47.t0 63.333
R259 a_476_47.n4 a_476_47.t3 63.321
R260 a_476_47.t1 a_476_47.n4 63.321
R261 a_956_413.t0 a_956_413.t1 98.5
R262 a_193_47.n1 a_193_47.t5 538.583
R263 a_193_47.n0 a_193_47.t2 373.664
R264 a_193_47.t1 a_193_47.n3 278.596
R265 a_193_47.n0 a_193_47.t4 264.028
R266 a_193_47.n3 a_193_47.t0 150.413
R267 a_193_47.n1 a_193_47.t3 135.794
R268 a_193_47.n2 a_193_47.n0 27.501
R269 a_193_47.n2 a_193_47.n1 10.05
R270 a_193_47.n3 a_193_47.n2 6.187
R271 a_1136_413.t0 a_1136_413.t1 98.5
R272 CLK.n0 CLK.t0 270.454
R273 CLK.n0 CLK.t1 235.108
R274 CLK.n1 CLK.n0 76
R275 CLK.n1 CLK 7.68
R276 CLK CLK.n1 4.754
R277 a_27_47.n0 a_27_47.t3 346.686
R278 a_27_47.n3 a_27_47.t7 263.171
R279 a_27_47.t0 a_27_47.n5 243.779
R280 a_27_47.n1 a_27_47.t2 235.952
R281 a_27_47.n1 a_27_47.t4 232.166
R282 a_27_47.n3 a_27_47.t5 227.825
R283 a_27_47.n4 a_27_47.t1 195.494
R284 a_27_47.n0 a_27_47.t6 158.045
R285 a_27_47.n4 a_27_47.n3 76
R286 a_27_47.n5 a_27_47.n4 35.339
R287 a_27_47.n2 a_27_47.n0 6.892
R288 a_27_47.n5 a_27_47.n2 6.181
R289 a_27_47.n2 a_27_47.n1 4.65
R290 a_381_47.n1 a_381_47.n0 405.201
R291 a_381_47.n1 a_381_47.t0 95.021
R292 a_381_47.n0 a_381_47.t3 63.333
R293 a_381_47.t1 a_381_47.n1 31.613
R294 a_381_47.n0 a_381_47.t2 26.77
R295 a_1056_47.t0 a_1056_47.t1 60
R296 D.n0 D.t0 264.028
R297 D.n0 D.t1 174.054
R298 D.n1 D.n0 76
R299 D.n1 D 8.585
R300 D D.n1 2.029
R301 SET_B.n0 SET_B.t0 401.403
R302 SET_B.n1 SET_B.t3 386.89
R303 SET_B.n1 SET_B.t1 148.348
R304 SET_B.n0 SET_B.t2 141.967
R305 SET_B.n2 SET_B.n1 98.281
R306 SET_B.n2 SET_B.n0 6.974
R307 SET_B SET_B.n2 3.246
R308 a_1224_47.t0 a_1224_47.t1 60
R309 a_562_413.t0 a_562_413.t1 211.071
R310 a_1296_47.t0 a_1296_47.t1 60
R311 a_796_47.t0 a_796_47.t1 60
C0 VPB VPWR 0.22fF
C1 VGND Q 0.48fF
C2 VPWR Q 0.74fF
C3 VPWR VGND 0.14fF
C4 SET_B VGND 0.48fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__dfxbp_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__dfxbp_1 VGND VPWR Q_N D CLK Q VNB VPB
X0 Q.t1 a_1059_315.t2 VGND.t1 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 a_891_413.t2 a_193_47.t2 a_634_159.t3 VNB.t12 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X2 a_561_413.t0 a_27_47.t2 a_466_413.t0 VPB.t5 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3 VPWR.t4 CLK.t0 a_27_47.t0 VPB.t9 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X4 a_381_47.t2 D.t0 VPWR.t8 VPB.t10 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 VGND.t4 a_634_159.t4 a_592_47.t0 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 a_466_413.t3 a_193_47.t3 a_381_47.t1 VPB.t13 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7 VPWR.t7 a_634_159.t5 a_561_413.t1 VPB.t8 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 a_634_159.t1 a_466_413.t4 VGND.t9 VNB.t11 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X9 Q.t0 a_1059_315.t3 VPWR.t2 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 VGND.t3 a_1059_315.t4 a_1490_369.t1 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11 a_634_159.t2 a_466_413.t5 VPWR.t5 VPB.t6 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X12 a_975_413.t1 a_193_47.t4 a_891_413.t3 VPB.t12 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13 VGND.t2 a_1059_315.t5 a_1017_47.t0 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14 a_193_47.t0 a_27_47.t3 VGND.t5 VNB.t5 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15 a_891_413.t0 a_27_47.t4 a_634_159.t0 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16 a_592_47.t1 a_193_47.t5 a_466_413.t2 VNB.t13 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X17 VPWR.t9 a_891_413.t4 a_1059_315.t0 VPB.t11 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X18 a_1017_47.t1 a_27_47.t5 a_891_413.t1 VNB.t6 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X19 VPWR.t1 a_1059_315.t6 a_975_413.t0 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20 a_466_413.t1 a_27_47.t6 a_381_47.t0 VNB.t7 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X21 a_193_47.t1 a_27_47.t7 VPWR.t3 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X22 VGND.t0 a_891_413.t5 a_1059_315.t1 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X23 Q_N.t1 a_1490_369.t2 VGND.t8 VNB.t10 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X24 a_381_47.t3 D.t1 VGND.t7 VNB.t9 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X25 Q_N.t0 a_1490_369.t3 VPWR.t6 VPB.t7 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X26 VGND.t6 CLK.t1 a_27_47.t1 VNB.t8 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X27 VPWR.t0 a_1059_315.t7 a_1490_369.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
R0 a_1059_315.n3 a_1059_315.t5 382.743
R1 a_1059_315.n0 a_1059_315.t7 258.795
R2 a_1059_315.n1 a_1059_315.t3 213.539
R3 a_1059_315.n0 a_1059_315.t4 166.387
R4 a_1059_315.n1 a_1059_315.t2 139.779
R5 a_1059_315.n3 a_1059_315.t6 138.53
R6 a_1059_315.n1 a_1059_315.n0 129.263
R7 a_1059_315.t0 a_1059_315.n4 128.779
R8 a_1059_315.n2 a_1059_315.t1 103.313
R9 a_1059_315.n4 a_1059_315.n3 97.957
R10 a_1059_315.n2 a_1059_315.n1 97.915
R11 a_1059_315.n4 a_1059_315.n2 16.622
R12 VGND.n6 VGND.t2 158.499
R13 VGND.n25 VGND.t7 150.527
R14 VGND.n2 VGND.n1 126.005
R15 VGND.n3 VGND.n0 111.467
R16 VGND.n30 VGND.n29 107.239
R17 VGND.n17 VGND.n16 107.029
R18 VGND.n16 VGND.t9 74.865
R19 VGND.n0 VGND.t3 54.285
R20 VGND.n16 VGND.t4 40
R21 VGND.n29 VGND.t5 38.571
R22 VGND.n29 VGND.t6 38.571
R23 VGND.n0 VGND.t8 25.934
R24 VGND.n1 VGND.t1 24.923
R25 VGND.n1 VGND.t0 24.923
R26 VGND.n3 VGND.n2 6.015
R27 VGND.n5 VGND.n4 4.65
R28 VGND.n7 VGND.n6 4.65
R29 VGND.n9 VGND.n8 4.65
R30 VGND.n11 VGND.n10 4.65
R31 VGND.n13 VGND.n12 4.65
R32 VGND.n15 VGND.n14 4.65
R33 VGND.n18 VGND.n17 4.65
R34 VGND.n20 VGND.n19 4.65
R35 VGND.n22 VGND.n21 4.65
R36 VGND.n24 VGND.n23 4.65
R37 VGND.n26 VGND.n25 4.65
R38 VGND.n28 VGND.n27 4.65
R39 VGND.n31 VGND.n30 3.932
R40 VGND.n5 VGND.n3 0.14
R41 VGND.n31 VGND.n28 0.137
R42 VGND VGND.n31 0.123
R43 VGND.n7 VGND.n5 0.119
R44 VGND.n9 VGND.n7 0.119
R45 VGND.n11 VGND.n9 0.119
R46 VGND.n13 VGND.n11 0.119
R47 VGND.n15 VGND.n13 0.119
R48 VGND.n18 VGND.n15 0.119
R49 VGND.n20 VGND.n18 0.119
R50 VGND.n22 VGND.n20 0.119
R51 VGND.n24 VGND.n22 0.119
R52 VGND.n26 VGND.n24 0.119
R53 VGND.n28 VGND.n26 0.119
R54 Q.n0 Q.t0 219.77
R55 Q.n0 Q.t1 82.859
R56 Q Q.n0 5.75
R57 VNB.t5 VNB.t9 6082.35
R58 VNB.t1 VNB.t0 5386.59
R59 VNB.t3 VNB.t2 4545.05
R60 VNB VNB.t8 4270.59
R61 VNB.t9 VNB.t7 3623.53
R62 VNB.t12 VNB.t6 3429.41
R63 VNB.t13 VNB.t4 3202.94
R64 VNB.t7 VNB.t13 3202.94
R65 VNB.t4 VNB.t11 3130.33
R66 VNB.t6 VNB.t1 3073.53
R67 VNB.t8 VNB.t5 2717.65
R68 VNB.t11 VNB.t12 2363.68
R69 VNB.t2 VNB.t10 2296.7
R70 VNB.t0 VNB.t3 2030.77
R71 a_193_47.n1 a_193_47.t5 407.215
R72 a_193_47.n1 a_193_47.t3 273.571
R73 a_193_47.t1 a_193_47.n3 246.213
R74 a_193_47.n0 a_193_47.t4 232.651
R75 a_193_47.n0 a_193_47.t2 222.372
R76 a_193_47.n3 a_193_47.t0 201.643
R77 a_193_47.n2 a_193_47.n1 90.25
R78 a_193_47.n2 a_193_47.n0 6.797
R79 a_193_47.n3 a_193_47.n2 5.609
R80 a_634_159.n1 a_634_159.t5 406.399
R81 a_634_159.n3 a_634_159.n2 381.512
R82 a_634_159.n1 a_634_159.t4 130.052
R83 a_634_159.n2 a_634_159.n0 121.487
R84 a_634_159.n2 a_634_159.n1 104.16
R85 a_634_159.n3 a_634_159.t0 89.119
R86 a_634_159.n0 a_634_159.t3 71.666
R87 a_634_159.t2 a_634_159.n3 37.523
R88 a_634_159.n0 a_634_159.t1 28.437
R89 a_891_413.n3 a_891_413.n2 403.558
R90 a_891_413.n1 a_891_413.t4 212.079
R91 a_891_413.n2 a_891_413.n1 175.108
R92 a_891_413.n2 a_891_413.n0 166.287
R93 a_891_413.n1 a_891_413.t5 141.239
R94 a_891_413.n0 a_891_413.t1 76.666
R95 a_891_413.n3 a_891_413.t3 63.321
R96 a_891_413.t0 a_891_413.n3 63.321
R97 a_891_413.n0 a_891_413.t2 50
R98 a_27_47.n2 a_27_47.t5 443.438
R99 a_27_47.n3 a_27_47.t6 270.054
R100 a_27_47.n4 a_27_47.t7 263.171
R101 a_27_47.n2 a_27_47.t4 254.388
R102 a_27_47.t0 a_27_47.n6 243.779
R103 a_27_47.n4 a_27_47.t3 227.825
R104 a_27_47.n5 a_27_47.t1 195.494
R105 a_27_47.n0 a_27_47.t2 142.671
R106 a_27_47.n1 a_27_47.n2 112.935
R107 a_27_47.n5 a_27_47.n4 76
R108 a_27_47.n6 a_27_47.n5 35.339
R109 a_27_47.n6 a_27_47.n1 6.379
R110 a_27_47.n1 a_27_47.n0 4.695
R111 a_27_47.n0 a_27_47.n3 2.98
R112 a_466_413.n3 a_466_413.n2 403.181
R113 a_466_413.n0 a_466_413.t4 230.482
R114 a_466_413.n2 a_466_413.n1 205.859
R115 a_466_413.n0 a_466_413.t5 196.013
R116 a_466_413.n2 a_466_413.n0 92.738
R117 a_466_413.n3 a_466_413.t3 79.738
R118 a_466_413.t0 a_466_413.n3 72.702
R119 a_466_413.n1 a_466_413.t2 70
R120 a_466_413.n1 a_466_413.t1 45
R121 a_561_413.t0 a_561_413.t1 171.202
R122 VPB.t1 VPB.t11 624.454
R123 VPB.t2 VPB.t0 556.386
R124 VPB.t3 VPB.t10 556.386
R125 VPB.t8 VPB.t6 390.654
R126 VPB.t12 VPB.t1 337.383
R127 VPB.t5 VPB.t8 304.828
R128 VPB.t0 VPB.t7 287.071
R129 VPB.t6 VPB.t4 281.152
R130 VPB.t13 VPB.t5 281.152
R131 VPB.t10 VPB.t13 251.557
R132 VPB.t11 VPB.t2 248.598
R133 VPB.t4 VPB.t12 248.598
R134 VPB.t9 VPB.t3 248.598
R135 VPB VPB.t9 142.056
R136 CLK.n0 CLK.t0 294.554
R137 CLK.n0 CLK.t1 211.008
R138 CLK CLK.n0 77.969
R139 VPWR.n6 VPWR.t1 375.232
R140 VPWR.n26 VPWR.t8 374.175
R141 VPWR.n31 VPWR.n30 311.893
R142 VPWR.n1 VPWR.n0 186.917
R143 VPWR.n15 VPWR.n14 174.594
R144 VPWR.n3 VPWR.n2 144.296
R145 VPWR.n14 VPWR.t7 113.978
R146 VPWR.n2 VPWR.t0 61.922
R147 VPWR.n30 VPWR.t3 41.554
R148 VPWR.n30 VPWR.t4 41.554
R149 VPWR.n14 VPWR.t5 35.46
R150 VPWR.n2 VPWR.t6 30.231
R151 VPWR.n0 VPWR.t2 26.595
R152 VPWR.n0 VPWR.t9 26.595
R153 VPWR.n16 VPWR.n15 16.188
R154 VPWR.n3 VPWR.n1 6.769
R155 VPWR.n5 VPWR.n4 4.65
R156 VPWR.n7 VPWR.n6 4.65
R157 VPWR.n9 VPWR.n8 4.65
R158 VPWR.n11 VPWR.n10 4.65
R159 VPWR.n13 VPWR.n12 4.65
R160 VPWR.n17 VPWR.n16 4.65
R161 VPWR.n19 VPWR.n18 4.65
R162 VPWR.n21 VPWR.n20 4.65
R163 VPWR.n23 VPWR.n22 4.65
R164 VPWR.n25 VPWR.n24 4.65
R165 VPWR.n27 VPWR.n26 4.65
R166 VPWR.n29 VPWR.n28 4.65
R167 VPWR.n32 VPWR.n31 3.932
R168 VPWR.n5 VPWR.n3 0.14
R169 VPWR.n32 VPWR.n29 0.137
R170 VPWR VPWR.n32 0.123
R171 VPWR.n7 VPWR.n5 0.119
R172 VPWR.n9 VPWR.n7 0.119
R173 VPWR.n11 VPWR.n9 0.119
R174 VPWR.n13 VPWR.n11 0.119
R175 VPWR.n17 VPWR.n13 0.119
R176 VPWR.n19 VPWR.n17 0.119
R177 VPWR.n21 VPWR.n19 0.119
R178 VPWR.n23 VPWR.n21 0.119
R179 VPWR.n25 VPWR.n23 0.119
R180 VPWR.n27 VPWR.n25 0.119
R181 VPWR.n29 VPWR.n27 0.119
R182 D.n0 D.t1 302.729
R183 D.n0 D.t0 212.756
R184 D D.n0 94.057
R185 a_381_47.n1 a_381_47.n0 511.303
R186 a_381_47.n0 a_381_47.t0 90
R187 a_381_47.t1 a_381_47.n1 65.666
R188 a_381_47.n1 a_381_47.t2 63.321
R189 a_381_47.n0 a_381_47.t3 31.393
R190 a_592_47.t0 a_592_47.t1 99.726
R191 a_1490_369.t0 a_1490_369.n1 243.368
R192 a_1490_369.n0 a_1490_369.t3 236.932
R193 a_1490_369.n0 a_1490_369.t2 164.632
R194 a_1490_369.n1 a_1490_369.t1 162.124
R195 a_1490_369.n1 a_1490_369.n0 97.527
R196 a_975_413.t0 a_975_413.t1 197
R197 a_1017_47.t0 a_1017_47.t1 93.059
R198 Q_N Q_N.t1 167.063
R199 Q_N Q_N.t0 135.522
C0 VPWR VGND 0.12fF
C1 VPB VPWR 0.18fF
C2 Q VGND 0.11fF
C3 Q_N VPWR 0.17fF
C4 Q VPWR 0.16fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__dfxbp_2.ext - technology: sky130A

.subckt sky130_fd_sc_hd__dfxbp_2 VGND VPWR Q_N D CLK Q VNB VPB
X0 Q.t3 a_1059_315.t2 VGND.t5 VNB.t10 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 a_891_413.t3 a_193_47.t2 a_634_159.t3 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X2 a_561_413.t1 a_27_47.t2 a_466_413.t1 VPB.t12 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3 VPWR.t8 CLK.t0 a_27_47.t0 VPB.t13 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X4 a_381_47.t1 D.t0 VPWR.t10 VPB.t9 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 VGND.t3 a_1059_315.t3 a_1589_47.t0 VNB.t9 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 VGND.t9 a_634_159.t4 a_592_47.t0 VNB.t13 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7 VPWR.t0 a_1589_47.t2 Q_N.t3 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 VPWR.t6 a_1059_315.t4 Q.t1 VPB.t6 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 VGND.t0 a_1589_47.t3 Q_N.t1 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 a_466_413.t2 a_193_47.t3 a_381_47.t3 VPB.t15 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11 VPWR.t2 a_634_159.t5 a_561_413.t0 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12 a_634_159.t1 a_466_413.t4 VGND.t8 VNB.t12 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X13 Q.t0 a_1059_315.t5 VPWR.t5 VPB.t5 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14 a_634_159.t2 a_466_413.t5 VPWR.t9 VPB.t8 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X15 a_975_413.t1 a_193_47.t4 a_891_413.t2 VPB.t14 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16 Q_N.t2 a_1589_47.t4 VPWR.t1 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17 VGND.t6 a_1059_315.t6 a_1017_47.t0 VNB.t8 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18 a_193_47.t0 a_27_47.t3 VGND.t1 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19 a_891_413.t0 a_27_47.t4 a_634_159.t0 VPB.t11 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20 a_592_47.t1 a_193_47.t5 a_466_413.t3 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X21 VPWR.t7 a_891_413.t4 a_1059_315.t0 VPB.t7 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X22 VPWR.t3 a_1059_315.t7 a_1589_47.t1 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X23 Q_N.t0 a_1589_47.t5 VGND.t7 VNB.t11 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X24 a_1017_47.t1 a_27_47.t5 a_891_413.t1 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X25 VPWR.t4 a_1059_315.t8 a_975_413.t0 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X26 a_466_413.t0 a_27_47.t6 a_381_47.t2 VNB.t5 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X27 a_193_47.t1 a_27_47.t7 VPWR.t11 VPB.t10 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X28 VGND.t2 a_891_413.t5 a_1059_315.t1 VNB.t6 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X29 VGND.t4 a_1059_315.t9 Q.t2 VNB.t7 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X30 a_381_47.t0 D.t1 VGND.t10 VNB.t14 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X31 VGND.t11 CLK.t1 a_27_47.t1 VNB.t15 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
R0 a_1059_315.n5 a_1059_315.t6 382.743
R1 a_1059_315.n0 a_1059_315.t7 258.795
R2 a_1059_315.n3 a_1059_315.t5 213.539
R3 a_1059_315.n2 a_1059_315.t4 212.079
R4 a_1059_315.n0 a_1059_315.t3 167.834
R5 a_1059_315.n1 a_1059_315.n0 140.218
R6 a_1059_315.n3 a_1059_315.t2 139.779
R7 a_1059_315.n1 a_1059_315.t9 139.779
R8 a_1059_315.n5 a_1059_315.t8 138.53
R9 a_1059_315.t0 a_1059_315.n6 128.779
R10 a_1059_315.n4 a_1059_315.t1 103.313
R11 a_1059_315.n6 a_1059_315.n5 97.957
R12 a_1059_315.n4 a_1059_315.n3 97.915
R13 a_1059_315.n3 a_1059_315.n2 59.884
R14 a_1059_315.n6 a_1059_315.n4 16.622
R15 a_1059_315.n2 a_1059_315.n1 1.46
R16 VGND.n16 VGND.t6 158.499
R17 VGND.n35 VGND.t10 150.527
R18 VGND.n5 VGND.t4 143.775
R19 VGND.n11 VGND.n10 126.005
R20 VGND.n2 VGND.t0 114.941
R21 VGND.n40 VGND.n39 107.239
R22 VGND.n27 VGND.n26 107.029
R23 VGND.n26 VGND.t8 74.865
R24 VGND.n1 VGND.n0 64.44
R25 VGND.n0 VGND.t3 57.793
R26 VGND.n26 VGND.t9 40
R27 VGND.n39 VGND.t1 38.571
R28 VGND.n39 VGND.t11 38.571
R29 VGND.n10 VGND.t5 24.923
R30 VGND.n10 VGND.t2 24.923
R31 VGND.n0 VGND.t7 24.767
R32 VGND.n6 VGND.n5 7.905
R33 VGND.n4 VGND.n3 4.65
R34 VGND.n7 VGND.n6 4.65
R35 VGND.n9 VGND.n8 4.65
R36 VGND.n13 VGND.n12 4.65
R37 VGND.n15 VGND.n14 4.65
R38 VGND.n17 VGND.n16 4.65
R39 VGND.n19 VGND.n18 4.65
R40 VGND.n21 VGND.n20 4.65
R41 VGND.n23 VGND.n22 4.65
R42 VGND.n25 VGND.n24 4.65
R43 VGND.n28 VGND.n27 4.65
R44 VGND.n30 VGND.n29 4.65
R45 VGND.n32 VGND.n31 4.65
R46 VGND.n34 VGND.n33 4.65
R47 VGND.n36 VGND.n35 4.65
R48 VGND.n38 VGND.n37 4.65
R49 VGND.n41 VGND.n40 3.932
R50 VGND.n2 VGND.n1 3.742
R51 VGND.n12 VGND.n11 1.882
R52 VGND.n4 VGND.n2 0.245
R53 VGND.n41 VGND.n38 0.137
R54 VGND VGND.n41 0.123
R55 VGND.n7 VGND.n4 0.119
R56 VGND.n9 VGND.n7 0.119
R57 VGND.n13 VGND.n9 0.119
R58 VGND.n15 VGND.n13 0.119
R59 VGND.n17 VGND.n15 0.119
R60 VGND.n19 VGND.n17 0.119
R61 VGND.n21 VGND.n19 0.119
R62 VGND.n23 VGND.n21 0.119
R63 VGND.n25 VGND.n23 0.119
R64 VGND.n28 VGND.n25 0.119
R65 VGND.n30 VGND.n28 0.119
R66 VGND.n32 VGND.n30 0.119
R67 VGND.n34 VGND.n32 0.119
R68 VGND.n36 VGND.n34 0.119
R69 VGND.n38 VGND.n36 0.119
R70 Q.n1 Q.n0 187.307
R71 Q Q.n2 93.663
R72 Q.n0 Q.t1 26.595
R73 Q.n0 Q.t0 26.595
R74 Q.n2 Q.t2 24.923
R75 Q.n2 Q.t3 24.923
R76 Q Q.n1 12.024
R77 VNB.t3 VNB.t14 6082.35
R78 VNB.t8 VNB.t6 5386.59
R79 VNB.t7 VNB.t9 4859.34
R80 VNB VNB.t15 4270.59
R81 VNB.t14 VNB.t5 3623.53
R82 VNB.t0 VNB.t4 3429.41
R83 VNB.t1 VNB.t13 3202.94
R84 VNB.t5 VNB.t1 3202.94
R85 VNB.t13 VNB.t12 3130.33
R86 VNB.t4 VNB.t8 3073.53
R87 VNB.t15 VNB.t3 2717.65
R88 VNB.t12 VNB.t0 2363.68
R89 VNB.t9 VNB.t11 2345.05
R90 VNB.t11 VNB.t2 2030.77
R91 VNB.t10 VNB.t7 2030.77
R92 VNB.t6 VNB.t10 2030.77
R93 a_193_47.n1 a_193_47.t5 407.215
R94 a_193_47.n1 a_193_47.t3 273.571
R95 a_193_47.t1 a_193_47.n3 246.213
R96 a_193_47.n0 a_193_47.t4 232.651
R97 a_193_47.n0 a_193_47.t2 222.372
R98 a_193_47.n3 a_193_47.t0 201.643
R99 a_193_47.n2 a_193_47.n1 90.25
R100 a_193_47.n2 a_193_47.n0 6.797
R101 a_193_47.n3 a_193_47.n2 5.609
R102 a_634_159.n1 a_634_159.t5 406.399
R103 a_634_159.n3 a_634_159.n2 381.512
R104 a_634_159.n1 a_634_159.t4 130.052
R105 a_634_159.n2 a_634_159.n0 121.487
R106 a_634_159.n2 a_634_159.n1 104.16
R107 a_634_159.n3 a_634_159.t0 89.119
R108 a_634_159.n0 a_634_159.t3 71.666
R109 a_634_159.t2 a_634_159.n3 37.523
R110 a_634_159.n0 a_634_159.t1 28.437
R111 a_891_413.n3 a_891_413.n2 403.558
R112 a_891_413.n1 a_891_413.t4 212.079
R113 a_891_413.n2 a_891_413.n1 175.108
R114 a_891_413.n2 a_891_413.n0 166.287
R115 a_891_413.n1 a_891_413.t5 141.239
R116 a_891_413.n0 a_891_413.t1 76.666
R117 a_891_413.n3 a_891_413.t2 63.321
R118 a_891_413.t0 a_891_413.n3 63.321
R119 a_891_413.n0 a_891_413.t3 50
R120 a_27_47.n2 a_27_47.t5 443.438
R121 a_27_47.n3 a_27_47.t6 270.054
R122 a_27_47.n4 a_27_47.t7 263.171
R123 a_27_47.n2 a_27_47.t4 254.388
R124 a_27_47.t0 a_27_47.n6 243.779
R125 a_27_47.n4 a_27_47.t3 227.825
R126 a_27_47.n5 a_27_47.t1 195.494
R127 a_27_47.n0 a_27_47.t2 142.671
R128 a_27_47.n1 a_27_47.n2 112.935
R129 a_27_47.n5 a_27_47.n4 76
R130 a_27_47.n6 a_27_47.n5 35.339
R131 a_27_47.n6 a_27_47.n1 6.379
R132 a_27_47.n1 a_27_47.n0 4.695
R133 a_27_47.n0 a_27_47.n3 2.98
R134 a_466_413.n3 a_466_413.n2 403.181
R135 a_466_413.n0 a_466_413.t4 230.482
R136 a_466_413.n2 a_466_413.n1 205.859
R137 a_466_413.n0 a_466_413.t5 196.013
R138 a_466_413.n2 a_466_413.n0 92.738
R139 a_466_413.n3 a_466_413.t2 79.738
R140 a_466_413.t1 a_466_413.n3 72.702
R141 a_466_413.n1 a_466_413.t3 70
R142 a_466_413.n1 a_466_413.t0 45
R143 a_561_413.t0 a_561_413.t1 171.202
R144 VPB.t3 VPB.t7 624.454
R145 VPB.t6 VPB.t4 600.778
R146 VPB.t10 VPB.t9 556.386
R147 VPB.t2 VPB.t8 390.654
R148 VPB.t14 VPB.t3 337.383
R149 VPB.t12 VPB.t2 304.828
R150 VPB.t4 VPB.t1 287.071
R151 VPB.t8 VPB.t11 281.152
R152 VPB.t15 VPB.t12 281.152
R153 VPB.t9 VPB.t15 251.557
R154 VPB.t1 VPB.t0 248.598
R155 VPB.t5 VPB.t6 248.598
R156 VPB.t7 VPB.t5 248.598
R157 VPB.t11 VPB.t14 248.598
R158 VPB.t13 VPB.t10 248.598
R159 VPB VPB.t13 142.056
R160 CLK.n0 CLK.t0 294.554
R161 CLK.n0 CLK.t1 211.008
R162 CLK CLK.n0 77.969
R163 VPWR.n16 VPWR.t4 375.232
R164 VPWR.n36 VPWR.t10 374.175
R165 VPWR.n41 VPWR.n40 311.893
R166 VPWR.n5 VPWR.t6 215.014
R167 VPWR.n11 VPWR.n10 186.917
R168 VPWR.n25 VPWR.n24 174.594
R169 VPWR.n2 VPWR.t0 157.829
R170 VPWR.n1 VPWR.n0 140.41
R171 VPWR.n24 VPWR.t2 113.978
R172 VPWR.n0 VPWR.t3 61.922
R173 VPWR.n40 VPWR.t11 41.554
R174 VPWR.n40 VPWR.t8 41.554
R175 VPWR.n24 VPWR.t9 35.46
R176 VPWR.n0 VPWR.t1 30.231
R177 VPWR.n10 VPWR.t5 26.595
R178 VPWR.n10 VPWR.t7 26.595
R179 VPWR.n26 VPWR.n25 16.188
R180 VPWR.n4 VPWR.n3 4.65
R181 VPWR.n7 VPWR.n6 4.65
R182 VPWR.n9 VPWR.n8 4.65
R183 VPWR.n13 VPWR.n12 4.65
R184 VPWR.n15 VPWR.n14 4.65
R185 VPWR.n17 VPWR.n16 4.65
R186 VPWR.n19 VPWR.n18 4.65
R187 VPWR.n21 VPWR.n20 4.65
R188 VPWR.n23 VPWR.n22 4.65
R189 VPWR.n27 VPWR.n26 4.65
R190 VPWR.n29 VPWR.n28 4.65
R191 VPWR.n31 VPWR.n30 4.65
R192 VPWR.n33 VPWR.n32 4.65
R193 VPWR.n35 VPWR.n34 4.65
R194 VPWR.n37 VPWR.n36 4.65
R195 VPWR.n39 VPWR.n38 4.65
R196 VPWR.n42 VPWR.n41 3.932
R197 VPWR.n2 VPWR.n1 3.905
R198 VPWR.n12 VPWR.n11 2.635
R199 VPWR.n6 VPWR.n5 1.882
R200 VPWR.n4 VPWR.n2 0.223
R201 VPWR.n42 VPWR.n39 0.137
R202 VPWR VPWR.n42 0.123
R203 VPWR.n7 VPWR.n4 0.119
R204 VPWR.n9 VPWR.n7 0.119
R205 VPWR.n13 VPWR.n9 0.119
R206 VPWR.n15 VPWR.n13 0.119
R207 VPWR.n17 VPWR.n15 0.119
R208 VPWR.n19 VPWR.n17 0.119
R209 VPWR.n21 VPWR.n19 0.119
R210 VPWR.n23 VPWR.n21 0.119
R211 VPWR.n27 VPWR.n23 0.119
R212 VPWR.n29 VPWR.n27 0.119
R213 VPWR.n31 VPWR.n29 0.119
R214 VPWR.n33 VPWR.n31 0.119
R215 VPWR.n35 VPWR.n33 0.119
R216 VPWR.n37 VPWR.n35 0.119
R217 VPWR.n39 VPWR.n37 0.119
R218 D.n0 D.t1 302.729
R219 D.n0 D.t0 212.756
R220 D D.n0 94.057
R221 a_381_47.n1 a_381_47.n0 511.303
R222 a_381_47.n1 a_381_47.t2 90
R223 a_381_47.n0 a_381_47.t3 65.666
R224 a_381_47.n0 a_381_47.t1 63.321
R225 a_381_47.n2 a_381_47.t0 26.393
R226 a_381_47.n3 a_381_47.n2 14.4
R227 a_381_47.n2 a_381_47.n1 5
R228 a_1589_47.t1 a_1589_47.n2 243.368
R229 a_1589_47.n0 a_1589_47.t2 212.079
R230 a_1589_47.n1 a_1589_47.t4 212.079
R231 a_1589_47.n2 a_1589_47.t0 161.917
R232 a_1589_47.n0 a_1589_47.t3 139.779
R233 a_1589_47.n1 a_1589_47.t5 139.779
R234 a_1589_47.n2 a_1589_47.n1 111.448
R235 a_1589_47.n1 a_1589_47.n0 61.345
R236 a_592_47.t0 a_592_47.t1 99.726
R237 Q_N Q_N.n1 145.582
R238 Q_N Q_N.n0 108.927
R239 Q_N.n0 Q_N.t3 26.595
R240 Q_N.n0 Q_N.t2 26.595
R241 Q_N.n1 Q_N.t1 24.923
R242 Q_N.n1 Q_N.t0 24.923
R243 a_975_413.t0 a_975_413.t1 197
R244 a_1017_47.t0 a_1017_47.t1 93.059
C0 VPWR VPB 0.21fF
C1 VGND Q_N 0.21fF
C2 VPWR Q_N 0.32fF
C3 VGND Q 0.15fF
C4 VPWR Q 0.25fF
C5 VPWR VGND 0.17fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__dfxtp_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__dfxtp_1 Q CLK D VPWR VGND VNB VPB
X0 Q.t0 a_1059_315.t2 VGND.t4 VNB.t9 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 a_891_413.t3 a_193_47.t2 a_634_159.t3 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X2 a_561_413.t0 a_27_47.t2 a_466_413.t0 VPB.t8 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3 VPWR.t0 CLK.t0 a_27_47.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X4 Q.t1 a_1059_315.t3 VPWR.t3 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 a_381_47.t1 D.t0 VPWR.t1 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 VGND.t1 a_634_159.t4 a_592_47.t0 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7 VPWR.t5 a_891_413.t4 a_1059_315.t0 VPB.t5 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 a_466_413.t2 a_193_47.t3 a_381_47.t3 VPB.t11 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9 VPWR.t7 a_634_159.t5 a_561_413.t1 VPB.t9 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10 a_634_159.t1 a_466_413.t4 VGND.t6 VNB.t10 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X11 a_634_159.t2 a_466_413.t5 VPWR.t2 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X12 a_975_413.t1 a_193_47.t4 a_891_413.t2 VPB.t10 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13 VGND.t5 a_1059_315.t4 a_1017_47.t0 VNB.t8 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14 a_193_47.t0 a_27_47.t3 VGND.t2 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15 a_891_413.t0 a_27_47.t4 a_634_159.t0 VPB.t7 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16 a_592_47.t1 a_193_47.t5 a_466_413.t3 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X17 a_1017_47.t1 a_27_47.t5 a_891_413.t1 VNB.t5 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X18 VPWR.t4 a_1059_315.t5 a_975_413.t0 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19 a_466_413.t1 a_27_47.t6 a_381_47.t2 VNB.t6 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X20 a_193_47.t1 a_27_47.t7 VPWR.t6 VPB.t6 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X21 VGND.t0 a_891_413.t5 a_1059_315.t1 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X22 a_381_47.t0 D.t1 VGND.t3 VNB.t7 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23 VGND.t7 CLK.t1 a_27_47.t1 VNB.t11 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
R0 a_1059_315.n2 a_1059_315.t4 382.743
R1 a_1059_315.n0 a_1059_315.t3 241.534
R2 a_1059_315.n0 a_1059_315.t2 169.234
R3 a_1059_315.n2 a_1059_315.t5 138.53
R4 a_1059_315.t0 a_1059_315.n3 128.779
R5 a_1059_315.n1 a_1059_315.t1 103.313
R6 a_1059_315.n1 a_1059_315.n0 97.915
R7 a_1059_315.n3 a_1059_315.n2 97.786
R8 a_1059_315.n3 a_1059_315.n1 16.622
R9 VGND.n1 VGND.t5 158.499
R10 VGND.n20 VGND.t3 150.527
R11 VGND.n2 VGND.n0 131.571
R12 VGND.n25 VGND.n24 107.239
R13 VGND.n12 VGND.n11 107.029
R14 VGND.n11 VGND.t6 74.865
R15 VGND.n11 VGND.t1 40
R16 VGND.n24 VGND.t2 38.571
R17 VGND.n24 VGND.t7 38.571
R18 VGND.n0 VGND.t4 24.923
R19 VGND.n0 VGND.t0 24.923
R20 VGND.n4 VGND.n3 4.65
R21 VGND.n6 VGND.n5 4.65
R22 VGND.n8 VGND.n7 4.65
R23 VGND.n10 VGND.n9 4.65
R24 VGND.n13 VGND.n12 4.65
R25 VGND.n15 VGND.n14 4.65
R26 VGND.n17 VGND.n16 4.65
R27 VGND.n19 VGND.n18 4.65
R28 VGND.n21 VGND.n20 4.65
R29 VGND.n23 VGND.n22 4.65
R30 VGND.n2 VGND.n1 4.018
R31 VGND.n26 VGND.n25 3.932
R32 VGND.n4 VGND.n2 0.214
R33 VGND.n26 VGND.n23 0.137
R34 VGND VGND.n26 0.123
R35 VGND.n6 VGND.n4 0.119
R36 VGND.n8 VGND.n6 0.119
R37 VGND.n10 VGND.n8 0.119
R38 VGND.n13 VGND.n10 0.119
R39 VGND.n15 VGND.n13 0.119
R40 VGND.n17 VGND.n15 0.119
R41 VGND.n19 VGND.n17 0.119
R42 VGND.n21 VGND.n19 0.119
R43 VGND.n23 VGND.n21 0.119
R44 Q.n0 Q.t1 221.7
R45 Q.n0 Q.t0 82.859
R46 Q Q.n0 5.75
R47 VNB.t4 VNB.t7 6082.35
R48 VNB.t8 VNB.t0 5354.23
R49 VNB VNB.t11 4270.59
R50 VNB.t7 VNB.t6 3623.53
R51 VNB.t2 VNB.t5 3429.41
R52 VNB.t3 VNB.t1 3202.94
R53 VNB.t6 VNB.t3 3202.94
R54 VNB.t1 VNB.t10 3130.33
R55 VNB.t5 VNB.t8 3073.53
R56 VNB.t11 VNB.t4 2717.65
R57 VNB.t10 VNB.t2 2363.68
R58 VNB.t0 VNB.t9 2030.77
R59 a_193_47.n1 a_193_47.t5 407.215
R60 a_193_47.n1 a_193_47.t3 273.571
R61 a_193_47.t1 a_193_47.n3 246.213
R62 a_193_47.n0 a_193_47.t4 232.651
R63 a_193_47.n0 a_193_47.t2 222.372
R64 a_193_47.n3 a_193_47.t0 201.643
R65 a_193_47.n2 a_193_47.n1 90.25
R66 a_193_47.n2 a_193_47.n0 6.797
R67 a_193_47.n3 a_193_47.n2 5.609
R68 a_634_159.n1 a_634_159.t5 406.399
R69 a_634_159.n3 a_634_159.n2 381.512
R70 a_634_159.n1 a_634_159.t4 130.052
R71 a_634_159.n2 a_634_159.n0 121.487
R72 a_634_159.n2 a_634_159.n1 104.16
R73 a_634_159.n3 a_634_159.t0 89.119
R74 a_634_159.n0 a_634_159.t3 71.666
R75 a_634_159.t2 a_634_159.n3 37.523
R76 a_634_159.n0 a_634_159.t1 28.437
R77 a_891_413.n3 a_891_413.n2 403.558
R78 a_891_413.n1 a_891_413.t4 212.079
R79 a_891_413.n2 a_891_413.n1 174.914
R80 a_891_413.n2 a_891_413.n0 166.287
R81 a_891_413.n1 a_891_413.t5 141.239
R82 a_891_413.n0 a_891_413.t1 76.666
R83 a_891_413.n3 a_891_413.t2 63.321
R84 a_891_413.t0 a_891_413.n3 63.321
R85 a_891_413.n0 a_891_413.t3 50
R86 a_27_47.n2 a_27_47.t5 443.438
R87 a_27_47.n3 a_27_47.t6 270.054
R88 a_27_47.n4 a_27_47.t7 263.171
R89 a_27_47.n2 a_27_47.t4 254.388
R90 a_27_47.t0 a_27_47.n6 243.779
R91 a_27_47.n4 a_27_47.t3 227.825
R92 a_27_47.n5 a_27_47.t1 195.494
R93 a_27_47.n0 a_27_47.t2 142.671
R94 a_27_47.n1 a_27_47.n2 112.935
R95 a_27_47.n5 a_27_47.n4 76
R96 a_27_47.n6 a_27_47.n5 35.339
R97 a_27_47.n6 a_27_47.n1 6.379
R98 a_27_47.n1 a_27_47.n0 4.695
R99 a_27_47.n0 a_27_47.n3 2.98
R100 a_466_413.n3 a_466_413.n2 403.181
R101 a_466_413.n0 a_466_413.t4 230.482
R102 a_466_413.n2 a_466_413.n1 205.859
R103 a_466_413.n0 a_466_413.t5 196.013
R104 a_466_413.n2 a_466_413.n0 92.738
R105 a_466_413.n3 a_466_413.t2 79.738
R106 a_466_413.t0 a_466_413.n3 72.702
R107 a_466_413.n1 a_466_413.t3 70
R108 a_466_413.n1 a_466_413.t1 45
R109 a_561_413.t0 a_561_413.t1 171.202
R110 VPB.t3 VPB.t5 621.495
R111 VPB.t6 VPB.t1 556.386
R112 VPB.t9 VPB.t2 390.654
R113 VPB.t10 VPB.t3 337.383
R114 VPB.t8 VPB.t9 304.828
R115 VPB.t2 VPB.t7 281.152
R116 VPB.t11 VPB.t8 281.152
R117 VPB.t1 VPB.t11 251.557
R118 VPB.t5 VPB.t4 248.598
R119 VPB.t7 VPB.t10 248.598
R120 VPB.t0 VPB.t6 248.598
R121 VPB VPB.t0 142.056
R122 CLK.n0 CLK.t0 294.554
R123 CLK.n0 CLK.t1 211.008
R124 CLK CLK.n0 77.969
R125 VPWR.n1 VPWR.t4 375.232
R126 VPWR.n21 VPWR.t1 374.175
R127 VPWR.n26 VPWR.n25 311.893
R128 VPWR.n2 VPWR.n0 192.981
R129 VPWR.n10 VPWR.n9 174.594
R130 VPWR.n9 VPWR.t7 113.978
R131 VPWR.n25 VPWR.t6 41.554
R132 VPWR.n25 VPWR.t0 41.554
R133 VPWR.n9 VPWR.t2 35.46
R134 VPWR.n0 VPWR.t3 26.595
R135 VPWR.n0 VPWR.t5 26.595
R136 VPWR.n11 VPWR.n10 16.188
R137 VPWR.n4 VPWR.n3 4.65
R138 VPWR.n6 VPWR.n5 4.65
R139 VPWR.n8 VPWR.n7 4.65
R140 VPWR.n12 VPWR.n11 4.65
R141 VPWR.n14 VPWR.n13 4.65
R142 VPWR.n16 VPWR.n15 4.65
R143 VPWR.n18 VPWR.n17 4.65
R144 VPWR.n20 VPWR.n19 4.65
R145 VPWR.n22 VPWR.n21 4.65
R146 VPWR.n24 VPWR.n23 4.65
R147 VPWR.n2 VPWR.n1 3.996
R148 VPWR.n27 VPWR.n26 3.932
R149 VPWR.n4 VPWR.n2 0.225
R150 VPWR.n27 VPWR.n24 0.137
R151 VPWR VPWR.n27 0.123
R152 VPWR.n6 VPWR.n4 0.119
R153 VPWR.n8 VPWR.n6 0.119
R154 VPWR.n12 VPWR.n8 0.119
R155 VPWR.n14 VPWR.n12 0.119
R156 VPWR.n16 VPWR.n14 0.119
R157 VPWR.n18 VPWR.n16 0.119
R158 VPWR.n20 VPWR.n18 0.119
R159 VPWR.n22 VPWR.n20 0.119
R160 VPWR.n24 VPWR.n22 0.119
R161 D.n0 D.t1 302.729
R162 D.n0 D.t0 212.756
R163 D D.n0 94.057
R164 a_381_47.n1 a_381_47.n0 511.303
R165 a_381_47.n1 a_381_47.t2 90
R166 a_381_47.n0 a_381_47.t3 65.666
R167 a_381_47.n0 a_381_47.t1 63.321
R168 a_381_47.n2 a_381_47.t0 26.393
R169 a_381_47.n3 a_381_47.n2 14.4
R170 a_381_47.n2 a_381_47.n1 5
R171 a_592_47.t0 a_592_47.t1 99.726
R172 a_975_413.t0 a_975_413.t1 197
R173 a_1017_47.t0 a_1017_47.t1 93.059
C0 VGND Q 0.11fF
C1 VPWR Q 0.16fF
C2 VPB VPWR 0.15fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__dfxtp_2.ext - technology: sky130A

.subckt sky130_fd_sc_hd__dfxtp_2 Q CLK D VPWR VGND VNB VPB
X0 Q.t2 a_1059_315.t2 VGND.t3 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 a_891_413.t3 a_193_47.t2 a_634_159.t3 VNB.t11 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X2 VPWR.t2 a_1059_315.t3 Q.t0 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 a_561_413.t0 a_27_47.t2 a_466_413.t0 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 VPWR.t6 CLK.t0 a_27_47.t0 VPB.t10 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X5 Q.t3 a_1059_315.t4 VPWR.t1 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 a_381_47.t3 D.t0 VPWR.t5 VPB.t7 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7 VGND.t0 a_634_159.t4 a_592_47.t1 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 VGND.t1 a_1059_315.t5 Q.t1 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 VPWR.t7 a_891_413.t4 a_1059_315.t0 VPB.t11 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 a_466_413.t2 a_193_47.t3 a_381_47.t1 VPB.t9 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11 VPWR.t8 a_634_159.t5 a_561_413.t1 VPB.t12 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12 a_634_159.t1 a_466_413.t4 VGND.t5 VNB.t7 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X13 a_634_159.t2 a_466_413.t5 VPWR.t4 VPB.t6 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X14 a_975_413.t1 a_193_47.t4 a_891_413.t2 VPB.t8 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15 VGND.t2 a_1059_315.t6 a_1017_47.t1 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16 a_193_47.t0 a_27_47.t3 VGND.t4 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17 a_891_413.t0 a_27_47.t4 a_634_159.t0 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18 a_592_47.t0 a_193_47.t5 a_466_413.t3 VNB.t12 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X19 a_1017_47.t0 a_27_47.t5 a_891_413.t1 VNB.t5 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X20 VPWR.t0 a_1059_315.t7 a_975_413.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21 a_466_413.t1 a_27_47.t6 a_381_47.t0 VNB.t6 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X22 a_193_47.t1 a_27_47.t7 VPWR.t3 VPB.t5 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X23 VGND.t7 a_891_413.t5 a_1059_315.t1 VNB.t9 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X24 a_381_47.t2 D.t1 VGND.t6 VNB.t8 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X25 VGND.t8 CLK.t1 a_27_47.t1 VNB.t10 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
R0 a_1059_315.n3 a_1059_315.t6 382.743
R1 a_1059_315.n1 a_1059_315.t4 213.539
R2 a_1059_315.n0 a_1059_315.t3 212.079
R3 a_1059_315.n0 a_1059_315.t5 141.239
R4 a_1059_315.n1 a_1059_315.t2 139.779
R5 a_1059_315.n3 a_1059_315.t7 138.53
R6 a_1059_315.t0 a_1059_315.n4 128.779
R7 a_1059_315.n2 a_1059_315.t1 103.313
R8 a_1059_315.n2 a_1059_315.n1 97.915
R9 a_1059_315.n4 a_1059_315.n3 97.786
R10 a_1059_315.n1 a_1059_315.n0 59.884
R11 a_1059_315.n4 a_1059_315.n2 16.622
R12 VGND.n5 VGND.t2 158.499
R13 VGND.n2 VGND.t1 152.87
R14 VGND.n24 VGND.t6 150.527
R15 VGND.n1 VGND.n0 126.005
R16 VGND.n29 VGND.n28 107.239
R17 VGND.n16 VGND.n15 107.029
R18 VGND.n15 VGND.t5 74.865
R19 VGND.n15 VGND.t0 40
R20 VGND.n28 VGND.t4 38.571
R21 VGND.n28 VGND.t8 38.571
R22 VGND.n0 VGND.t3 24.923
R23 VGND.n0 VGND.t7 24.923
R24 VGND.n2 VGND.n1 6.252
R25 VGND.n4 VGND.n3 4.65
R26 VGND.n6 VGND.n5 4.65
R27 VGND.n8 VGND.n7 4.65
R28 VGND.n10 VGND.n9 4.65
R29 VGND.n12 VGND.n11 4.65
R30 VGND.n14 VGND.n13 4.65
R31 VGND.n17 VGND.n16 4.65
R32 VGND.n19 VGND.n18 4.65
R33 VGND.n21 VGND.n20 4.65
R34 VGND.n23 VGND.n22 4.65
R35 VGND.n25 VGND.n24 4.65
R36 VGND.n27 VGND.n26 4.65
R37 VGND.n30 VGND.n29 3.932
R38 VGND.n4 VGND.n2 0.279
R39 VGND.n30 VGND.n27 0.137
R40 VGND VGND.n30 0.123
R41 VGND.n6 VGND.n4 0.119
R42 VGND.n8 VGND.n6 0.119
R43 VGND.n10 VGND.n8 0.119
R44 VGND.n12 VGND.n10 0.119
R45 VGND.n14 VGND.n12 0.119
R46 VGND.n17 VGND.n14 0.119
R47 VGND.n19 VGND.n17 0.119
R48 VGND.n21 VGND.n19 0.119
R49 VGND.n23 VGND.n21 0.119
R50 VGND.n25 VGND.n23 0.119
R51 VGND.n27 VGND.n25 0.119
R52 Q.n1 Q.n0 189.237
R53 Q Q.n2 93.663
R54 Q.n0 Q.t0 26.595
R55 Q.n0 Q.t3 26.595
R56 Q.n2 Q.t1 24.923
R57 Q.n2 Q.t2 24.923
R58 Q Q.n1 12.024
R59 VNB.t4 VNB.t8 6082.35
R60 VNB.t1 VNB.t9 5354.23
R61 VNB VNB.t10 4270.59
R62 VNB.t8 VNB.t6 3623.53
R63 VNB.t11 VNB.t5 3429.41
R64 VNB.t12 VNB.t0 3202.94
R65 VNB.t6 VNB.t12 3202.94
R66 VNB.t0 VNB.t7 3130.33
R67 VNB.t5 VNB.t1 3073.53
R68 VNB.t10 VNB.t4 2717.65
R69 VNB.t7 VNB.t11 2363.68
R70 VNB.t3 VNB.t2 2030.77
R71 VNB.t9 VNB.t3 2030.77
R72 a_193_47.n1 a_193_47.t5 407.215
R73 a_193_47.n1 a_193_47.t3 273.571
R74 a_193_47.t1 a_193_47.n3 246.213
R75 a_193_47.n0 a_193_47.t4 232.651
R76 a_193_47.n0 a_193_47.t2 222.372
R77 a_193_47.n3 a_193_47.t0 201.643
R78 a_193_47.n2 a_193_47.n1 90.25
R79 a_193_47.n2 a_193_47.n0 6.797
R80 a_193_47.n3 a_193_47.n2 5.609
R81 a_634_159.n1 a_634_159.t5 406.399
R82 a_634_159.n3 a_634_159.n2 381.512
R83 a_634_159.n1 a_634_159.t4 130.052
R84 a_634_159.n2 a_634_159.n0 121.487
R85 a_634_159.n2 a_634_159.n1 104.16
R86 a_634_159.n3 a_634_159.t0 89.119
R87 a_634_159.n0 a_634_159.t3 71.666
R88 a_634_159.t2 a_634_159.n3 37.523
R89 a_634_159.n0 a_634_159.t1 28.437
R90 a_891_413.n3 a_891_413.n2 403.558
R91 a_891_413.n1 a_891_413.t4 212.079
R92 a_891_413.n2 a_891_413.n1 174.914
R93 a_891_413.n2 a_891_413.n0 166.287
R94 a_891_413.n1 a_891_413.t5 141.239
R95 a_891_413.n0 a_891_413.t1 76.666
R96 a_891_413.n3 a_891_413.t2 63.321
R97 a_891_413.t0 a_891_413.n3 63.321
R98 a_891_413.n0 a_891_413.t3 50
R99 VPWR.n5 VPWR.t0 375.232
R100 VPWR.n25 VPWR.t5 374.175
R101 VPWR.n30 VPWR.n29 311.893
R102 VPWR.n2 VPWR.t2 219.222
R103 VPWR.n1 VPWR.n0 186.917
R104 VPWR.n14 VPWR.n13 174.594
R105 VPWR.n13 VPWR.t8 113.978
R106 VPWR.n29 VPWR.t3 41.554
R107 VPWR.n29 VPWR.t6 41.554
R108 VPWR.n13 VPWR.t4 35.46
R109 VPWR.n0 VPWR.t1 26.595
R110 VPWR.n0 VPWR.t7 26.595
R111 VPWR.n15 VPWR.n14 16.188
R112 VPWR.n2 VPWR.n1 6.997
R113 VPWR.n4 VPWR.n3 4.65
R114 VPWR.n6 VPWR.n5 4.65
R115 VPWR.n8 VPWR.n7 4.65
R116 VPWR.n10 VPWR.n9 4.65
R117 VPWR.n12 VPWR.n11 4.65
R118 VPWR.n16 VPWR.n15 4.65
R119 VPWR.n18 VPWR.n17 4.65
R120 VPWR.n20 VPWR.n19 4.65
R121 VPWR.n22 VPWR.n21 4.65
R122 VPWR.n24 VPWR.n23 4.65
R123 VPWR.n26 VPWR.n25 4.65
R124 VPWR.n28 VPWR.n27 4.65
R125 VPWR.n31 VPWR.n30 3.932
R126 VPWR.n4 VPWR.n2 0.288
R127 VPWR.n31 VPWR.n28 0.137
R128 VPWR VPWR.n31 0.123
R129 VPWR.n6 VPWR.n4 0.119
R130 VPWR.n8 VPWR.n6 0.119
R131 VPWR.n10 VPWR.n8 0.119
R132 VPWR.n12 VPWR.n10 0.119
R133 VPWR.n16 VPWR.n12 0.119
R134 VPWR.n18 VPWR.n16 0.119
R135 VPWR.n20 VPWR.n18 0.119
R136 VPWR.n22 VPWR.n20 0.119
R137 VPWR.n24 VPWR.n22 0.119
R138 VPWR.n26 VPWR.n24 0.119
R139 VPWR.n28 VPWR.n26 0.119
R140 VPB.t0 VPB.t11 621.495
R141 VPB.t5 VPB.t7 556.386
R142 VPB.t12 VPB.t6 390.654
R143 VPB.t8 VPB.t0 337.383
R144 VPB.t3 VPB.t12 304.828
R145 VPB.t6 VPB.t4 281.152
R146 VPB.t9 VPB.t3 281.152
R147 VPB.t7 VPB.t9 251.557
R148 VPB.t1 VPB.t2 248.598
R149 VPB.t11 VPB.t1 248.598
R150 VPB.t4 VPB.t8 248.598
R151 VPB.t10 VPB.t5 248.598
R152 VPB VPB.t10 142.056
R153 a_27_47.n2 a_27_47.t5 443.438
R154 a_27_47.n3 a_27_47.t6 270.054
R155 a_27_47.n4 a_27_47.t7 263.171
R156 a_27_47.n2 a_27_47.t4 254.388
R157 a_27_47.t0 a_27_47.n6 243.779
R158 a_27_47.n4 a_27_47.t3 227.825
R159 a_27_47.n5 a_27_47.t1 195.494
R160 a_27_47.n0 a_27_47.t2 142.671
R161 a_27_47.n1 a_27_47.n2 112.935
R162 a_27_47.n5 a_27_47.n4 76
R163 a_27_47.n6 a_27_47.n5 35.339
R164 a_27_47.n6 a_27_47.n1 6.379
R165 a_27_47.n1 a_27_47.n0 4.695
R166 a_27_47.n0 a_27_47.n3 2.98
R167 a_466_413.n3 a_466_413.n2 403.181
R168 a_466_413.n0 a_466_413.t4 230.482
R169 a_466_413.n2 a_466_413.n1 205.859
R170 a_466_413.n0 a_466_413.t5 196.013
R171 a_466_413.n2 a_466_413.n0 92.738
R172 a_466_413.n3 a_466_413.t2 79.738
R173 a_466_413.t0 a_466_413.n3 72.702
R174 a_466_413.n1 a_466_413.t3 70
R175 a_466_413.n1 a_466_413.t1 45
R176 a_561_413.t0 a_561_413.t1 171.202
R177 CLK.n0 CLK.t0 294.554
R178 CLK.n0 CLK.t1 211.008
R179 CLK CLK.n0 77.969
R180 D.n0 D.t1 302.729
R181 D.n0 D.t0 212.756
R182 D D.n0 94.057
R183 a_381_47.n1 a_381_47.n0 511.303
R184 a_381_47.n0 a_381_47.t0 90
R185 a_381_47.t1 a_381_47.n1 65.666
R186 a_381_47.n1 a_381_47.t3 63.321
R187 a_381_47.n0 a_381_47.t2 31.393
R188 a_592_47.t1 a_592_47.t0 99.726
R189 a_975_413.t0 a_975_413.t1 197
R190 a_1017_47.t1 a_1017_47.t0 93.059
C0 VPB VPWR 0.17fF
C1 VGND Q 0.15fF
C2 VPWR Q 0.25fF
C3 VPWR VGND 0.11fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__dfxtp_4.ext - technology: sky130A

.subckt sky130_fd_sc_hd__dfxtp_4 VGND VPWR D CLK Q VNB VPB
X0 Q.t3 a_1062_300.t2 VPWR.t8 VPB.t10 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_1020_47.t0 a_27_47.t2 a_891_413.t3 VNB.t7 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X2 a_572_47.t1 a_193_47.t2 a_475_413.t2 VNB.t14 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X3 VPWR.t4 a_1062_300.t3 a_975_413.t0 VPB.t9 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 a_634_183.t1 a_475_413.t4 VGND.t4 VNB.t13 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X5 VPWR.t0 CLK.t0 a_27_47.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X6 a_381_47.t0 D.t0 VPWR.t3 VPB.t5 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7 a_475_413.t0 a_27_47.t3 a_381_47.t2 VNB.t6 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X8 VGND.t10 a_1062_300.t4 a_1020_47.t1 VNB.t12 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9 VPWR.t1 a_634_183.t4 a_568_413.t0 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10 Q.t7 a_1062_300.t5 VGND.t9 VNB.t11 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 a_568_413.t1 a_27_47.t4 a_475_413.t1 VPB.t11 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12 a_634_183.t0 a_475_413.t5 VPWR.t10 VPB.t14 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X13 a_975_413.t1 a_193_47.t3 a_891_413.t0 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14 a_193_47.t1 a_27_47.t5 VGND.t5 VNB.t5 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15 a_891_413.t2 a_27_47.t6 a_634_183.t2 VPB.t12 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16 Q.t6 a_1062_300.t6 VGND.t8 VNB.t10 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X17 VGND.t2 a_891_413.t4 a_1062_300.t0 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X18 VPWR.t7 a_1062_300.t7 Q.t2 VPB.t8 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X19 VGND.t7 a_1062_300.t8 Q.t5 VNB.t9 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X20 Q.t1 a_1062_300.t9 VPWR.t6 VPB.t7 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X21 a_193_47.t0 a_27_47.t7 VPWR.t9 VPB.t13 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X22 VGND.t6 a_1062_300.t10 Q.t4 VNB.t8 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X23 a_381_47.t1 D.t1 VGND.t3 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24 VPWR.t2 a_891_413.t5 a_1062_300.t1 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X25 a_891_413.t1 a_193_47.t4 a_634_183.t3 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X26 a_475_413.t3 a_193_47.t5 a_381_47.t3 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X27 VGND.t1 a_634_183.t5 a_572_47.t0 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X28 VGND.t0 CLK.t1 a_27_47.t1 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X29 VPWR.t5 a_1062_300.t11 Q.t0 VPB.t6 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
R0 a_1062_300.n12 a_1062_300.t4 359.398
R1 a_1062_300.n0 a_1062_300.t11 212.079
R2 a_1062_300.n2 a_1062_300.t2 212.079
R3 a_1062_300.n5 a_1062_300.t7 212.079
R4 a_1062_300.n8 a_1062_300.t9 212.079
R5 a_1062_300.n12 a_1062_300.t3 163.385
R6 a_1062_300.n0 a_1062_300.t8 139.779
R7 a_1062_300.n2 a_1062_300.t5 139.779
R8 a_1062_300.n5 a_1062_300.t10 139.779
R9 a_1062_300.n8 a_1062_300.t6 139.779
R10 a_1062_300.t1 a_1062_300.n13 130.613
R11 a_1062_300.n11 a_1062_300.t0 119.251
R12 a_1062_300.n13 a_1062_300.n12 102.763
R13 a_1062_300.n4 a_1062_300.n1 101.6
R14 a_1062_300.n4 a_1062_300.n3 76
R15 a_1062_300.n7 a_1062_300.n6 76
R16 a_1062_300.n10 a_1062_300.n9 76
R17 a_1062_300.n11 a_1062_300.n10 41.411
R18 a_1062_300.n13 a_1062_300.n11 34.919
R19 a_1062_300.n7 a_1062_300.n4 25.6
R20 a_1062_300.n10 a_1062_300.n7 25.6
R21 a_1062_300.n1 a_1062_300.n0 20.448
R22 a_1062_300.n9 a_1062_300.n8 16.796
R23 a_1062_300.n3 a_1062_300.n2 8.763
R24 a_1062_300.n6 a_1062_300.n5 5.112
R25 VPWR.n10 VPWR.t4 380.825
R26 VPWR.n31 VPWR.t3 374.175
R27 VPWR.n36 VPWR.n35 311.893
R28 VPWR.n2 VPWR.t5 211.729
R29 VPWR.n6 VPWR.n5 177.655
R30 VPWR.n1 VPWR.n0 176.853
R31 VPWR.n20 VPWR.n19 174.594
R32 VPWR.n19 VPWR.t1 113.978
R33 VPWR.n35 VPWR.t9 41.554
R34 VPWR.n35 VPWR.t0 41.554
R35 VPWR.n19 VPWR.t10 35.46
R36 VPWR.n5 VPWR.t2 33.49
R37 VPWR.n5 VPWR.t6 30.535
R38 VPWR.n0 VPWR.t7 29.55
R39 VPWR.n0 VPWR.t8 26.595
R40 VPWR.n21 VPWR.n20 16.188
R41 VPWR.n4 VPWR.n3 4.65
R42 VPWR.n7 VPWR.n6 4.65
R43 VPWR.n9 VPWR.n8 4.65
R44 VPWR.n12 VPWR.n11 4.65
R45 VPWR.n14 VPWR.n13 4.65
R46 VPWR.n16 VPWR.n15 4.65
R47 VPWR.n18 VPWR.n17 4.65
R48 VPWR.n22 VPWR.n21 4.65
R49 VPWR.n24 VPWR.n23 4.65
R50 VPWR.n26 VPWR.n25 4.65
R51 VPWR.n28 VPWR.n27 4.65
R52 VPWR.n30 VPWR.n29 4.65
R53 VPWR.n32 VPWR.n31 4.65
R54 VPWR.n34 VPWR.n33 4.65
R55 VPWR.n2 VPWR.n1 4.392
R56 VPWR.n37 VPWR.n36 3.932
R57 VPWR.n11 VPWR.n10 3.388
R58 VPWR.n4 VPWR.n2 0.258
R59 VPWR.n37 VPWR.n34 0.137
R60 VPWR VPWR.n37 0.123
R61 VPWR.n7 VPWR.n4 0.119
R62 VPWR.n9 VPWR.n7 0.119
R63 VPWR.n12 VPWR.n9 0.119
R64 VPWR.n14 VPWR.n12 0.119
R65 VPWR.n16 VPWR.n14 0.119
R66 VPWR.n18 VPWR.n16 0.119
R67 VPWR.n22 VPWR.n18 0.119
R68 VPWR.n24 VPWR.n22 0.119
R69 VPWR.n26 VPWR.n24 0.119
R70 VPWR.n28 VPWR.n26 0.119
R71 VPWR.n30 VPWR.n28 0.119
R72 VPWR.n32 VPWR.n30 0.119
R73 VPWR.n34 VPWR.n32 0.119
R74 Q.n7 Q.n6 292.5
R75 Q.n8 Q.n7 146.531
R76 Q.n5 Q.n4 107.635
R77 Q Q.n0 93.646
R78 Q.n1 Q.n0 92.5
R79 Q.n5 Q.n3 74.164
R80 Q.n3 Q.n2 52.342
R81 Q.n3 Q.n1 42.208
R82 Q.n6 Q.n5 42.208
R83 Q.n7 Q.t2 26.595
R84 Q.n7 Q.t1 26.595
R85 Q.n4 Q.t0 26.595
R86 Q.n4 Q.t3 26.595
R87 Q.n0 Q.t4 24.923
R88 Q.n0 Q.t6 24.923
R89 Q.n2 Q.t5 24.923
R90 Q.n2 Q.t7 24.923
R91 Q.n1 Q 11.844
R92 Q.n8 Q 9.965
R93 Q.n6 Q 5.922
R94 Q Q.n8 2.967
R95 VPB.t9 VPB.t2 639.252
R96 VPB.t13 VPB.t5 556.386
R97 VPB.t1 VPB.t14 390.654
R98 VPB.t3 VPB.t9 346.261
R99 VPB.t11 VPB.t1 284.112
R100 VPB.t2 VPB.t7 281.152
R101 VPB.t14 VPB.t12 281.152
R102 VPB.t5 VPB.t4 278.193
R103 VPB.t4 VPB.t11 275.233
R104 VPB.t8 VPB.t10 257.476
R105 VPB.t10 VPB.t6 248.598
R106 VPB.t7 VPB.t8 248.598
R107 VPB.t12 VPB.t3 248.598
R108 VPB.t0 VPB.t13 248.598
R109 VPB VPB.t0 142.056
R110 a_27_47.n1 a_27_47.t3 501.814
R111 a_27_47.n0 a_27_47.t2 448.258
R112 a_27_47.n3 a_27_47.t7 263.171
R113 a_27_47.n0 a_27_47.t6 254.388
R114 a_27_47.t0 a_27_47.n5 243.779
R115 a_27_47.n3 a_27_47.t5 227.825
R116 a_27_47.n4 a_27_47.t1 195.494
R117 a_27_47.n1 a_27_47.t4 148.348
R118 a_27_47.n2 a_27_47.n0 112.768
R119 a_27_47.n2 a_27_47.n1 87.5
R120 a_27_47.n4 a_27_47.n3 76
R121 a_27_47.n5 a_27_47.n4 35.339
R122 a_27_47.n5 a_27_47.n2 6.618
R123 a_891_413.n3 a_891_413.n2 409.581
R124 a_891_413.n1 a_891_413.t5 212.079
R125 a_891_413.n2 a_891_413.n1 197.671
R126 a_891_413.n2 a_891_413.n0 164.781
R127 a_891_413.n1 a_891_413.t4 139.779
R128 a_891_413.n0 a_891_413.t1 73.333
R129 a_891_413.t0 a_891_413.n3 63.321
R130 a_891_413.n3 a_891_413.t2 63.321
R131 a_891_413.n0 a_891_413.t3 48.333
R132 a_1020_47.t1 a_1020_47.t0 93.059
R133 VNB.t5 VNB.t4 6082.35
R134 VNB.t12 VNB.t3 5483.65
R135 VNB VNB.t0 4270.59
R136 VNB.t1 VNB.t13 4003.85
R137 VNB.t2 VNB.t7 3332.35
R138 VNB.t14 VNB.t1 3170.59
R139 VNB.t6 VNB.t14 3105.88
R140 VNB.t7 VNB.t12 3073.53
R141 VNB.t4 VNB.t6 3073.53
R142 VNB.t0 VNB.t5 2717.65
R143 VNB.t13 VNB.t2 2363.68
R144 VNB.t3 VNB.t10 2296.7
R145 VNB.t8 VNB.t11 2103.3
R146 VNB.t11 VNB.t9 2030.77
R147 VNB.t10 VNB.t8 2030.77
R148 a_193_47.t0 a_193_47.n3 278.596
R149 a_193_47.n0 a_193_47.t3 272.659
R150 a_193_47.n1 a_193_47.t5 269.802
R151 a_193_47.n1 a_193_47.t2 205.234
R152 a_193_47.n0 a_193_47.t4 195.261
R153 a_193_47.n3 a_193_47.t1 150.413
R154 a_193_47.n2 a_193_47.n0 14.334
R155 a_193_47.n3 a_193_47.n2 5.797
R156 a_193_47.n2 a_193_47.n1 4.65
R157 a_475_413.n3 a_475_413.n2 400.546
R158 a_475_413.n0 a_475_413.t4 226.539
R159 a_475_413.n2 a_475_413.n1 208.495
R160 a_475_413.n0 a_475_413.t5 196.013
R161 a_475_413.n2 a_475_413.n0 92.738
R162 a_475_413.n3 a_475_413.t3 75.047
R163 a_475_413.t1 a_475_413.n3 72.702
R164 a_475_413.n1 a_475_413.t0 61.666
R165 a_475_413.n1 a_475_413.t2 48.333
R166 a_572_47.t0 a_572_47.t1 98.059
R167 a_975_413.t0 a_975_413.t1 204.035
R168 VGND.n2 VGND.t7 193.413
R169 VGND.n11 VGND.t10 158.553
R170 VGND.n31 VGND.t3 150.527
R171 VGND.n6 VGND.n5 116.217
R172 VGND.n1 VGND.n0 115.841
R173 VGND.n36 VGND.n35 107.239
R174 VGND.n23 VGND.n22 107.029
R175 VGND.n22 VGND.t1 87.142
R176 VGND.n22 VGND.t4 66.294
R177 VGND.n35 VGND.t5 38.571
R178 VGND.n35 VGND.t0 38.571
R179 VGND.n5 VGND.t2 31.384
R180 VGND.n5 VGND.t8 28.615
R181 VGND.n0 VGND.t6 26.769
R182 VGND.n0 VGND.t9 25.846
R183 VGND.n2 VGND.n1 4.772
R184 VGND.n4 VGND.n3 4.65
R185 VGND.n8 VGND.n7 4.65
R186 VGND.n10 VGND.n9 4.65
R187 VGND.n13 VGND.n12 4.65
R188 VGND.n15 VGND.n14 4.65
R189 VGND.n17 VGND.n16 4.65
R190 VGND.n19 VGND.n18 4.65
R191 VGND.n21 VGND.n20 4.65
R192 VGND.n24 VGND.n23 4.65
R193 VGND.n26 VGND.n25 4.65
R194 VGND.n28 VGND.n27 4.65
R195 VGND.n30 VGND.n29 4.65
R196 VGND.n32 VGND.n31 4.65
R197 VGND.n34 VGND.n33 4.65
R198 VGND.n37 VGND.n36 3.932
R199 VGND.n7 VGND.n6 3.011
R200 VGND.n12 VGND.n11 3.011
R201 VGND.n4 VGND.n2 0.254
R202 VGND.n37 VGND.n34 0.137
R203 VGND VGND.n37 0.123
R204 VGND.n8 VGND.n4 0.119
R205 VGND.n10 VGND.n8 0.119
R206 VGND.n13 VGND.n10 0.119
R207 VGND.n15 VGND.n13 0.119
R208 VGND.n17 VGND.n15 0.119
R209 VGND.n19 VGND.n17 0.119
R210 VGND.n21 VGND.n19 0.119
R211 VGND.n24 VGND.n21 0.119
R212 VGND.n26 VGND.n24 0.119
R213 VGND.n28 VGND.n26 0.119
R214 VGND.n30 VGND.n28 0.119
R215 VGND.n32 VGND.n30 0.119
R216 VGND.n34 VGND.n32 0.119
R217 a_634_183.n1 a_634_183.t4 433.799
R218 a_634_183.n3 a_634_183.n2 381.512
R219 a_634_183.n1 a_634_183.t5 128.098
R220 a_634_183.n2 a_634_183.n0 125.628
R221 a_634_183.n2 a_634_183.n1 109.306
R222 a_634_183.n3 a_634_183.t2 89.119
R223 a_634_183.n0 a_634_183.t3 63.333
R224 a_634_183.t0 a_634_183.n3 37.523
R225 a_634_183.n0 a_634_183.t1 36.77
R226 CLK.n0 CLK.t0 294.554
R227 CLK.n0 CLK.t1 211.008
R228 CLK.n1 CLK.n0 76
R229 CLK.n1 CLK 10.422
R230 CLK CLK.n1 2.011
R231 D.n0 D.t1 305.623
R232 D.n0 D.t0 215.65
R233 D D.n0 78.514
R234 a_381_47.n1 a_381_47.n0 514.934
R235 a_381_47.n1 a_381_47.t3 86.773
R236 a_381_47.t0 a_381_47.n1 63.321
R237 a_381_47.n0 a_381_47.t2 58.333
R238 a_381_47.n0 a_381_47.t1 34.726
R239 a_568_413.t0 a_568_413.t1 154.785
C0 VGND Q 0.36fF
C1 VPWR Q 0.55fF
C2 VPWR VGND 0.13fF
C3 VPB VPWR 0.18fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__diode_2.ext - technology: sky130A

.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VPWR VPB VNB
D0 VNB DIODE sky130_fd_pr__diode_pw2nd_05v5 pj=5.36e+06u area=4.347e+11p
R0 DIODE DIODE.t0 0.938
R1 DIODE.t0 DIODE 0.786
R2 VNB.n1 VNB 3882.35
R3 VNB.n1 VNB.n0 2348.31
R4 VNB VNB.n1 741.573
C0 DIODE VPWR 0.13fF
C1 DIODE VGND 0.13fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__dlclkp_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__dlclkp_1 GATE GCLK CLK VGND VPWR VNB VPB
X0 a_381_369.t0 GATE.t0 VPWR.t4 VPB.t5 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1 a_476_413.t1 a_193_47.t2 a_381_369.t1 VPB.t8 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 a_957_369.t1 a_642_307.t2 VPWR.t7 VPB.t9 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X3 VPWR.t5 CLK.t0 a_27_47.t1 VPB.t6 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X4 a_1042_47.t1 a_642_307.t3 a_957_369.t0 VNB.t6 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 GCLK.t1 a_957_369.t3 VPWR.t2 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 VGND.t1 CLK.t1 a_1042_47.t0 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7 a_193_47.t0 a_27_47.t2 VGND.t0 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 a_651_47.t0 a_193_47.t3 a_476_413.t0 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=390000u l=150000u
X9 a_193_47.t1 a_27_47.t3 VPWR.t3 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X10 GCLK.t0 a_957_369.t4 VGND.t5 VNB.t8 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 VPWR.t0 a_642_307.t4 a_600_413.t1 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12 a_476_413.t2 a_27_47.t4 a_396_119.t0 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13 VPWR.t6 CLK.t2 a_957_369.t2 VPB.t7 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X14 a_642_307.t0 a_476_413.t4 VGND.t4 VNB.t7 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X15 a_600_413.t0 a_27_47.t5 a_476_413.t3 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16 VPWR.t1 a_476_413.t5 a_642_307.t1 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17 VGND.t3 a_642_307.t5 a_651_47.t1 VNB.t5 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18 VGND.t2 CLK.t3 a_27_47.t0 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19 a_396_119.t1 GATE.t1 VGND.t6 VNB.t9 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
R0 GATE.n0 GATE.t1 189.586
R1 GATE.n0 GATE.t0 183.159
R2 GATE.n1 GATE.n0 76
R3  GATE.n1 59.264
R4 GATE.n1 GATE 12.288
R5 VPWR.n14 VPWR.t4 438.422
R6 VPWR.n6 VPWR.t0 373.741
R7 VPWR.n1 VPWR.n0 312.71
R8 VPWR.n19 VPWR.n18 311.893
R9 VPWR.n3 VPWR.n2 311.754
R10 VPWR.n2 VPWR.t6 58.484
R11 VPWR.n0 VPWR.t7 53.867
R12 VPWR.n18 VPWR.t3 41.554
R13 VPWR.n18 VPWR.t5 41.554
R14 VPWR.n0 VPWR.t1 36.222
R15 VPWR.n2 VPWR.t2 31.605
R16 VPWR.n5 VPWR.n4 4.65
R17 VPWR.n7 VPWR.n6 4.65
R18 VPWR.n9 VPWR.n8 4.65
R19 VPWR.n11 VPWR.n10 4.65
R20 VPWR.n13 VPWR.n12 4.65
R21 VPWR.n15 VPWR.n14 4.65
R22 VPWR.n17 VPWR.n16 4.65
R23 VPWR.n20 VPWR.n19 3.932
R24 VPWR.n3 VPWR.n1 3.803
R25 VPWR.n5 VPWR.n3 0.155
R26 VPWR.n20 VPWR.n17 0.137
R27 VPWR VPWR.n20 0.121
R28 VPWR.n7 VPWR.n5 0.119
R29 VPWR.n9 VPWR.n7 0.119
R30 VPWR.n11 VPWR.n9 0.119
R31 VPWR.n13 VPWR.n11 0.119
R32 VPWR.n15 VPWR.n13 0.119
R33 VPWR.n17 VPWR.n15 0.119
R34 a_381_369.t0 a_381_369.t1 132.285
R35 VPB.t3 VPB.t5 574.276
R36 VPB.t0 VPB.t1 562.305
R37 VPB.t9 VPB.t7 464.641
R38 VPB.t8 VPB.t4 372.972
R39 VPB.t5 VPB.t8 290.192
R40 VPB.t7 VPB.t2 281.152
R41 VPB.t1 VPB.t9 281.152
R42 VPB.t6 VPB.t3 256.591
R43 VPB.t4 VPB.t0 213.084
R44 VPB VPB.t6 198.552
R45 a_193_47.n0 a_193_47.t3 290.244
R46 a_193_47.n0 a_193_47.t2 234.881
R47 a_193_47.t1 a_193_47.n1 216.28
R48 a_193_47.n1 a_193_47.t0 204.248
R49 a_193_47.n1 a_193_47.n0 96.376
R50 a_476_413.n3 a_476_413.n2 434.713
R51 a_476_413.n1 a_476_413.t5 234.481
R52 a_476_413.n2 a_476_413.n0 180.544
R53 a_476_413.n1 a_476_413.t4 162.181
R54 a_476_413.n0 a_476_413.t2 152.793
R55 a_476_413.t1 a_476_413.n3 121.952
R56 a_476_413.n3 a_476_413.t3 98.5
R57 a_476_413.n2 a_476_413.n1 93.454
R58 a_476_413.n0 a_476_413.t0 46.154
R59 a_642_307.t1 a_642_307.n4 460.314
R60 a_642_307.n2 a_642_307.t5 370.701
R61 a_642_307.n0 a_642_307.t2 299.374
R62 a_642_307.n0 a_642_307.t3 292.948
R63 a_642_307.n2 a_642_307.t4 165.339
R64 a_642_307.n1 a_642_307.t0 152.029
R65 a_642_307.n3 a_642_307.n2 95.587
R66 a_642_307.n1 a_642_307.n0 76
R67 a_642_307.n4 a_642_307.n1 31.504
R68 a_642_307.n4 a_642_307.n3 0.193
R69 a_957_369.n0 a_957_369.t3 241.534
R70 a_957_369.n2 a_957_369.n1 233.057
R71 a_957_369.n1 a_957_369.t0 211.828
R72 a_957_369.n0 a_957_369.t4 169.234
R73 a_957_369.t1 a_957_369.n2 118.507
R74 a_957_369.n2 a_957_369.t2 76.953
R75 a_957_369.n1 a_957_369.n0 76
R76 CLK.n1 CLK.t0 259.402
R77 CLK.n0 CLK.t2 259.044
R78 CLK.n3 CLK.t3 230.191
R79 CLK.n0 CLK.t1 228.686
R80 CLK.n4 CLK.n0 17.062
R81 CLK.n2 CLK.n1 10.516
R82 CLK.n4 CLK.n3 8.764
R83 CLK CLK.n6 7.836
R84 CLK.n3 CLK.n2 4.381
R85 CLK.n6 CLK.n5 3.134
R86 CLK.n5 CLK.n4 1.306
R87 a_27_47.n0 a_27_47.t4 747.099
R88 a_27_47.t4 a_27_47.t5 660.339
R89 a_27_47.t1 a_27_47.n2 289.299
R90 a_27_47.n1 a_27_47.t3 266.384
R91 a_27_47.n2 a_27_47.t0 208.015
R92 a_27_47.n0 a_27_47.t2 91.58
R93 a_27_47.n1 a_27_47.n0 84.832
R94 a_27_47.n2 a_27_47.n1 76
R95 a_1042_47.t0 a_1042_47.t1 60
R96 VNB VNB.t3 6438.23
R97 VNB.t2 VNB.t9 5684.28
R98 VNB.t7 VNB.t6 5321.88
R99 VNB.t1 VNB.t0 4215.27
R100 VNB.t3 VNB.t2 2717.65
R101 VNB.t0 VNB.t5 2696.77
R102 VNB.t5 VNB.t7 2566.51
R103 VNB.t9 VNB.t1 2521.88
R104 VNB.t6 VNB.t4 2329.41
R105 VNB.t4 VNB.t8 2255.35
R106 GCLK.n0 GCLK.t1 538.75
R107 GCLK GCLK.t1 531.565
R108 GCLK GCLK.t0 157.328
R109 GCLK.n0 GCLK 77.492
R110 GCLK GCLK.n0 6.037
R111 VGND.n12 VGND.t6 172.631
R112 VGND.n3 VGND.n0 119.198
R113 VGND.n2 VGND.n1 117.417
R114 VGND.n17 VGND.n16 106.463
R115 VGND.n1 VGND.t3 70.329
R116 VGND.n0 VGND.t1 52.857
R117 VGND.n16 VGND.t0 38.571
R118 VGND.n16 VGND.t2 38.571
R119 VGND.n0 VGND.t5 27.362
R120 VGND.n1 VGND.t4 24.924
R121 VGND.n13 VGND.n12 4.65
R122 VGND.n15 VGND.n14 4.65
R123 VGND.n5 VGND.n4 4.65
R124 VGND.n7 VGND.n6 4.65
R125 VGND.n9 VGND.n8 4.65
R126 VGND.n11 VGND.n10 4.65
R127 VGND.n18 VGND.n17 3.932
R128 VGND.n3 VGND.n2 3.79
R129 VGND.n5 VGND.n3 0.144
R130 VGND.n18 VGND.n15 0.137
R131 VGND VGND.n18 0.121
R132 VGND.n7 VGND.n5 0.119
R133 VGND.n9 VGND.n7 0.119
R134 VGND.n11 VGND.n9 0.119
R135 VGND.n13 VGND.n11 0.119
R136 VGND.n15 VGND.n13 0.119
R137 a_651_47.t1 a_651_47.t0 88.152
R138 a_600_413.t0 a_600_413.t1 98.5
R139 a_396_119.t0 a_396_119.t1 121.299
R140 a_396_119.n0 a_396_119.t0 29.538
C0 GATE VGND 0.11fF
C1 CLK VGND 0.26fF
C2 CLK VPWR 0.19fF
C3 VPB VPWR 0.13fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__dlclkp_2.ext - technology: sky130A

.subckt sky130_fd_sc_hd__dlclkp_2 GATE GCLK CLK VGND VPWR VNB VPB
X0 a_381_369.t1 GATE.t0 VPWR.t8 VPB.t10 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1 a_957_369.t1 a_643_307.t2 VPWR.t2 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X2 a_601_413.t0 a_27_47.t2 a_477_413.t1 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3 a_397_119.t1 GATE.t1 VGND.t7 VNB.t10 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 VPWR.t3 CLK.t0 a_27_47.t0 VPB.t5 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X5 a_1041_47.t0 a_643_307.t3 a_957_369.t0 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 a_477_413.t0 a_193_47.t2 a_381_369.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7 VPWR.t5 a_957_369.t3 GCLK.t3 VPB.t7 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 GCLK.t2 a_957_369.t4 VPWR.t6 VPB.t8 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 VGND.t5 CLK.t1 a_1041_47.t1 VNB.t8 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10 a_193_47.t0 a_27_47.t3 VGND.t0 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11 a_652_47.t0 a_193_47.t3 a_477_413.t3 VNB.t5 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=390000u l=150000u
X12 VGND.t4 a_957_369.t5 GCLK.t1 VNB.t7 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 VPWR.t4 CLK.t2 a_957_369.t2 VPB.t6 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X14 a_193_47.t1 a_27_47.t4 VPWR.t0 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X15 GCLK.t0 a_957_369.t6 VGND.t3 VNB.t6 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X16 a_477_413.t2 a_27_47.t5 a_397_119.t0 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17 VPWR.t1 a_477_413.t4 a_643_307.t0 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X18 VGND.t1 a_643_307.t4 a_652_47.t1 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19 VPWR.t7 a_643_307.t5 a_601_413.t1 VPB.t9 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20 a_643_307.t1 a_477_413.t5 VGND.t2 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X21 VGND.t6 CLK.t3 a_27_47.t1 VNB.t9 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
R0 GATE.n0 GATE.t1 189.422
R1 GATE.n0 GATE.t0 183.694
R2 GATE.n1 GATE.n0 76
R3 GATE.n1 GATE 12.288
R4  GATE.n1 11.264
R5 VPWR.n20 VPWR.t8 438.422
R6 VPWR.n12 VPWR.t7 373.741
R7 VPWR.n8 VPWR.n7 312.71
R8 VPWR.n25 VPWR.n24 311.893
R9 VPWR.n1 VPWR.n0 308.042
R10 VPWR.n2 VPWR.t5 159.676
R11 VPWR.n0 VPWR.t4 60.023
R12 VPWR.n7 VPWR.t2 60.023
R13 VPWR.n24 VPWR.t0 41.554
R14 VPWR.n24 VPWR.t3 41.554
R15 VPWR.n0 VPWR.t6 31.605
R16 VPWR.n7 VPWR.t1 31.605
R17 VPWR.n4 VPWR.n3 4.65
R18 VPWR.n6 VPWR.n5 4.65
R19 VPWR.n9 VPWR.n8 4.65
R20 VPWR.n11 VPWR.n10 4.65
R21 VPWR.n13 VPWR.n12 4.65
R22 VPWR.n15 VPWR.n14 4.65
R23 VPWR.n17 VPWR.n16 4.65
R24 VPWR.n19 VPWR.n18 4.65
R25 VPWR.n21 VPWR.n20 4.65
R26 VPWR.n23 VPWR.n22 4.65
R27 VPWR.n26 VPWR.n25 3.932
R28 VPWR.n2 VPWR.n1 3.815
R29 VPWR.n4 VPWR.n2 0.24
R30 VPWR.n26 VPWR.n23 0.137
R31 VPWR VPWR.n26 0.121
R32 VPWR.n6 VPWR.n4 0.119
R33 VPWR.n9 VPWR.n6 0.119
R34 VPWR.n11 VPWR.n9 0.119
R35 VPWR.n13 VPWR.n11 0.119
R36 VPWR.n15 VPWR.n13 0.119
R37 VPWR.n17 VPWR.n15 0.119
R38 VPWR.n19 VPWR.n17 0.119
R39 VPWR.n21 VPWR.n19 0.119
R40 VPWR.n23 VPWR.n21 0.119
R41 a_381_369.t1 a_381_369.t0 134.63
R42 VPB.t1 VPB.t10 574.276
R43 VPB.t9 VPB.t2 556.386
R44 VPB.t4 VPB.t6 461.682
R45 VPB.t0 VPB.t3 372.972
R46 VPB.t10 VPB.t0 293.247
R47 VPB.t6 VPB.t8 284.112
R48 VPB.t2 VPB.t4 284.112
R49 VPB.t5 VPB.t1 256.591
R50 VPB.t8 VPB.t7 248.598
R51 VPB.t3 VPB.t9 213.084
R52 VPB VPB.t5 195.498
R53 a_643_307.t0 a_643_307.n4 466.769
R54 a_643_307.n3 a_643_307.t4 370.701
R55 a_643_307.n0 a_643_307.t2 299.374
R56 a_643_307.n0 a_643_307.t3 292.948
R57 a_643_307.n3 a_643_307.t5 165.339
R58 a_643_307.n1 a_643_307.t1 151.427
R59 a_643_307.n4 a_643_307.n3 95.393
R60 a_643_307.n1 a_643_307.n0 76
R61 a_643_307.n2 a_643_307.n1 30.742
R62 a_643_307.n4 a_643_307.n2 0.193
R63 a_957_369.n3 a_957_369.n2 233.409
R64 a_957_369.n2 a_957_369.t0 213.241
R65 a_957_369.n0 a_957_369.t3 212.079
R66 a_957_369.n1 a_957_369.t4 212.079
R67 a_957_369.n0 a_957_369.t5 139.779
R68 a_957_369.n1 a_957_369.t6 139.779
R69 a_957_369.t1 a_957_369.n3 120.046
R70 a_957_369.n2 a_957_369.n1 84.763
R71 a_957_369.n3 a_957_369.t2 73.875
R72 a_957_369.n1 a_957_369.n0 61.345
R73 a_27_47.n0 a_27_47.t5 748.705
R74 a_27_47.t5 a_27_47.t2 660.339
R75 a_27_47.t0 a_27_47.n2 289.299
R76 a_27_47.n1 a_27_47.t4 266.384
R77 a_27_47.n2 a_27_47.t1 208.015
R78 a_27_47.n0 a_27_47.t3 91.58
R79 a_27_47.n1 a_27_47.n0 84.832
R80 a_27_47.n2 a_27_47.n1 76
R81 a_477_413.n3 a_477_413.n2 434.336
R82 a_477_413.n1 a_477_413.t4 235.131
R83 a_477_413.n2 a_477_413.n0 180.168
R84 a_477_413.n1 a_477_413.t5 162.831
R85 a_477_413.n0 a_477_413.t2 152.793
R86 a_477_413.t0 a_477_413.n3 121.952
R87 a_477_413.n3 a_477_413.t1 98.5
R88 a_477_413.n2 a_477_413.n1 93.648
R89 a_477_413.n0 a_477_413.t3 46.154
R90 a_601_413.t0 a_601_413.t1 98.5
R91 VGND.n22 VGND.t7 174.06
R92 VGND.n12 VGND.n11 117.045
R93 VGND.n2 VGND.n1 114.711
R94 VGND.n27 VGND.n26 106.463
R95 VGND.n0 VGND.t4 101.097
R96 VGND.n11 VGND.t1 67.978
R97 VGND.n1 VGND.t5 55.714
R98 VGND.n26 VGND.t0 38.571
R99 VGND.n26 VGND.t6 38.571
R100 VGND.n1 VGND.t3 25.934
R101 VGND.n11 VGND.t2 24.923
R102 VGND.n23 VGND.n22 4.65
R103 VGND.n25 VGND.n24 4.65
R104 VGND.n4 VGND.n3 4.65
R105 VGND.n6 VGND.n5 4.65
R106 VGND.n8 VGND.n7 4.65
R107 VGND.n10 VGND.n9 4.65
R108 VGND.n13 VGND.n12 4.65
R109 VGND.n15 VGND.n14 4.65
R110 VGND.n17 VGND.n16 4.65
R111 VGND.n19 VGND.n18 4.65
R112 VGND.n21 VGND.n20 4.65
R113 VGND.n28 VGND.n27 3.932
R114 VGND.n4 VGND.n0 0.781
R115 VGND.n3 VGND.n2 0.752
R116 VGND.n28 VGND.n25 0.137
R117 VGND VGND.n28 0.121
R118 VGND.n6 VGND.n4 0.119
R119 VGND.n8 VGND.n6 0.119
R120 VGND.n10 VGND.n8 0.119
R121 VGND.n13 VGND.n10 0.119
R122 VGND.n15 VGND.n13 0.119
R123 VGND.n17 VGND.n15 0.119
R124 VGND.n19 VGND.n17 0.119
R125 VGND.n21 VGND.n19 0.119
R126 VGND.n23 VGND.n21 0.119
R127 VGND.n25 VGND.n23 0.119
R128 a_397_119.t0 a_397_119.t1 121.299
R129 a_397_119.n0 a_397_119.t0 29.538
R130 VNB VNB.t9 6438.23
R131 VNB.t1 VNB.t10 5707.56
R132 VNB.t4 VNB.t3 5321.88
R133 VNB.t0 VNB.t5 4215.27
R134 VNB.t9 VNB.t1 2717.65
R135 VNB.t5 VNB.t2 2696.77
R136 VNB.t10 VNB.t0 2521.88
R137 VNB.t2 VNB.t4 2518.16
R138 VNB.t3 VNB.t8 2329.41
R139 VNB.t8 VNB.t6 2269.18
R140 VNB.t6 VNB.t7 2030.77
R141 CLK.n1 CLK.t0 259.743
R142 CLK.n0 CLK.t2 259.044
R143 CLK.n3 CLK.t3 230.645
R144 CLK.n0 CLK.t1 228.686
R145 CLK.n4 CLK.n0 16.975
R146 CLK.n2 CLK.n1 10.711
R147 CLK.n4 CLK.n3 8.764
R148 CLK CLK.n6 8
R149 CLK.n3 CLK.n2 4.462
R150 CLK.n6 CLK.n5 3.2
R151 CLK.n5 CLK.n4 1.333
R152 a_1041_47.t0 a_1041_47.t1 60
R153 a_193_47.n0 a_193_47.t3 275.728
R154 a_193_47.n0 a_193_47.t2 234.881
R155 a_193_47.t1 a_193_47.n1 216.28
R156 a_193_47.n1 a_193_47.t0 204.248
R157 a_193_47.n1 a_193_47.n0 94.192
R158 GCLK GCLK.n0 300.469
R159 GCLK.n2 GCLK.n0 292.5
R160 GCLK GCLK.n1 92.713
R161 GCLK.n2 GCLK 74.298
R162 GCLK.n0 GCLK.t3 26.595
R163 GCLK.n0 GCLK.t2 26.595
R164 GCLK.n1 GCLK.t1 24.923
R165 GCLK.n1 GCLK.t0 24.923
R166 GCLK GCLK.n2 6.037
R167 a_652_47.t1 a_652_47.t0 88.152
C0 VGND GCLK 0.17fF
C1 VPWR GCLK 0.23fF
C2 GATE VGND 0.14fF
C3 CLK VGND 0.26fF
C4 CLK VPWR 0.19fF
C5 VPB VPWR 0.15fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__dlclkp_4.ext - technology: sky130A

.subckt sky130_fd_sc_hd__dlclkp_4 CLK GCLK GATE VPWR VGND VNB VPB
X0 a_575_47.t1 a_193_47.t2 a_477_413.t3 VNB.t12 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X1 a_381_369.t0 GATE.t0 VPWR.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X2 a_1046_47.t0 a_627_153.t2 a_953_297.t0 VNB.t9 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 a_953_297.t1 a_627_153.t3 VPWR.t9 VPB.t10 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 VPWR.t4 a_953_297.t3 GCLK.t7 VPB.t5 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 GCLK.t3 a_953_297.t4 VGND.t9 VNB.t7 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 VPWR.t10 a_627_153.t4 a_585_413.t0 VPB.t11 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7 GCLK.t6 a_953_297.t5 VPWR.t5 VPB.t6 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 VPWR.t1 CLK.t0 a_27_47.t1 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X9 VPWR.t2 CLK.t1 a_953_297.t2 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 GCLK.t5 a_953_297.t6 VPWR.t6 VPB.t7 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 a_477_413.t2 a_193_47.t3 a_381_369.t1 VPB.t12 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12 VPWR.t7 a_953_297.t7 GCLK.t4 VPB.t8 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13 a_585_413.t1 a_27_47.t2 a_477_413.t0 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14 a_477_413.t1 a_27_47.t3 a_381_47.t1 VNB.t5 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X15 VPWR.t8 a_477_413.t4 a_627_153.t1 VPB.t9 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16 a_193_47.t0 a_27_47.t4 VGND.t4 VNB.t6 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17 GCLK.t2 a_953_297.t8 VGND.t8 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X18 a_193_47.t1 a_27_47.t5 VPWR.t3 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X19 VGND.t5 a_477_413.t5 a_627_153.t0 VNB.t8 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X20 VGND.t7 a_953_297.t9 GCLK.t1 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X21 VGND.t6 a_953_297.t10 GCLK.t0 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X22 a_381_47.t0 GATE.t1 VGND.t0 VNB.t11 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23 VGND.t2 CLK.t2 a_1046_47.t1 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X24 VGND.t1 a_627_153.t5 a_575_47.t0 VNB.t10 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X25 VGND.t3 CLK.t3 a_27_47.t0 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
R0 a_193_47.n0 a_193_47.t2 435.762
R1 a_193_47.t1 a_193_47.n1 242.337
R2 a_193_47.n0 a_193_47.t3 219.041
R3 a_193_47.n1 a_193_47.t0 177.44
R4 a_193_47.n1 a_193_47.n0 126.524
R5 a_477_413.n3 a_477_413.n2 412.318
R6 a_477_413.n0 a_477_413.t4 212.079
R7 a_477_413.n2 a_477_413.n1 188.499
R8 a_477_413.n2 a_477_413.n0 171.241
R9 a_477_413.n0 a_477_413.t5 143.43
R10 a_477_413.n3 a_477_413.t2 119.607
R11 a_477_413.t0 a_477_413.n3 63.321
R12 a_477_413.n1 a_477_413.t3 48.333
R13 a_477_413.n1 a_477_413.t1 46.666
R14 a_575_47.t0 a_575_47.t1 93.059
R15 VNB VNB.t4 6438.23
R16 VNB.t6 VNB.t11 6082.35
R17 VNB.t10 VNB.t8 5321.88
R18 VNB.t8 VNB.t9 4545.05
R19 VNB.t11 VNB.t5 3461.76
R20 VNB.t12 VNB.t10 3073.53
R21 VNB.t5 VNB.t12 2814.71
R22 VNB.t4 VNB.t6 2717.65
R23 VNB.t7 VNB.t1 2465.93
R24 VNB.t0 VNB.t2 2030.77
R25 VNB.t1 VNB.t0 2030.77
R26 VNB.t3 VNB.t7 2030.77
R27 VNB.t9 VNB.t3 2030.77
R28 GATE.n0 GATE.t1 800.12
R29 GATE.n0 GATE.t0 367.926
R30 GATE GATE.n0 89.056
R31 VPWR.n26 VPWR.t0 438.422
R32 VPWR.n18 VPWR.t10 369.332
R33 VPWR.n14 VPWR.n13 312.71
R34 VPWR.n31 VPWR.n0 311.893
R35 VPWR.n2 VPWR.n1 311.207
R36 VPWR.n7 VPWR.n6 168.598
R37 VPWR.n3 VPWR.t4 155.241
R38 VPWR.n0 VPWR.t3 41.554
R39 VPWR.n0 VPWR.t1 41.554
R40 VPWR.n13 VPWR.t9 39.4
R41 VPWR.n6 VPWR.t6 32.505
R42 VPWR.n6 VPWR.t2 32.505
R43 VPWR.n13 VPWR.t8 29.55
R44 VPWR.n1 VPWR.t5 26.595
R45 VPWR.n1 VPWR.t7 26.595
R46 VPWR.n32 VPWR.n31 26.108
R47 VPWR.n31 VPWR.n30 4.65
R48 VPWR.n5 VPWR.n4 4.65
R49 VPWR.n8 VPWR.n7 4.65
R50 VPWR.n10 VPWR.n9 4.65
R51 VPWR.n12 VPWR.n11 4.65
R52 VPWR.n15 VPWR.n14 4.65
R53 VPWR.n17 VPWR.n16 4.65
R54 VPWR.n19 VPWR.n18 4.65
R55 VPWR.n21 VPWR.n20 4.65
R56 VPWR.n23 VPWR.n22 4.65
R57 VPWR.n25 VPWR.n24 4.65
R58 VPWR.n27 VPWR.n26 4.65
R59 VPWR.n29 VPWR.n28 4.65
R60 VPWR.n3 VPWR.n2 3.904
R61 VPWR.n5 VPWR.n3 0.224
R62 VPWR.n8 VPWR.n5 0.119
R63 VPWR.n10 VPWR.n8 0.119
R64 VPWR.n12 VPWR.n10 0.119
R65 VPWR.n15 VPWR.n12 0.119
R66 VPWR.n17 VPWR.n15 0.119
R67 VPWR.n19 VPWR.n17 0.119
R68 VPWR.n21 VPWR.n19 0.119
R69 VPWR.n23 VPWR.n21 0.119
R70 VPWR.n25 VPWR.n23 0.119
R71 VPWR.n27 VPWR.n25 0.119
R72 VPWR.n29 VPWR.n27 0.119
R73 VPWR.n30 VPWR.n29 0.119
R74 VPWR.n30 VPWR 0.118
R75 VPWR VPWR.n32 0.02
R76 VPWR.n32 VPWR 0.001
R77 a_381_369.t0 a_381_369.t1 134.63
R78 VPB.t11 VPB.t9 580.062
R79 VPB.t4 VPB.t0 556.386
R80 VPB.t10 VPB.t2 488.317
R81 VPB.t12 VPB.t3 319.626
R82 VPB.t7 VPB.t8 301.869
R83 VPB.t9 VPB.t10 295.95
R84 VPB.t2 VPB.t7 284.112
R85 VPB.t0 VPB.t12 284.112
R86 VPB.t6 VPB.t5 248.598
R87 VPB.t8 VPB.t6 248.598
R88 VPB.t1 VPB.t4 248.598
R89 VPB.t3 VPB.t11 213.084
R90 VPB VPB.t1 189.408
R91 a_627_153.t1 a_627_153.n4 466.769
R92 a_627_153.n3 a_627_153.t5 353.754
R93 a_627_153.n0 a_627_153.t2 291.116
R94 a_627_153.n0 a_627_153.t3 263.388
R95 a_627_153.n3 a_627_153.t4 149.821
R96 a_627_153.n1 a_627_153.t0 145.846
R97 a_627_153.n1 a_627_153.n0 99.466
R98 a_627_153.n4 a_627_153.n3 96.945
R99 a_627_153.n2 a_627_153.n1 16.78
R100 a_627_153.n4 a_627_153.n2 0.969
R101 a_953_297.n0 a_953_297.t3 212.079
R102 a_953_297.n1 a_953_297.t5 212.079
R103 a_953_297.n2 a_953_297.t7 212.079
R104 a_953_297.n3 a_953_297.t6 212.079
R105 a_953_297.n5 a_953_297.t0 162.54
R106 a_953_297.n0 a_953_297.t10 139.779
R107 a_953_297.n1 a_953_297.t8 139.779
R108 a_953_297.n2 a_953_297.t9 139.779
R109 a_953_297.n3 a_953_297.t4 139.779
R110 a_953_297.n6 a_953_297.n5 129.171
R111 a_953_297.n6 a_953_297.t2 96.53
R112 a_953_297.n5 a_953_297.n4 67.003
R113 a_953_297.n1 a_953_297.n0 61.345
R114 a_953_297.n2 a_953_297.n1 61.345
R115 a_953_297.t1 a_953_297.n6 36.445
R116 a_953_297.n4 a_953_297.n2 34.464
R117 a_953_297.n4 a_953_297.n3 28.826
R118 a_1046_47.t0 a_1046_47.t1 49.846
R119 GCLK GCLK.n1 298.9
R120 GCLK.n5 GCLK.n4 292.5
R121 GCLK.n4 GCLK.n3 147.123
R122 GCLK.n6 GCLK.n0 141.038
R123 GCLK GCLK.n7 50.358
R124 GCLK.n1 GCLK.t4 44.325
R125 GCLK.n0 GCLK.t1 41.538
R126 GCLK.n1 GCLK.t5 26.595
R127 GCLK.n4 GCLK.t7 26.595
R128 GCLK.n4 GCLK.t6 26.595
R129 GCLK.n0 GCLK.t3 24.923
R130 GCLK.n7 GCLK.t0 24.923
R131 GCLK.n7 GCLK.t2 24.923
R132 GCLK.n2 GCLK 9.6
R133 GCLK.n6 GCLK 7.098
R134 GCLK GCLK.n5 5.003
R135 GCLK.n3 GCLK.n2 4.776
R136 GCLK.n5 GCLK 2.909
R137 GCLK.n2 GCLK 2.56
R138 GCLK.n3 GCLK 2.4
R139 GCLK GCLK.n6 0.814
R140 VGND.n19 VGND.t1 148.073
R141 VGND.n27 VGND.t0 145.59
R142 VGND.n15 VGND.t5 137.633
R143 VGND.n3 VGND.n2 114.711
R144 VGND.n1 VGND.t6 111.393
R145 VGND.n9 VGND.n8 109.871
R146 VGND.n32 VGND.n0 107.239
R147 VGND.n0 VGND.t4 38.571
R148 VGND.n0 VGND.t3 38.571
R149 VGND.n33 VGND.n32 26.108
R150 VGND.n2 VGND.t8 24.923
R151 VGND.n2 VGND.t7 24.923
R152 VGND.n8 VGND.t9 24.923
R153 VGND.n8 VGND.t2 24.923
R154 VGND.n32 VGND.n31 4.65
R155 VGND.n5 VGND.n4 4.65
R156 VGND.n7 VGND.n6 4.65
R157 VGND.n10 VGND.n9 4.65
R158 VGND.n12 VGND.n11 4.65
R159 VGND.n14 VGND.n13 4.65
R160 VGND.n16 VGND.n15 4.65
R161 VGND.n18 VGND.n17 4.65
R162 VGND.n20 VGND.n19 4.65
R163 VGND.n22 VGND.n21 4.65
R164 VGND.n24 VGND.n23 4.65
R165 VGND.n26 VGND.n25 4.65
R166 VGND.n28 VGND.n27 4.65
R167 VGND.n30 VGND.n29 4.65
R168 VGND.n4 VGND.n3 3.388
R169 VGND.n5 VGND.n1 0.753
R170 VGND.n7 VGND.n5 0.119
R171 VGND.n10 VGND.n7 0.119
R172 VGND.n12 VGND.n10 0.119
R173 VGND.n14 VGND.n12 0.119
R174 VGND.n16 VGND.n14 0.119
R175 VGND.n18 VGND.n16 0.119
R176 VGND.n20 VGND.n18 0.119
R177 VGND.n22 VGND.n20 0.119
R178 VGND.n24 VGND.n22 0.119
R179 VGND.n26 VGND.n24 0.119
R180 VGND.n28 VGND.n26 0.119
R181 VGND.n30 VGND.n28 0.119
R182 VGND.n31 VGND.n30 0.119
R183 VGND.n31 VGND 0.118
R184 VGND VGND.n33 0.02
R185 VGND.n33 VGND 0.001
R186 a_585_413.t0 a_585_413.t1 98.5
R187 CLK.n3 CLK.t0 259.402
R188 CLK.n0 CLK.t1 241.534
R189 CLK.n5 CLK.t3 230.191
R190 CLK.n0 CLK.t2 169.234
R191 CLK.n7 CLK.n0 99.052
R192 CLK.n4 CLK.n3 10.516
R193 CLK.n6 CLK.n5 8.764
R194 CLK.n1 CLK 8
R195 CLK.n5 CLK.n4 4.381
R196 CLK CLK.n7 3.42
R197 CLK.n2 CLK.n1 3.2
R198 CLK.n6 CLK.n2 1.333
R199 CLK.n7 CLK.n6 1.061
R200 a_27_47.n0 a_27_47.t5 263.171
R201 a_27_47.n2 a_27_47.t3 258.418
R202 a_27_47.t1 a_27_47.n3 245.105
R203 a_27_47.n0 a_27_47.t4 227.825
R204 a_27_47.n2 a_27_47.t2 225.22
R205 a_27_47.n1 a_27_47.t0 196.895
R206 a_27_47.n3 a_27_47.n2 88.532
R207 a_27_47.n1 a_27_47.n0 76
R208 a_27_47.n3 a_27_47.n1 38.923
R209 a_381_47.n0 a_381_47.t1 86.666
R210 a_381_47.n0 a_381_47.t0 26.393
R211 a_381_47.n1 a_381_47.n0 14.4
C0 VGND CLK 0.26fF
C1 VPWR CLK 0.16fF
C2 VPWR VPB 0.17fF
C3 VGND GCLK 0.42fF
C4 VPWR GCLK 0.51fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__dlrbn_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__dlrbn_1 RESET_B Q_N Q D GATE_N VGND VPWR VNB VPB
X0 Q.t0 a_724_21.t3 VGND.t4 VNB.t6 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 VPWR.t8 D.t0 a_299_47.t1 VPB.t9 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X2 a_561_413.t3 a_27_47.t2 a_465_47.t1 VNB.t10 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X3 a_465_47.t0 a_299_47.t2 VGND.t0 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 Q.t1 a_724_21.t4 VPWR.t1 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 a_561_413.t0 a_193_47.t2 a_465_369.t1 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 a_724_21.t0 a_561_413.t4 VPWR.t0 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 VGND.t2 a_724_21.t5 a_659_47.t0 VNB.t5 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 VPWR.t4 GATE_N.t0 a_27_47.t0 VPB.t5 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X9 Q_N.t1 a_1308_47.t2 VPWR.t5 VPB.t6 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 a_659_47.t1 a_193_47.t3 a_561_413.t1 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X11 VPWR.t3 a_724_21.t6 a_682_413.t0 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12 VGND.t3 a_724_21.t7 a_1308_47.t0 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13 a_193_47.t0 a_27_47.t3 VGND.t8 VNB.t11 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14 a_682_413.t1 a_27_47.t4 a_561_413.t2 VPB.t10 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15 VPWR.t7 RESET_B.t0 a_724_21.t2 VPB.t8 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16 a_942_47.t1 a_561_413.t5 a_724_21.t1 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X17 VPWR.t2 a_724_21.t8 a_1308_47.t1 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X18 a_193_47.t1 a_27_47.t5 VPWR.t9 VPB.t11 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X19 Q_N.t0 a_1308_47.t3 VGND.t6 VNB.t8 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X20 VGND.t1 D.t1 a_299_47.t0 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21 VGND.t7 RESET_B.t1 a_942_47.t0 VNB.t9 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X22 a_465_369.t0 a_299_47.t3 VPWR.t6 VPB.t7 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X23 VGND.t5 GATE_N.t1 a_27_47.t1 VNB.t7 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
R0 a_724_21.n3 a_724_21.t5 368.328
R1 a_724_21.n0 a_724_21.t8 247.54
R2 a_724_21.n2 a_724_21.t1 228.301
R3 a_724_21.n1 a_724_21.t4 212.079
R4 a_724_21.n0 a_724_21.t7 154.354
R5 a_724_21.n5 a_724_21.n4 151.979
R6 a_724_21.n3 a_724_21.t6 149.821
R7 a_724_21.n1 a_724_21.t3 139.779
R8 a_724_21.n1 a_724_21.n0 118.309
R9 a_724_21.n4 a_724_21.n3 112.864
R10 a_724_21.n2 a_724_21.n1 97.178
R11 a_724_21.n4 a_724_21.n2 65.208
R12 a_724_21.t0 a_724_21.n5 34.475
R13 a_724_21.n5 a_724_21.t2 26.595
R14 VGND.n13 VGND.t2 148.331
R15 VGND.n4 VGND.n1 110.989
R16 VGND.n29 VGND.n0 107.239
R17 VGND.n22 VGND.n21 106.463
R18 VGND.n3 VGND.n2 92.5
R19 VGND.n6 VGND.n5 92.5
R20 VGND.n1 VGND.t3 54.285
R21 VGND.n21 VGND.t0 38.571
R22 VGND.n21 VGND.t1 38.571
R23 VGND.n0 VGND.t8 38.571
R24 VGND.n0 VGND.t5 38.571
R25 VGND.n5 VGND.t7 35.076
R26 VGND.n2 VGND.t4 27.692
R27 VGND.n30 VGND.n29 26.108
R28 VGND.n1 VGND.t6 25.934
R29 VGND.n4 VGND.n3 4.939
R30 VGND.n29 VGND.n28 4.65
R31 VGND.n8 VGND.n7 4.65
R32 VGND.n10 VGND.n9 4.65
R33 VGND.n12 VGND.n11 4.65
R34 VGND.n14 VGND.n13 4.65
R35 VGND.n16 VGND.n15 4.65
R36 VGND.n18 VGND.n17 4.65
R37 VGND.n20 VGND.n19 4.65
R38 VGND.n23 VGND.n22 4.65
R39 VGND.n25 VGND.n24 4.65
R40 VGND.n27 VGND.n26 4.65
R41 VGND.n7 VGND.n6 1.571
R42 VGND.n8 VGND.n4 0.144
R43 VGND.n10 VGND.n8 0.119
R44 VGND.n12 VGND.n10 0.119
R45 VGND.n14 VGND.n12 0.119
R46 VGND.n16 VGND.n14 0.119
R47 VGND.n18 VGND.n16 0.119
R48 VGND.n20 VGND.n18 0.119
R49 VGND.n23 VGND.n20 0.119
R50 VGND.n25 VGND.n23 0.119
R51 VGND.n27 VGND.n25 0.119
R52 VGND.n28 VGND.n27 0.119
R53 VGND.n28 VGND 0.118
R54 VGND VGND.n30 0.02
R55 VGND.n30 VGND 0.001
R56 Q.n0 Q.t1 172.943
R57 Q.n1 Q.t0 117.423
R58 Q Q.n0 10.226
R59 Q Q.n1 10.2
R60 Q.n1 Q 3.4
R61 Q.n0 Q 3.303
R62 VNB.t11 VNB.t3 6082.35
R63 VNB.t5 VNB.t2 5321.88
R64 VNB.t6 VNB.t4 4545.05
R65 VNB VNB.t7 4238.23
R66 VNB.t9 VNB.t6 4061.54
R67 VNB.t0 VNB.t10 3494.12
R68 VNB.t1 VNB.t5 3073.53
R69 VNB.t10 VNB.t1 2782.35
R70 VNB.t3 VNB.t0 2717.65
R71 VNB.t7 VNB.t11 2717.65
R72 VNB.t4 VNB.t8 2296.7
R73 VNB.t2 VNB.t9 2224.18
R74 D.n0 D.t0 327.642
R75 D.n0 D.t1 157.336
R76 D D.n0 78.594
R77 a_299_47.n0 a_299_47.t3 373.281
R78 a_299_47.t1 a_299_47.n1 292.715
R79 a_299_47.n1 a_299_47.t0 182.645
R80 a_299_47.n0 a_299_47.t2 132.281
R81 a_299_47.n1 a_299_47.n0 80.46
R82 VPWR.n8 VPWR.t0 576.219
R83 VPWR.n10 VPWR.t3 375.732
R84 VPWR.n26 VPWR.n0 311.893
R85 VPWR.n3 VPWR.n2 170.129
R86 VPWR.n19 VPWR.n18 165.066
R87 VPWR.n1 VPWR.t7 75.845
R88 VPWR.n1 VPWR.t1 60.085
R89 VPWR.n2 VPWR.t2 58.484
R90 VPWR.n18 VPWR.t6 41.554
R91 VPWR.n18 VPWR.t8 41.554
R92 VPWR.n0 VPWR.t9 41.554
R93 VPWR.n0 VPWR.t4 41.554
R94 VPWR.n2 VPWR.t5 31.605
R95 VPWR.n27 VPWR.n26 26.108
R96 VPWR.n3 VPWR.n1 6.877
R97 VPWR.n26 VPWR.n25 4.65
R98 VPWR.n5 VPWR.n4 4.65
R99 VPWR.n7 VPWR.n6 4.65
R100 VPWR.n9 VPWR.n8 4.65
R101 VPWR.n11 VPWR.n10 4.65
R102 VPWR.n13 VPWR.n12 4.65
R103 VPWR.n15 VPWR.n14 4.65
R104 VPWR.n17 VPWR.n16 4.65
R105 VPWR.n20 VPWR.n19 4.65
R106 VPWR.n22 VPWR.n21 4.65
R107 VPWR.n24 VPWR.n23 4.65
R108 VPWR.n5 VPWR.n3 0.145
R109 VPWR.n7 VPWR.n5 0.119
R110 VPWR.n9 VPWR.n7 0.119
R111 VPWR.n11 VPWR.n9 0.119
R112 VPWR.n13 VPWR.n11 0.119
R113 VPWR.n15 VPWR.n13 0.119
R114 VPWR.n17 VPWR.n15 0.119
R115 VPWR.n20 VPWR.n17 0.119
R116 VPWR.n22 VPWR.n20 0.119
R117 VPWR.n24 VPWR.n22 0.119
R118 VPWR.n25 VPWR.n24 0.119
R119 VPWR.n25 VPWR 0.118
R120 VPWR VPWR.n27 0.02
R121 VPWR.n27 VPWR 0.001
R122 VPB.t4 VPB.t2 556.386
R123 VPB.t3 VPB.t1 556.386
R124 VPB.t11 VPB.t9 556.386
R125 VPB.t8 VPB.t4 497.196
R126 VPB.t0 VPB.t10 358.099
R127 VPB.t7 VPB.t0 284.112
R128 VPB.t2 VPB.t6 281.152
R129 VPB.t1 VPB.t8 272.274
R130 VPB.t9 VPB.t7 248.598
R131 VPB.t5 VPB.t11 248.598
R132 VPB.t10 VPB.t3 213.084
R133 VPB VPB.t5 139.096
R134 a_27_47.t0 a_27_47.n3 265.057
R135 a_27_47.n1 a_27_47.t5 263.171
R136 a_27_47.n0 a_27_47.t4 240.108
R137 a_27_47.n0 a_27_47.t2 239.726
R138 a_27_47.n1 a_27_47.t3 227.825
R139 a_27_47.n2 a_27_47.t1 196.895
R140 a_27_47.n2 a_27_47.n1 76
R141 a_27_47.n3 a_27_47.n2 18.97
R142 a_27_47.n3 a_27_47.n0 11.268
R143 a_465_47.n0 a_465_47.t1 88.333
R144 a_465_47.n0 a_465_47.t0 26.393
R145 a_465_47.n1 a_465_47.n0 14.4
R146 a_561_413.n3 a_561_413.n2 400.17
R147 a_561_413.n0 a_561_413.t4 212.079
R148 a_561_413.n2 a_561_413.n0 171.139
R149 a_561_413.n2 a_561_413.n1 166.462
R150 a_561_413.n0 a_561_413.t5 139.779
R151 a_561_413.t0 a_561_413.n3 121.952
R152 a_561_413.n3 a_561_413.t2 91.464
R153 a_561_413.n1 a_561_413.t1 46.666
R154 a_561_413.n1 a_561_413.t3 46.666
R155 a_193_47.n0 a_193_47.t3 464.325
R156 a_193_47.n0 a_193_47.t2 242.606
R157 a_193_47.n1 a_193_47.t0 230.004
R158 a_193_47.t1 a_193_47.n1 121.759
R159 a_193_47.n1 a_193_47.n0 99.063
R160 a_465_369.t0 a_465_369.t1 134.63
R161 a_659_47.t0 a_659_47.t1 93.059
R162 GATE_N.n0 GATE_N.t0 269.919
R163 GATE_N.n0 GATE_N.t1 234.573
R164 GATE_N.n1 GATE_N.n0 76
R165 GATE_N GATE_N.n1 10.971
R166 GATE_N.n1 GATE_N 6.791
R167 a_1308_47.t1 a_1308_47.n1 377.062
R168 a_1308_47.n0 a_1308_47.t2 237.733
R169 a_1308_47.n1 a_1308_47.t0 218.035
R170 a_1308_47.n0 a_1308_47.t3 165.433
R171 a_1308_47.n1 a_1308_47.n0 99.272
R172 Q_N.n1 Q_N.t1 172.965
R173 Q_N.n0 Q_N.t0 117.423
R174 Q_N Q_N.n0 95.163
R175 Q_N.n1 Q_N 12.564
R176 Q_N Q_N.n1 4.065
R177 Q_N.n0 Q_N 0.246
R178 a_682_413.t0 a_682_413.t1 98.5
R179 RESET_B.n0 RESET_B.t0 241.534
R180 RESET_B.n0 RESET_B.t1 169.234
R181 RESET_B.n1 RESET_B.n0 76
R182 RESET_B.n1 RESET_B 10.278
R183 RESET_B RESET_B.n1 7.563
R184 a_942_47.t0 a_942_47.t1 57.23
C0 VPWR Q_N 0.12fF
C1 VPWR Q 0.15fF
C2 VPWR VGND 0.14fF
C3 VPB VPWR 0.16fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__dlrbn_2.ext - technology: sky130A

.subckt sky130_fd_sc_hd__dlrbn_2 D GATE_N Q RESET_B Q_N VPWR VGND VNB VPB
X0 VPWR.t4 D.t0 a_299_47.t1 VPB.t5 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1 a_561_413.t1 a_27_47.t2 a_465_47.t0 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X2 a_465_47.t1 a_299_47.t2 VGND.t1 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3 Q_N.t1 a_1313_47.t2 VPWR.t10 VPB.t12 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 Q_N.t3 a_1313_47.t3 VGND.t10 VNB.t13 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 a_561_413.t2 a_193_47.t2 a_465_369.t1 VPB.t6 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 a_724_21.t1 a_561_413.t4 VPWR.t2 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 VGND.t6 a_724_21.t3 a_659_47.t0 VNB.t9 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 VPWR.t5 GATE_N.t0 a_27_47.t0 VPB.t7 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X9 VPWR.t11 a_1313_47.t4 Q_N.t0 VPB.t13 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 VGND.t7 a_724_21.t4 a_1313_47.t0 VNB.t10 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11 a_659_47.t1 a_193_47.t3 a_561_413.t3 VNB.t6 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X12 VPWR.t6 a_724_21.t5 a_682_413.t1 VPB.t8 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13 VGND.t5 a_1313_47.t5 Q_N.t2 VNB.t8 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14 a_193_47.t1 a_27_47.t3 VGND.t0 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15 a_682_413.t0 a_27_47.t4 a_561_413.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16 Q.t3 a_724_21.t6 VGND.t8 VNB.t11 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X17 a_942_47.t0 a_561_413.t5 a_724_21.t0 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X18 VPWR.t7 a_724_21.t7 a_1313_47.t1 VPB.t9 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X19 VPWR.t8 a_724_21.t8 Q.t1 VPB.t10 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X20 a_193_47.t0 a_27_47.t5 VPWR.t0 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X21 Q.t0 a_724_21.t9 VPWR.t9 VPB.t11 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X22 VPWR.t3 RESET_B.t0 a_724_21.t2 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X23 VGND.t3 D.t1 a_299_47.t0 VNB.t5 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24 VGND.t2 RESET_B.t1 a_942_47.t1 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X25 VGND.t9 a_724_21.t10 Q.t2 VNB.t12 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X26 a_465_369.t0 a_299_47.t3 VPWR.t1 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X27 VGND.t4 GATE_N.t1 a_27_47.t1 VNB.t7 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
R0 D.n0 D.t0 327.642
R1 D.n0 D.t1 157.336
R2 D D.n0 78.594
R3 a_299_47.n0 a_299_47.t3 373.281
R4 a_299_47.t1 a_299_47.n1 292.715
R5 a_299_47.n1 a_299_47.t0 182.645
R6 a_299_47.n0 a_299_47.t2 132.281
R7 a_299_47.n1 a_299_47.n0 80.46
R8 VPWR.n14 VPWR.t2 561.48
R9 VPWR.n17 VPWR.t6 355.821
R10 VPWR.n34 VPWR.n33 311.893
R11 VPWR.n5 VPWR.t8 196.751
R12 VPWR.n10 VPWR.n9 168.909
R13 VPWR.n1 VPWR.n0 166.336
R14 VPWR.n27 VPWR.n26 165.066
R15 VPWR.n2 VPWR.t11 154.717
R16 VPWR.n0 VPWR.t7 58.484
R17 VPWR.n26 VPWR.t1 41.554
R18 VPWR.n26 VPWR.t4 41.554
R19 VPWR.n33 VPWR.t0 41.554
R20 VPWR.n33 VPWR.t5 41.554
R21 VPWR.n0 VPWR.t10 31.605
R22 VPWR.n9 VPWR.t9 26.595
R23 VPWR.n9 VPWR.t3 26.595
R24 VPWR.n4 VPWR.n3 4.65
R25 VPWR.n6 VPWR.n5 4.65
R26 VPWR.n8 VPWR.n7 4.65
R27 VPWR.n11 VPWR.n10 4.65
R28 VPWR.n13 VPWR.n12 4.65
R29 VPWR.n16 VPWR.n15 4.65
R30 VPWR.n19 VPWR.n18 4.65
R31 VPWR.n21 VPWR.n20 4.65
R32 VPWR.n23 VPWR.n22 4.65
R33 VPWR.n25 VPWR.n24 4.65
R34 VPWR.n28 VPWR.n27 4.65
R35 VPWR.n30 VPWR.n29 4.65
R36 VPWR.n32 VPWR.n31 4.65
R37 VPWR.n35 VPWR.n34 3.932
R38 VPWR.n2 VPWR.n1 3.764
R39 VPWR.n15 VPWR.n14 1.05
R40 VPWR.n4 VPWR.n2 0.244
R41 VPWR.n35 VPWR.n32 0.137
R42 VPWR VPWR.n35 0.121
R43 VPWR.n6 VPWR.n4 0.119
R44 VPWR.n8 VPWR.n6 0.119
R45 VPWR.n11 VPWR.n8 0.119
R46 VPWR.n13 VPWR.n11 0.119
R47 VPWR.n16 VPWR.n13 0.119
R48 VPWR.n19 VPWR.n16 0.119
R49 VPWR.n21 VPWR.n19 0.119
R50 VPWR.n23 VPWR.n21 0.119
R51 VPWR.n25 VPWR.n23 0.119
R52 VPWR.n28 VPWR.n25 0.119
R53 VPWR.n30 VPWR.n28 0.119
R54 VPWR.n32 VPWR.n30 0.119
R55 VPWR.n18 VPWR.n17 0.095
R56 VPB.t10 VPB.t9 562.305
R57 VPB.t8 VPB.t3 556.386
R58 VPB.t1 VPB.t5 556.386
R59 VPB.t6 VPB.t0 358.099
R60 VPB.t2 VPB.t6 284.112
R61 VPB.t9 VPB.t12 281.152
R62 VPB.t11 VPB.t10 281.152
R63 VPB.t12 VPB.t13 251.557
R64 VPB.t4 VPB.t11 248.598
R65 VPB.t3 VPB.t4 248.598
R66 VPB.t5 VPB.t2 248.598
R67 VPB.t7 VPB.t1 248.598
R68 VPB.t0 VPB.t8 213.084
R69 VPB VPB.t7 189.408
R70 a_27_47.t0 a_27_47.n3 263.929
R71 a_27_47.n1 a_27_47.t5 263.171
R72 a_27_47.n0 a_27_47.t4 240.108
R73 a_27_47.n0 a_27_47.t2 239.726
R74 a_27_47.n1 a_27_47.t3 227.825
R75 a_27_47.n2 a_27_47.t1 195.572
R76 a_27_47.n2 a_27_47.n1 76
R77 a_27_47.n3 a_27_47.n2 18.495
R78 a_27_47.n3 a_27_47.n0 11.268
R79 a_465_47.n0 a_465_47.t0 88.333
R80 a_465_47.n0 a_465_47.t1 26.393
R81 a_465_47.n1 a_465_47.n0 14.4
R82 a_561_413.n3 a_561_413.n2 422.17
R83 a_561_413.n0 a_561_413.t4 212.079
R84 a_561_413.n2 a_561_413.n1 190.005
R85 a_561_413.n2 a_561_413.n0 172.656
R86 a_561_413.n0 a_561_413.t5 139.779
R87 a_561_413.n3 a_561_413.t2 121.952
R88 a_561_413.t0 a_561_413.n3 91.464
R89 a_561_413.n1 a_561_413.t3 46.666
R90 a_561_413.n1 a_561_413.t1 46.666
R91 VNB VNB.t7 6438.23
R92 VNB.t0 VNB.t5 6082.35
R93 VNB.t9 VNB.t3 5321.88
R94 VNB.t12 VNB.t10 4593.41
R95 VNB.t2 VNB.t1 3494.12
R96 VNB.t6 VNB.t9 3073.53
R97 VNB.t1 VNB.t6 2782.35
R98 VNB.t5 VNB.t2 2717.65
R99 VNB.t7 VNB.t0 2717.65
R100 VNB.t10 VNB.t13 2296.7
R101 VNB.t11 VNB.t12 2296.7
R102 VNB.t13 VNB.t8 2054.95
R103 VNB.t4 VNB.t11 2030.77
R104 VNB.t3 VNB.t4 2030.77
R105 VGND.n5 VGND.t9 190.514
R106 VGND.n17 VGND.t6 148.331
R107 VGND.n2 VGND.t5 111.582
R108 VGND.n1 VGND.n0 108.447
R109 VGND.n33 VGND.n32 107.239
R110 VGND.n26 VGND.n25 106.463
R111 VGND.n10 VGND.n9 92.5
R112 VGND.n0 VGND.t7 54.285
R113 VGND.n25 VGND.t1 38.571
R114 VGND.n25 VGND.t3 38.571
R115 VGND.n32 VGND.t0 38.571
R116 VGND.n32 VGND.t4 38.571
R117 VGND.n0 VGND.t10 25.934
R118 VGND.n9 VGND.t8 24.923
R119 VGND.n9 VGND.t2 24.923
R120 VGND.n4 VGND.n3 4.65
R121 VGND.n6 VGND.n5 4.65
R122 VGND.n8 VGND.n7 4.65
R123 VGND.n12 VGND.n11 4.65
R124 VGND.n14 VGND.n13 4.65
R125 VGND.n16 VGND.n15 4.65
R126 VGND.n18 VGND.n17 4.65
R127 VGND.n20 VGND.n19 4.65
R128 VGND.n22 VGND.n21 4.65
R129 VGND.n24 VGND.n23 4.65
R130 VGND.n27 VGND.n26 4.65
R131 VGND.n29 VGND.n28 4.65
R132 VGND.n31 VGND.n30 4.65
R133 VGND.n34 VGND.n33 3.932
R134 VGND.n2 VGND.n1 3.764
R135 VGND.n11 VGND.n10 0.561
R136 VGND.n4 VGND.n2 0.244
R137 VGND.n34 VGND.n31 0.137
R138 VGND VGND.n34 0.121
R139 VGND.n6 VGND.n4 0.119
R140 VGND.n8 VGND.n6 0.119
R141 VGND.n12 VGND.n8 0.119
R142 VGND.n14 VGND.n12 0.119
R143 VGND.n16 VGND.n14 0.119
R144 VGND.n18 VGND.n16 0.119
R145 VGND.n20 VGND.n18 0.119
R146 VGND.n22 VGND.n20 0.119
R147 VGND.n24 VGND.n22 0.119
R148 VGND.n27 VGND.n24 0.119
R149 VGND.n29 VGND.n27 0.119
R150 VGND.n31 VGND.n29 0.119
R151 a_1313_47.t1 a_1313_47.n2 240.007
R152 a_1313_47.n1 a_1313_47.t2 239.038
R153 a_1313_47.n0 a_1313_47.t4 221.719
R154 a_1313_47.n1 a_1313_47.t3 166.738
R155 a_1313_47.n2 a_1313_47.t0 149.883
R156 a_1313_47.n0 a_1313_47.t5 149.419
R157 a_1313_47.n2 a_1313_47.n1 99.272
R158 a_1313_47.n1 a_1313_47.n0 62.481
R159 Q_N.n4 Q_N.n3 142.958
R160 Q_N.n1 Q_N.n0 92.5
R161 Q_N.n3 Q_N.t0 27.58
R162 Q_N.n2 Q_N.n1 27.32
R163 Q_N.n3 Q_N.t1 26.595
R164 Q_N.n0 Q_N.t2 25.846
R165 Q_N.n0 Q_N.t3 24.923
R166 Q_N Q_N.n2 24.38
R167 Q_N.n2 Q_N 15.881
R168 Q_N.n4 Q_N 9.194
R169 Q_N Q_N.n4 7.483
R170 Q_N.n1 Q_N 6.776
R171 a_193_47.n0 a_193_47.t3 464.325
R172 a_193_47.n0 a_193_47.t2 242.606
R173 a_193_47.n1 a_193_47.t1 230.004
R174 a_193_47.t0 a_193_47.n1 121.759
R175 a_193_47.n1 a_193_47.n0 99.063
R176 a_465_369.t0 a_465_369.t1 134.63
R177 a_724_21.n5 a_724_21.t3 368.328
R178 a_724_21.n0 a_724_21.t7 247.54
R179 a_724_21.n1 a_724_21.t8 212.079
R180 a_724_21.n2 a_724_21.t9 212.079
R181 a_724_21.n4 a_724_21.t0 209.214
R182 a_724_21.n0 a_724_21.t4 154.354
R183 a_724_21.n7 a_724_21.n6 153.497
R184 a_724_21.n5 a_724_21.t5 149.821
R185 a_724_21.n1 a_724_21.t10 139.779
R186 a_724_21.n2 a_724_21.t6 139.779
R187 a_724_21.n1 a_724_21.n0 119.769
R188 a_724_21.n6 a_724_21.n5 107.827
R189 a_724_21.n4 a_724_21.n3 76
R190 a_724_21.n3 a_724_21.n1 60.615
R191 a_724_21.n6 a_724_21.n4 57.563
R192 a_724_21.n7 a_724_21.t2 26.595
R193 a_724_21.t1 a_724_21.n7 26.595
R194 a_724_21.n3 a_724_21.n2 8.763
R195 a_659_47.t0 a_659_47.t1 93.059
R196 GATE_N.n0 GATE_N.t0 269.919
R197 GATE_N.n0 GATE_N.t1 234.573
R198 GATE_N.n1 GATE_N.n0 76
R199 GATE_N GATE_N.n1 10.971
R200 GATE_N.n1 GATE_N 6.791
R201 a_682_413.t0 a_682_413.t1 98.5
R202 Q.n1 Q.n0 146.368
R203 Q.n3 Q.n2 92.5
R204 Q Q.n1 41.61
R205 Q.n0 Q.t0 36.445
R206 Q.n2 Q.t3 34.153
R207 Q.n0 Q.t1 27.58
R208 Q.n2 Q.t2 25.846
R209 Q Q.n3 19.104
R210 Q.n3 Q 7.63
R211 Q.n1 Q 3.988
R212 a_942_47.t0 a_942_47.t1 49.846
R213 RESET_B.n0 RESET_B.t0 241.534
R214 RESET_B.n0 RESET_B.t1 169.234
R215 RESET_B RESET_B.n0 86.278
C0 VPB VPWR 0.18fF
C1 VGND Q_N 0.20fF
C2 VPWR Q_N 0.31fF
C3 VPWR Q 0.20fF
C4 VPWR VGND 0.15fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__dlrbp_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__dlrbp_1 GATE RESET_B Q_N Q D VGND VPWR VNB VPB
X0 a_560_47.t1 a_193_47.t2 a_465_47.t0 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X1 Q.t0 a_711_307.t3 VGND.t2 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 VPWR.t1 D.t0 a_299_47.t0 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X3 a_645_413.t1 a_193_47.t3 a_560_47.t2 VPB.t6 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 VPWR.t5 a_711_307.t4 a_645_413.t0 VPB.t5 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 a_465_47.t1 a_299_47.t2 VGND.t7 VNB.t10 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 VGND.t1 RESET_B.t0 a_941_47.t0 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 Q.t1 a_711_307.t5 VPWR.t3 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 a_560_47.t3 a_27_47.t2 a_465_369.t0 VPB.t10 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9 VPWR.t6 GATE.t0 a_27_47.t0 VPB.t7 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X10 VGND.t3 a_711_307.t6 a_658_47.t0 VNB.t8 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11 Q_N.t0 a_1308_47.t2 VPWR.t8 VPB.t9 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 a_658_47.t1 a_27_47.t3 a_560_47.t0 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X13 VGND.t4 a_711_307.t7 a_1308_47.t1 VNB.t9 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14 a_193_47.t0 a_27_47.t4 VGND.t0 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15 a_711_307.t2 a_560_47.t4 VPWR.t7 VPB.t8 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16 a_941_47.t1 a_560_47.t5 a_711_307.t1 VNB.t7 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X17 VPWR.t4 a_711_307.t8 a_1308_47.t0 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X18 a_193_47.t1 a_27_47.t5 VPWR.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X19 Q_N.t1 a_1308_47.t3 VGND.t8 VNB.t11 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X20 VGND.t6 D.t1 a_299_47.t1 VNB.t6 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21 VPWR.t2 RESET_B.t1 a_711_307.t0 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X22 a_465_369.t1 a_299_47.t3 VPWR.t9 VPB.t11 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X23 VGND.t5 GATE.t1 a_27_47.t1 VNB.t5 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
R0 a_193_47.n0 a_193_47.t2 261.236
R1 a_193_47.n1 a_193_47.t0 230.004
R2 a_193_47.n0 a_193_47.t3 224.251
R3 a_193_47.t1 a_193_47.n1 121.759
R4 a_193_47.n1 a_193_47.n0 12.644
R5 a_465_47.n0 a_465_47.t0 66.666
R6 a_465_47.n0 a_465_47.t1 26.393
R7 a_465_47.n1 a_465_47.n0 14.4
R8 a_560_47.n3 a_560_47.n2 407.446
R9 a_560_47.n0 a_560_47.t4 212.079
R10 a_560_47.n2 a_560_47.n1 193.393
R11 a_560_47.n2 a_560_47.n0 171.618
R12 a_560_47.n0 a_560_47.t5 141.969
R13 a_560_47.n1 a_560_47.t0 68.333
R14 a_560_47.t2 a_560_47.n3 63.321
R15 a_560_47.n3 a_560_47.t3 63.321
R16 a_560_47.n1 a_560_47.t1 45
R17 VNB.t1 VNB.t6 6082.35
R18 VNB.t8 VNB.t7 5321.88
R19 VNB.t2 VNB.t9 4545.05
R20 VNB VNB.t5 4238.23
R21 VNB.t3 VNB.t2 4158.24
R22 VNB.t4 VNB.t0 3170.59
R23 VNB.t0 VNB.t8 3073.53
R24 VNB.t10 VNB.t4 3073.53
R25 VNB.t6 VNB.t10 2717.65
R26 VNB.t5 VNB.t1 2717.65
R27 VNB.t9 VNB.t11 2296.7
R28 VNB.t7 VNB.t3 2151.65
R29 a_711_307.n3 a_711_307.t6 366.001
R30 a_711_307.n0 a_711_307.t8 269.919
R31 a_711_307.n2 a_711_307.t1 231.931
R32 a_711_307.n1 a_711_307.t5 212.079
R33 a_711_307.n0 a_711_307.t7 176.733
R34 a_711_307.n5 a_711_307.n4 153.497
R35 a_711_307.n3 a_711_307.t4 147.494
R36 a_711_307.n1 a_711_307.t3 139.779
R37 a_711_307.n1 a_711_307.n0 137.296
R38 a_711_307.n4 a_711_307.n3 112.46
R39 a_711_307.n2 a_711_307.n1 94.987
R40 a_711_307.n4 a_711_307.n2 69.219
R41 a_711_307.n5 a_711_307.t2 34.475
R42 a_711_307.t0 a_711_307.n5 26.595
R43 VGND.n12 VGND.t3 148.073
R44 VGND.n3 VGND.n0 110.988
R45 VGND.n28 VGND.n27 107.239
R46 VGND.n21 VGND.n20 106.463
R47 VGND.n2 VGND.n1 92.5
R48 VGND.n5 VGND.n4 92.5
R49 VGND.n0 VGND.t4 54.285
R50 VGND.n20 VGND.t7 38.571
R51 VGND.n20 VGND.t6 38.571
R52 VGND.n27 VGND.t0 38.571
R53 VGND.n27 VGND.t5 38.571
R54 VGND.n0 VGND.t8 25.934
R55 VGND.n1 VGND.t2 24.923
R56 VGND.n4 VGND.t1 24.923
R57 VGND.n7 VGND.n6 4.65
R58 VGND.n9 VGND.n8 4.65
R59 VGND.n11 VGND.n10 4.65
R60 VGND.n13 VGND.n12 4.65
R61 VGND.n15 VGND.n14 4.65
R62 VGND.n17 VGND.n16 4.65
R63 VGND.n19 VGND.n18 4.65
R64 VGND.n22 VGND.n21 4.65
R65 VGND.n24 VGND.n23 4.65
R66 VGND.n26 VGND.n25 4.65
R67 VGND.n3 VGND.n2 4.588
R68 VGND.n29 VGND.n28 3.932
R69 VGND.n7 VGND.n3 0.145
R70 VGND.n29 VGND.n26 0.137
R71 VGND VGND.n29 0.121
R72 VGND.n9 VGND.n7 0.119
R73 VGND.n11 VGND.n9 0.119
R74 VGND.n13 VGND.n11 0.119
R75 VGND.n15 VGND.n13 0.119
R76 VGND.n17 VGND.n15 0.119
R77 VGND.n19 VGND.n17 0.119
R78 VGND.n22 VGND.n19 0.119
R79 VGND.n24 VGND.n22 0.119
R80 VGND.n26 VGND.n24 0.119
R81 VGND.n6 VGND.n5 0.112
R82 Q.n0 Q.t1 172.935
R83 Q.n1 Q.t0 117.423
R84 Q Q.n0 9.355
R85 Q Q.n1 9.325
R86 Q.n1 Q 3.108
R87 Q.n0 Q 3.019
R88 D.n0 D.t0 327.642
R89 D.n0 D.t1 157.336
R90 D D.n0 78.594
R91 a_299_47.n0 a_299_47.t3 373.281
R92 a_299_47.t0 a_299_47.n1 292.715
R93 a_299_47.n1 a_299_47.t1 182.645
R94 a_299_47.n0 a_299_47.t2 132.281
R95 a_299_47.n1 a_299_47.n0 80.46
R96 VPWR.n10 VPWR.t7 561.48
R97 VPWR.n13 VPWR.t5 355.821
R98 VPWR.n30 VPWR.n29 311.893
R99 VPWR.n3 VPWR.n2 170.129
R100 VPWR.n23 VPWR.n22 165.066
R101 VPWR.n5 VPWR.n4 146.25
R102 VPWR.n1 VPWR.n0 146.25
R103 VPWR.n2 VPWR.t4 58.484
R104 VPWR.n22 VPWR.t9 41.554
R105 VPWR.n22 VPWR.t1 41.554
R106 VPWR.n29 VPWR.t0 41.554
R107 VPWR.n29 VPWR.t6 41.554
R108 VPWR.n2 VPWR.t8 31.605
R109 VPWR.n0 VPWR.t3 26.595
R110 VPWR.n4 VPWR.t2 26.595
R111 VPWR.n7 VPWR.n6 4.65
R112 VPWR.n9 VPWR.n8 4.65
R113 VPWR.n12 VPWR.n11 4.65
R114 VPWR.n15 VPWR.n14 4.65
R115 VPWR.n17 VPWR.n16 4.65
R116 VPWR.n19 VPWR.n18 4.65
R117 VPWR.n21 VPWR.n20 4.65
R118 VPWR.n24 VPWR.n23 4.65
R119 VPWR.n26 VPWR.n25 4.65
R120 VPWR.n28 VPWR.n27 4.65
R121 VPWR.n3 VPWR.n1 4.376
R122 VPWR.n31 VPWR.n30 3.932
R123 VPWR.n14 VPWR.n13 1.337
R124 VPWR.n11 VPWR.n10 0.668
R125 VPWR.n7 VPWR.n3 0.145
R126 VPWR.n31 VPWR.n28 0.137
R127 VPWR VPWR.n31 0.121
R128 VPWR.n9 VPWR.n7 0.119
R129 VPWR.n12 VPWR.n9 0.119
R130 VPWR.n15 VPWR.n12 0.119
R131 VPWR.n17 VPWR.n15 0.119
R132 VPWR.n19 VPWR.n17 0.119
R133 VPWR.n21 VPWR.n19 0.119
R134 VPWR.n24 VPWR.n21 0.119
R135 VPWR.n26 VPWR.n24 0.119
R136 VPWR.n28 VPWR.n26 0.119
R137 VPWR.n6 VPWR.n5 0.073
R138 VPB.t5 VPB.t8 583.021
R139 VPB.t4 VPB.t3 556.386
R140 VPB.t0 VPB.t1 556.386
R141 VPB.t2 VPB.t4 509.034
R142 VPB.t6 VPB.t5 284.112
R143 VPB.t11 VPB.t10 284.112
R144 VPB.t3 VPB.t9 281.152
R145 VPB.t8 VPB.t2 272.274
R146 VPB.t10 VPB.t6 248.598
R147 VPB.t1 VPB.t11 248.598
R148 VPB.t7 VPB.t0 248.598
R149 VPB VPB.t7 139.096
R150 a_645_413.t0 a_645_413.t1 154.785
R151 RESET_B.n0 RESET_B.t1 241.534
R152 RESET_B.n0 RESET_B.t0 169.234
R153 RESET_B.n1 RESET_B.n0 76
R154 RESET_B.n1 RESET_B 10.86
R155 RESET_B RESET_B.n1 6.981
R156 a_941_47.t0 a_941_47.t1 54.461
R157 a_27_47.n2 a_27_47.t3 448.863
R158 a_27_47.t0 a_27_47.n7 265.057
R159 a_27_47.n5 a_27_47.t5 263.171
R160 a_27_47.n1 a_27_47.t2 241
R161 a_27_47.n5 a_27_47.t4 227.825
R162 a_27_47.n6 a_27_47.t1 196.895
R163 a_27_47.n6 a_27_47.n5 76
R164 a_27_47.n7 a_27_47.n6 18.97
R165 a_27_47.n4 a_27_47.n3 15.872
R166 a_27_47.n3 a_27_47.n2 11.851
R167 a_27_47.n7 a_27_47.n4 9.604
R168 a_27_47.n4 a_27_47.n0 2.327
R169 a_27_47.n3 a_27_47.n1 1.606
R170 a_465_369.t1 a_465_369.t0 134.63
R171 GATE.n0 GATE.t0 272.06
R172 GATE.n0 GATE.t1 236.714
R173 GATE.n1 GATE.n0 76
R174 GATE GATE.n1 11.2
R175 GATE.n1 GATE 6.933
R176 a_658_47.t0 a_658_47.t1 93.059
R177 a_1308_47.t0 a_1308_47.n1 377.062
R178 a_1308_47.n0 a_1308_47.t2 238.589
R179 a_1308_47.n0 a_1308_47.t3 166.289
R180 a_1308_47.n1 a_1308_47.t1 159.243
R181 a_1308_47.n1 a_1308_47.n0 99.466
R182 Q_N.n1 Q_N.t0 172.965
R183 Q_N.n0 Q_N.t1 117.423
R184 Q_N Q_N.n0 97.723
R185 Q_N.n1 Q_N 12.564
R186 Q_N Q_N.n1 4.065
R187 Q_N.n0 Q_N 0.246
C0 VPB VPWR 0.16fF
C1 VPWR Q_N 0.12fF
C2 VPWR Q 0.13fF
C3 VPWR VGND 0.14fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__dlrbp_2.ext - technology: sky130A

.subckt sky130_fd_sc_hd__dlrbp_2 Q RESET_B Q_N D GATE VGND VPWR VNB VPB
X0 VPWR.t11 D.t0 a_299_47.t0 VPB.t13 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1 Q_N.t1 a_1316_47.t2 VGND.t1 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 a_645_413.t0 a_193_47.t2 a_561_413.t3 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3 VPWR.t5 a_711_307.t3 a_645_413.t1 VPB.t7 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 a_561_413.t2 a_193_47.t3 a_465_47.t1 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X5 a_465_47.t0 a_299_47.t2 VGND.t2 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 VGND.t4 a_711_307.t4 a_1316_47.t0 VNB.t7 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7 VPWR.t6 a_711_307.t5 a_1316_47.t1 VPB.t8 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X8 a_561_413.t0 a_27_47.t2 a_465_369.t0 VPB.t5 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9 a_711_307.t1 a_561_413.t4 VPWR.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 VGND.t5 a_711_307.t6 a_659_47.t1 VNB.t8 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11 VPWR.t9 GATE.t0 a_27_47.t0 VPB.t11 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X12 VPWR.t10 RESET_B.t0 a_711_307.t2 VPB.t12 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13 a_659_47.t0 a_27_47.t3 a_561_413.t1 VNB.t5 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X14 VGND.t6 a_711_307.t7 Q.t1 VNB.t9 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X15 VGND.t0 a_1316_47.t3 Q_N.t0 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X16 a_193_47.t0 a_27_47.t4 VGND.t3 VNB.t6 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17 VPWR.t7 a_711_307.t8 Q.t3 VPB.t9 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X18 VPWR.t1 a_1316_47.t4 Q_N.t3 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X19 a_942_47.t0 a_561_413.t5 a_711_307.t0 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X20 Q.t0 a_711_307.t9 VGND.t7 VNB.t10 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X21 Q_N.t2 a_1316_47.t5 VPWR.t2 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X22 a_193_47.t1 a_27_47.t5 VPWR.t4 VPB.t6 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X23 VGND.t9 RESET_B.t1 a_942_47.t1 VNB.t12 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X24 VGND.t10 D.t1 a_299_47.t1 VNB.t13 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X25 Q.t2 a_711_307.t10 VPWR.t8 VPB.t10 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X26 a_465_369.t1 a_299_47.t3 VPWR.t3 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X27 VGND.t8 GATE.t1 a_27_47.t1 VNB.t11 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
R0 D.n0 D.t0 327.642
R1 D.n0 D.t1 157.336
R2 D D.n0 78.594
R3 a_299_47.n0 a_299_47.t3 373.281
R4 a_299_47.t0 a_299_47.n1 292.715
R5 a_299_47.n1 a_299_47.t1 182.645
R6 a_299_47.n0 a_299_47.t2 132.281
R7 a_299_47.n1 a_299_47.n0 80.46
R8 VPWR.n14 VPWR.t0 561.48
R9 VPWR.n17 VPWR.t5 355.821
R10 VPWR.n34 VPWR.n33 311.893
R11 VPWR.n5 VPWR.t7 195.621
R12 VPWR.n1 VPWR.n0 166.336
R13 VPWR.n27 VPWR.n26 165.066
R14 VPWR.n10 VPWR.n9 161.185
R15 VPWR.n2 VPWR.t1 155.734
R16 VPWR.n0 VPWR.t6 56.945
R17 VPWR.n26 VPWR.t3 41.554
R18 VPWR.n26 VPWR.t11 41.554
R19 VPWR.n33 VPWR.t4 41.554
R20 VPWR.n33 VPWR.t9 41.554
R21 VPWR.n9 VPWR.t8 36.445
R22 VPWR.n0 VPWR.t2 33.144
R23 VPWR.n9 VPWR.t10 26.595
R24 VPWR.n4 VPWR.n3 4.65
R25 VPWR.n6 VPWR.n5 4.65
R26 VPWR.n8 VPWR.n7 4.65
R27 VPWR.n11 VPWR.n10 4.65
R28 VPWR.n13 VPWR.n12 4.65
R29 VPWR.n16 VPWR.n15 4.65
R30 VPWR.n19 VPWR.n18 4.65
R31 VPWR.n21 VPWR.n20 4.65
R32 VPWR.n23 VPWR.n22 4.65
R33 VPWR.n25 VPWR.n24 4.65
R34 VPWR.n28 VPWR.n27 4.65
R35 VPWR.n30 VPWR.n29 4.65
R36 VPWR.n32 VPWR.n31 4.65
R37 VPWR.n35 VPWR.n34 3.932
R38 VPWR.n2 VPWR.n1 3.742
R39 VPWR.n18 VPWR.n17 1.337
R40 VPWR.n15 VPWR.n14 1.05
R41 VPWR.n4 VPWR.n2 0.245
R42 VPWR.n35 VPWR.n32 0.137
R43 VPWR VPWR.n35 0.121
R44 VPWR.n6 VPWR.n4 0.119
R45 VPWR.n8 VPWR.n6 0.119
R46 VPWR.n11 VPWR.n8 0.119
R47 VPWR.n13 VPWR.n11 0.119
R48 VPWR.n16 VPWR.n13 0.119
R49 VPWR.n19 VPWR.n16 0.119
R50 VPWR.n21 VPWR.n19 0.119
R51 VPWR.n23 VPWR.n21 0.119
R52 VPWR.n25 VPWR.n23 0.119
R53 VPWR.n28 VPWR.n25 0.119
R54 VPWR.n30 VPWR.n28 0.119
R55 VPWR.n32 VPWR.n30 0.119
R56 VPB.t7 VPB.t0 594.859
R57 VPB.t9 VPB.t8 556.386
R58 VPB.t6 VPB.t13 556.386
R59 VPB.t4 VPB.t7 284.112
R60 VPB.t3 VPB.t5 284.112
R61 VPB.t8 VPB.t2 281.152
R62 VPB.t12 VPB.t10 278.193
R63 VPB.t10 VPB.t9 260.436
R64 VPB.t0 VPB.t12 254.517
R65 VPB.t2 VPB.t1 248.598
R66 VPB.t5 VPB.t4 248.598
R67 VPB.t13 VPB.t3 248.598
R68 VPB.t11 VPB.t6 248.598
R69 VPB VPB.t11 139.096
R70 a_1316_47.n1 a_1316_47.t5 300.445
R71 a_1316_47.t1 a_1316_47.n3 245.874
R72 a_1316_47.n1 a_1316_47.t2 228.145
R73 a_1316_47.n0 a_1316_47.t4 221.719
R74 a_1316_47.n3 a_1316_47.t0 156.187
R75 a_1316_47.n0 a_1316_47.t3 149.419
R76 a_1316_47.n3 a_1316_47.n2 94.23
R77 a_1316_47.n2 a_1316_47.n0 83.903
R78 a_1316_47.n2 a_1316_47.n1 0.892
R79 VGND.n5 VGND.t6 189.881
R80 VGND.n17 VGND.t5 148.331
R81 VGND.n2 VGND.t0 112.437
R82 VGND.n1 VGND.n0 108.447
R83 VGND.n33 VGND.n32 107.239
R84 VGND.n26 VGND.n25 106.463
R85 VGND.n10 VGND.n9 92.5
R86 VGND.n0 VGND.t4 52.857
R87 VGND.n25 VGND.t2 38.571
R88 VGND.n25 VGND.t10 38.571
R89 VGND.n32 VGND.t3 38.571
R90 VGND.n32 VGND.t8 38.571
R91 VGND.n9 VGND.t7 34.153
R92 VGND.n0 VGND.t1 27.362
R93 VGND.n9 VGND.t9 24.923
R94 VGND.n4 VGND.n3 4.65
R95 VGND.n6 VGND.n5 4.65
R96 VGND.n8 VGND.n7 4.65
R97 VGND.n12 VGND.n11 4.65
R98 VGND.n14 VGND.n13 4.65
R99 VGND.n16 VGND.n15 4.65
R100 VGND.n18 VGND.n17 4.65
R101 VGND.n20 VGND.n19 4.65
R102 VGND.n22 VGND.n21 4.65
R103 VGND.n24 VGND.n23 4.65
R104 VGND.n27 VGND.n26 4.65
R105 VGND.n29 VGND.n28 4.65
R106 VGND.n31 VGND.n30 4.65
R107 VGND.n34 VGND.n33 3.932
R108 VGND.n2 VGND.n1 3.742
R109 VGND.n11 VGND.n10 0.336
R110 VGND.n4 VGND.n2 0.245
R111 VGND.n34 VGND.n31 0.137
R112 VGND VGND.n34 0.121
R113 VGND.n6 VGND.n4 0.119
R114 VGND.n8 VGND.n6 0.119
R115 VGND.n12 VGND.n8 0.119
R116 VGND.n14 VGND.n12 0.119
R117 VGND.n16 VGND.n14 0.119
R118 VGND.n18 VGND.n16 0.119
R119 VGND.n20 VGND.n18 0.119
R120 VGND.n22 VGND.n20 0.119
R121 VGND.n24 VGND.n22 0.119
R122 VGND.n27 VGND.n24 0.119
R123 VGND.n29 VGND.n27 0.119
R124 VGND.n31 VGND.n29 0.119
R125 Q_N.n4 Q_N.n3 142.894
R126 Q_N.n1 Q_N.n0 92.5
R127 Q_N.n2 Q_N.n1 30.885
R128 Q_N Q_N.n2 30.298
R129 Q_N.n3 Q_N.t3 26.595
R130 Q_N.n3 Q_N.t2 26.595
R131 Q_N.n0 Q_N.t0 24.923
R132 Q_N.n0 Q_N.t1 24.923
R133 Q_N.n2 Q_N 14.933
R134 Q_N.n4 Q_N 9.375
R135 Q_N Q_N.n4 7.629
R136 Q_N.n1 Q_N 6.912
R137 VNB.t6 VNB.t13 6082.35
R138 VNB.t8 VNB.t0 5321.88
R139 VNB.t9 VNB.t7 4545.05
R140 VNB VNB.t11 4238.23
R141 VNB.t3 VNB.t4 3494.12
R142 VNB.t5 VNB.t8 3073.53
R143 VNB.t4 VNB.t5 2782.35
R144 VNB.t13 VNB.t3 2717.65
R145 VNB.t11 VNB.t6 2717.65
R146 VNB.t7 VNB.t2 2296.7
R147 VNB.t12 VNB.t10 2272.53
R148 VNB.t10 VNB.t9 2127.47
R149 VNB.t0 VNB.t12 2079.12
R150 VNB.t2 VNB.t1 2030.77
R151 a_193_47.n0 a_193_47.t3 255.766
R152 a_193_47.n1 a_193_47.t0 230.004
R153 a_193_47.n0 a_193_47.t2 146.481
R154 a_193_47.t1 a_193_47.n1 121.759
R155 a_193_47.n1 a_193_47.n0 6.199
R156 a_561_413.n3 a_561_413.n2 407.446
R157 a_561_413.n0 a_561_413.t4 212.079
R158 a_561_413.n2 a_561_413.n1 188.122
R159 a_561_413.n2 a_561_413.n0 174.539
R160 a_561_413.n0 a_561_413.t5 139.779
R161 a_561_413.n3 a_561_413.t3 63.321
R162 a_561_413.t0 a_561_413.n3 63.321
R163 a_561_413.n1 a_561_413.t1 46.666
R164 a_561_413.n1 a_561_413.t2 46.666
R165 a_645_413.t0 a_645_413.t1 154.785
R166 a_711_307.n4 a_711_307.t6 366.001
R167 a_711_307.n0 a_711_307.t5 269.919
R168 a_711_307.n2 a_711_307.t10 212.079
R169 a_711_307.n1 a_711_307.t8 212.079
R170 a_711_307.n3 a_711_307.t0 204.937
R171 a_711_307.n0 a_711_307.t4 176.733
R172 a_711_307.n6 a_711_307.n5 153.497
R173 a_711_307.n4 a_711_307.t3 147.494
R174 a_711_307.n2 a_711_307.t9 139.779
R175 a_711_307.n1 a_711_307.t7 139.779
R176 a_711_307.n1 a_711_307.n0 137.296
R177 a_711_307.n5 a_711_307.n4 112.072
R178 a_711_307.n3 a_711_307.n2 76
R179 a_711_307.n2 a_711_307.n1 64.266
R180 a_711_307.n5 a_711_307.n3 58.82
R181 a_711_307.t1 a_711_307.n6 28.565
R182 a_711_307.n6 a_711_307.t2 26.595
R183 a_465_47.n0 a_465_47.t1 88.333
R184 a_465_47.n0 a_465_47.t0 26.393
R185 a_465_47.n1 a_465_47.n0 14.4
R186 a_27_47.n2 a_27_47.t3 450.47
R187 a_27_47.t0 a_27_47.n7 265.057
R188 a_27_47.n5 a_27_47.t5 263.171
R189 a_27_47.n1 a_27_47.t2 241
R190 a_27_47.n5 a_27_47.t4 227.825
R191 a_27_47.n6 a_27_47.t1 196.895
R192 a_27_47.n6 a_27_47.n5 76
R193 a_27_47.n7 a_27_47.n6 18.97
R194 a_27_47.n4 a_27_47.n3 15.872
R195 a_27_47.n3 a_27_47.n2 11.851
R196 a_27_47.n7 a_27_47.n4 9.604
R197 a_27_47.n4 a_27_47.n0 2.327
R198 a_27_47.n3 a_27_47.n1 1.606
R199 a_465_369.t1 a_465_369.t0 134.63
R200 a_659_47.t1 a_659_47.t0 93.059
R201 GATE.n0 GATE.t0 269.919
R202 GATE.n0 GATE.t1 234.573
R203 GATE.n1 GATE.n0 76
R204 GATE GATE.n1 10.971
R205 GATE.n1 GATE 6.791
R206 RESET_B.n0 RESET_B.t0 241.534
R207 RESET_B.n0 RESET_B.t1 169.234
R208 RESET_B RESET_B.n0 85.89
R209 Q.n1 Q.n0 146.375
R210 Q.n3 Q.n2 92.5
R211 Q Q.n1 37.799
R212 Q.n0 Q.t2 30.535
R213 Q.n2 Q.t0 28.615
R214 Q Q.n3 28.552
R215 Q.n0 Q.t3 26.595
R216 Q.n2 Q.t1 24.923
R217 Q.n3 Q 11.67
R218 Q.n1 Q 4.228
R219 a_942_47.t0 a_942_47.t1 51.692
C0 VGND Q_N 0.20fF
C1 VPWR Q_N 0.30fF
C2 VGND Q 0.12fF
C3 VPWR Q 0.22fF
C4 VPWR VGND 0.15fF
C5 VPB VPWR 0.18fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__dlrtn_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__dlrtn_1 RESET_B Q D GATE_N VGND VPWR VNB VPB
X0 VPWR.t6 D.t0 a_299_47.t1 VPB.t7 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1 a_561_413.t0 a_27_47.t2 a_465_47.t0 VNB.t6 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X2 a_465_47.t1 a_299_47.t2 VGND.t5 VNB.t7 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3 a_561_413.t2 a_193_47.t2 a_465_369.t0 VPB.t9 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 a_724_21.t1 a_561_413.t4 VPWR.t7 VPB.t8 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 VGND.t0 a_724_21.t3 a_659_47.t1 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 VPWR.t3 GATE_N.t0 a_27_47.t0 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X7 a_659_47.t0 a_193_47.t3 a_561_413.t3 VNB.t9 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X8 VPWR.t0 a_724_21.t4 a_682_413.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9 Q.t0 a_724_21.t5 VPWR.t1 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 a_193_47.t1 a_27_47.t3 VGND.t4 VNB.t5 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11 a_682_413.t1 a_27_47.t4 a_561_413.t1 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12 a_942_47.t0 a_561_413.t5 a_724_21.t0 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 a_193_47.t0 a_27_47.t5 VPWR.t4 VPB.t5 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X14 Q.t1 a_724_21.t6 VGND.t1 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X15 VPWR.t2 RESET_B.t0 a_724_21.t2 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16 VGND.t6 D.t1 a_299_47.t0 VNB.t8 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17 VGND.t2 RESET_B.t1 a_942_47.t1 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X18 a_465_369.t1 a_299_47.t3 VPWR.t5 VPB.t6 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X19 VGND.t3 GATE_N.t1 a_27_47.t1 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
R0 D.n0 D.t0 327.642
R1 D.n0 D.t1 157.336
R2 D D.n0 78.594
R3 a_299_47.n0 a_299_47.t3 373.281
R4 a_299_47.t1 a_299_47.n1 292.715
R5 a_299_47.n1 a_299_47.t0 182.645
R6 a_299_47.n0 a_299_47.t2 132.281
R7 a_299_47.n1 a_299_47.n0 80.46
R8 VPWR.n9 VPWR.t7 578.851
R9 VPWR.n11 VPWR.t0 374.358
R10 VPWR.n27 VPWR.n0 311.893
R11 VPWR.n2 VPWR.n1 292.665
R12 VPWR.n4 VPWR.n3 292.5
R13 VPWR.n20 VPWR.n19 165.066
R14 VPWR.n3 VPWR.t2 43.34
R15 VPWR.n19 VPWR.t5 41.554
R16 VPWR.n19 VPWR.t6 41.554
R17 VPWR.n0 VPWR.t4 41.554
R18 VPWR.n0 VPWR.t3 41.554
R19 VPWR.n1 VPWR.t1 26.595
R20 VPWR.n28 VPWR.n27 26.108
R21 VPWR.n27 VPWR.n26 4.65
R22 VPWR.n6 VPWR.n5 4.65
R23 VPWR.n8 VPWR.n7 4.65
R24 VPWR.n10 VPWR.n9 4.65
R25 VPWR.n12 VPWR.n11 4.65
R26 VPWR.n14 VPWR.n13 4.65
R27 VPWR.n16 VPWR.n15 4.65
R28 VPWR.n18 VPWR.n17 4.65
R29 VPWR.n21 VPWR.n20 4.65
R30 VPWR.n23 VPWR.n22 4.65
R31 VPWR.n25 VPWR.n24 4.65
R32 VPWR.n6 VPWR.n2 4.112
R33 VPWR.n5 VPWR.n4 1.146
R34 VPWR.n8 VPWR.n6 0.119
R35 VPWR.n10 VPWR.n8 0.119
R36 VPWR.n12 VPWR.n10 0.119
R37 VPWR.n14 VPWR.n12 0.119
R38 VPWR.n16 VPWR.n14 0.119
R39 VPWR.n18 VPWR.n16 0.119
R40 VPWR.n21 VPWR.n18 0.119
R41 VPWR.n23 VPWR.n21 0.119
R42 VPWR.n25 VPWR.n23 0.119
R43 VPWR.n26 VPWR.n25 0.119
R44 VPWR.n26 VPWR 0.118
R45 VPWR VPWR.n28 0.02
R46 VPWR.n28 VPWR 0.001
R47 VPB.t0 VPB.t8 556.386
R48 VPB.t5 VPB.t7 556.386
R49 VPB.t2 VPB.t1 541.588
R50 VPB.t9 VPB.t4 358.099
R51 VPB.t6 VPB.t9 284.112
R52 VPB.t8 VPB.t2 248.598
R53 VPB.t7 VPB.t6 248.598
R54 VPB.t3 VPB.t5 248.598
R55 VPB.t4 VPB.t0 213.084
R56 VPB VPB.t3 139.096
R57 a_27_47.t0 a_27_47.n3 269.575
R58 a_27_47.n1 a_27_47.t5 263.171
R59 a_27_47.n0 a_27_47.t4 240.108
R60 a_27_47.n0 a_27_47.t2 239.726
R61 a_27_47.n1 a_27_47.t3 227.825
R62 a_27_47.n2 a_27_47.t1 202.368
R63 a_27_47.n2 a_27_47.n1 76
R64 a_27_47.n3 a_27_47.n2 18.97
R65 a_27_47.n3 a_27_47.n0 11.268
R66 a_465_47.n0 a_465_47.t0 88.333
R67 a_465_47.n0 a_465_47.t1 26.393
R68 a_465_47.n1 a_465_47.n0 14.4
R69 a_561_413.n3 a_561_413.n2 454.57
R70 a_561_413.n0 a_561_413.t4 221.719
R71 a_561_413.n2 a_561_413.n1 188.773
R72 a_561_413.n2 a_561_413.n0 177.437
R73 a_561_413.n0 a_561_413.t5 149.419
R74 a_561_413.n3 a_561_413.t2 121.952
R75 a_561_413.t1 a_561_413.n3 91.464
R76 a_561_413.n1 a_561_413.t3 46.666
R77 a_561_413.n1 a_561_413.t0 46.666
R78 VNB.t5 VNB.t8 6082.35
R79 VNB.t0 VNB.t2 5321.88
R80 VNB.t3 VNB.t1 4424.17
R81 VNB VNB.t4 4238.23
R82 VNB.t7 VNB.t6 3494.12
R83 VNB.t9 VNB.t0 3073.53
R84 VNB.t6 VNB.t9 2782.35
R85 VNB.t8 VNB.t7 2717.65
R86 VNB.t4 VNB.t5 2717.65
R87 VNB.t2 VNB.t3 2030.77
R88 VGND.n4 VGND.t0 148.331
R89 VGND.n26 VGND.n25 107.239
R90 VGND.n2 VGND.n1 106.463
R91 VGND.n9 VGND.n8 92.598
R92 VGND.n7 VGND.n6 92.5
R93 VGND.n8 VGND.n7 74.769
R94 VGND.n7 VGND.t2 40.615
R95 VGND.n1 VGND.t5 38.571
R96 VGND.n1 VGND.t6 38.571
R97 VGND.n25 VGND.t4 38.571
R98 VGND.n25 VGND.t3 38.571
R99 VGND.n13 VGND.n12 34.635
R100 VGND.n18 VGND.n17 34.635
R101 VGND.n19 VGND.n18 34.635
R102 VGND.n24 VGND.n23 34.635
R103 VGND.n8 VGND.t1 25.846
R104 VGND.n19 VGND.n2 24.47
R105 VGND.n12 VGND.n11 24.33
R106 VGND.n26 VGND.n24 22.964
R107 VGND.n13 VGND.n4 22.588
R108 VGND.n17 VGND.n4 21.835
R109 VGND.n23 VGND.n2 19.952
R110 VGND.n9 VGND.n6 8.998
R111 VGND.n11 VGND.n10 4.65
R112 VGND.n12 VGND.n5 4.65
R113 VGND.n14 VGND.n13 4.65
R114 VGND.n15 VGND.n4 4.65
R115 VGND.n17 VGND.n16 4.65
R116 VGND.n18 VGND.n3 4.65
R117 VGND.n20 VGND.n19 4.65
R118 VGND.n21 VGND.n2 4.65
R119 VGND.n23 VGND.n22 4.65
R120 VGND.n24 VGND.n0 4.65
R121 VGND.n10 VGND.n9 4.133
R122 VGND.n27 VGND.n26 3.932
R123 VGND.n11 VGND.n6 1.347
R124 VGND.n27 VGND.n0 0.137
R125 VGND.n10 VGND.n5 0.119
R126 VGND.n14 VGND.n5 0.119
R127 VGND.n15 VGND.n14 0.119
R128 VGND.n16 VGND.n15 0.119
R129 VGND.n16 VGND.n3 0.119
R130 VGND.n20 VGND.n3 0.119
R131 VGND.n21 VGND.n20 0.119
R132 VGND.n22 VGND.n21 0.119
R133 VGND.n22 VGND.n0 0.119
R134 VGND VGND.n27 0.101
R135 a_193_47.n0 a_193_47.t3 464.325
R136 a_193_47.n0 a_193_47.t2 242.606
R137 a_193_47.n1 a_193_47.t1 230.004
R138 a_193_47.t0 a_193_47.n1 121.759
R139 a_193_47.n1 a_193_47.n0 99.063
R140 a_465_369.t1 a_465_369.t0 134.63
R141 a_724_21.n2 a_724_21.t3 368.328
R142 a_724_21.n0 a_724_21.t5 235.47
R143 a_724_21.n1 a_724_21.t0 181.805
R144 a_724_21.n0 a_724_21.t6 163.17
R145 a_724_21.n4 a_724_21.n3 152.768
R146 a_724_21.n2 a_724_21.t4 149.821
R147 a_724_21.n3 a_724_21.n2 111.684
R148 a_724_21.n1 a_724_21.n0 76
R149 a_724_21.n3 a_724_21.n1 50.684
R150 a_724_21.n4 a_724_21.t2 26.595
R151 a_724_21.t1 a_724_21.n4 26.595
R152 a_659_47.t1 a_659_47.t0 93.059
R153 GATE_N.n0 GATE_N.t0 269.919
R154 GATE_N.n0 GATE_N.t1 234.573
R155 GATE_N.n1 GATE_N.n0 76
R156 GATE_N GATE_N.n1 10.971
R157 GATE_N.n1 GATE_N 6.791
R158 a_682_413.t0 a_682_413.t1 98.5
R159 Q.n0 Q.t0 226.813
R160 Q.n1 Q.t1 117.423
R161 Q Q.n1 9.107
R162 Q Q.n0 8.551
R163 Q.n0 Q 7.973
R164 Q.n1 Q 7.63
R165 a_942_47.t0 a_942_47.t1 49.846
R166 RESET_B.n0 RESET_B.t0 241.534
R167 RESET_B.n0 RESET_B.t1 169.234
R168 RESET_B.n1 RESET_B.n0 76
R169 RESET_B.n1 RESET_B 10.666
R170 RESET_B RESET_B.n1 7.175
C0 VPWR VGND 0.11fF
C1 VPB VPWR 0.13fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__dlrtn_2.ext - technology: sky130A

.subckt sky130_fd_sc_hd__dlrtn_2 RESET_B Q D GATE_N VGND VPWR VNB VPB
X0 a_560_47.t0 a_27_47.t2 a_465_47.t1 VNB.t7 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X1 VPWR.t0 D.t0 a_299_47.t1 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X2 a_645_413.t1 a_27_47.t3 a_560_47.t1 VPB.t6 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3 VPWR.t2 a_711_307.t3 a_645_413.t0 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 a_465_47.t0 a_299_47.t2 VGND.t6 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 VPWR.t8 RESET_B.t0 a_711_307.t2 VPB.t10 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 a_560_47.t2 a_193_47.t2 a_465_369.t0 VPB.t9 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7 VPWR.t1 GATE_N.t0 a_27_47.t0 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X8 Q.t3 a_711_307.t4 VPWR.t3 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 VGND.t4 a_711_307.t5 a_658_47.t1 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10 a_658_47.t0 a_193_47.t3 a_560_47.t3 VNB.t9 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X11 VPWR.t4 a_711_307.t6 Q.t2 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 a_193_47.t0 a_27_47.t4 VGND.t5 VNB.t6 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13 a_711_307.t0 a_560_47.t4 VPWR.t7 VPB.t8 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14 Q.t1 a_711_307.t7 VGND.t2 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X15 a_941_47.t1 a_560_47.t5 a_711_307.t1 VNB.t8 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X16 a_193_47.t1 a_27_47.t5 VPWR.t5 VPB.t5 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X17 VGND.t3 a_711_307.t8 Q.t0 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X18 VGND.t0 D.t1 a_299_47.t0 VNB.t5 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19 VGND.t7 RESET_B.t1 a_941_47.t0 VNB.t10 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X20 a_465_369.t1 a_299_47.t3 VPWR.t6 VPB.t7 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X21 VGND.t1 GATE_N.t1 a_27_47.t1 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
R0 a_27_47.t0 a_27_47.n3 269.575
R1 a_27_47.n1 a_27_47.t5 263.171
R2 a_27_47.n0 a_27_47.t2 239.674
R3 a_27_47.n0 a_27_47.t3 232.156
R4 a_27_47.n1 a_27_47.t4 227.825
R5 a_27_47.n2 a_27_47.t1 202.368
R6 a_27_47.n2 a_27_47.n1 76
R7 a_27_47.n3 a_27_47.n2 18.97
R8 a_27_47.n3 a_27_47.n0 11.268
R9 a_465_47.n0 a_465_47.t1 66.666
R10 a_465_47.n0 a_465_47.t0 26.393
R11 a_465_47.n1 a_465_47.n0 14.4
R12 a_560_47.n3 a_560_47.n2 462.193
R13 a_560_47.n0 a_560_47.t4 268.312
R14 a_560_47.n2 a_560_47.n1 188.618
R15 a_560_47.n2 a_560_47.n0 176.796
R16 a_560_47.n0 a_560_47.t5 151.204
R17 a_560_47.t1 a_560_47.n3 63.321
R18 a_560_47.n3 a_560_47.t2 63.321
R19 a_560_47.n1 a_560_47.t0 60
R20 a_560_47.n1 a_560_47.t3 53.333
R21 VNB.t6 VNB.t5 6082.35
R22 VNB.t2 VNB.t8 5321.88
R23 VNB VNB.t1 4238.23
R24 VNB.t7 VNB.t9 3170.59
R25 VNB.t9 VNB.t2 3073.53
R26 VNB.t0 VNB.t7 3073.53
R27 VNB.t5 VNB.t0 2717.65
R28 VNB.t1 VNB.t6 2717.65
R29 VNB.t10 VNB.t3 2417.58
R30 VNB.t3 VNB.t4 2030.77
R31 VNB.t8 VNB.t10 2030.77
R32 D.n0 D.t0 327.642
R33 D.n0 D.t1 157.336
R34 D D.n0 78.594
R35 a_299_47.n0 a_299_47.t3 373.281
R36 a_299_47.t1 a_299_47.n1 289.243
R37 a_299_47.n1 a_299_47.t0 180.931
R38 a_299_47.n0 a_299_47.t2 132.281
R39 a_299_47.n1 a_299_47.n0 80.266
R40 VPWR.n10 VPWR.t7 578.851
R41 VPWR.n4 VPWR.t2 392.618
R42 VPWR.n23 VPWR.n22 311.893
R43 VPWR.n6 VPWR.t4 260.952
R44 VPWR.n2 VPWR.n1 165.066
R45 VPWR.n8 VPWR.n7 161.588
R46 VPWR.n1 VPWR.t6 41.554
R47 VPWR.n1 VPWR.t0 41.554
R48 VPWR.n22 VPWR.t5 41.554
R49 VPWR.n22 VPWR.t1 41.554
R50 VPWR.n15 VPWR.n14 34.635
R51 VPWR.n16 VPWR.n15 34.635
R52 VPWR.n21 VPWR.n20 34.635
R53 VPWR.n7 VPWR.t3 32.505
R54 VPWR.n7 VPWR.t8 32.505
R55 VPWR.n14 VPWR.n4 26.352
R56 VPWR.n20 VPWR.n2 25.976
R57 VPWR.n23 VPWR.n21 22.964
R58 VPWR.n10 VPWR.n9 20.329
R59 VPWR.n9 VPWR.n8 19.576
R60 VPWR.n16 VPWR.n2 19.576
R61 VPWR.n10 VPWR.n4 12.8
R62 VPWR.n9 VPWR.n5 4.65
R63 VPWR.n11 VPWR.n10 4.65
R64 VPWR.n12 VPWR.n4 4.65
R65 VPWR.n14 VPWR.n13 4.65
R66 VPWR.n15 VPWR.n3 4.65
R67 VPWR.n17 VPWR.n16 4.65
R68 VPWR.n18 VPWR.n2 4.65
R69 VPWR.n20 VPWR.n19 4.65
R70 VPWR.n21 VPWR.n0 4.65
R71 VPWR.n24 VPWR.n23 3.932
R72 VPWR.n8 VPWR.n6 3.832
R73 VPWR.n6 VPWR.n5 0.233
R74 VPWR.n24 VPWR.n0 0.137
R75 VPWR.n11 VPWR.n5 0.119
R76 VPWR.n12 VPWR.n11 0.119
R77 VPWR.n13 VPWR.n12 0.119
R78 VPWR.n13 VPWR.n3 0.119
R79 VPWR.n17 VPWR.n3 0.119
R80 VPWR.n18 VPWR.n17 0.119
R81 VPWR.n19 VPWR.n18 0.119
R82 VPWR.n19 VPWR.n0 0.119
R83 VPWR VPWR.n24 0.101
R84 VPB.t2 VPB.t8 583.021
R85 VPB.t5 VPB.t0 556.386
R86 VPB.t10 VPB.t3 284.112
R87 VPB.t6 VPB.t2 284.112
R88 VPB.t7 VPB.t9 284.112
R89 VPB.t3 VPB.t4 269.314
R90 VPB.t8 VPB.t10 248.598
R91 VPB.t9 VPB.t6 248.598
R92 VPB.t0 VPB.t7 248.598
R93 VPB.t1 VPB.t5 248.598
R94 VPB VPB.t1 139.096
R95 a_645_413.t0 a_645_413.t1 154.785
R96 a_711_307.n4 a_711_307.t5 366.001
R97 a_711_307.n2 a_711_307.t4 214.269
R98 a_711_307.n0 a_711_307.t6 212.079
R99 a_711_307.n3 a_711_307.t1 177.868
R100 a_711_307.n6 a_711_307.n5 152.768
R101 a_711_307.n4 a_711_307.t3 147.494
R102 a_711_307.n0 a_711_307.t8 139.779
R103 a_711_307.n1 a_711_307.t7 139.779
R104 a_711_307.n5 a_711_307.n4 110.909
R105 a_711_307.n3 a_711_307.n2 76
R106 a_711_307.n5 a_711_307.n3 71.134
R107 a_711_307.n1 a_711_307.n0 61.345
R108 a_711_307.n6 a_711_307.t2 26.595
R109 a_711_307.t0 a_711_307.n6 26.595
R110 a_711_307.n2 a_711_307.n1 2.921
R111 VGND.n6 VGND.t3 198.41
R112 VGND.n4 VGND.t4 148.073
R113 VGND.n23 VGND.n22 107.239
R114 VGND.n8 VGND.n7 106.463
R115 VGND.n2 VGND.n1 106.463
R116 VGND.n7 VGND.t2 39.692
R117 VGND.n1 VGND.t6 38.571
R118 VGND.n1 VGND.t0 38.571
R119 VGND.n22 VGND.t5 38.571
R120 VGND.n22 VGND.t1 38.571
R121 VGND.n10 VGND.n9 34.635
R122 VGND.n15 VGND.n14 34.635
R123 VGND.n16 VGND.n15 34.635
R124 VGND.n21 VGND.n20 34.635
R125 VGND.n7 VGND.t7 24.923
R126 VGND.n16 VGND.n2 24.47
R127 VGND.n23 VGND.n21 22.964
R128 VGND.n10 VGND.n4 22.588
R129 VGND.n14 VGND.n4 21.458
R130 VGND.n9 VGND.n8 19.952
R131 VGND.n20 VGND.n2 19.952
R132 VGND.n9 VGND.n5 4.65
R133 VGND.n11 VGND.n10 4.65
R134 VGND.n12 VGND.n4 4.65
R135 VGND.n14 VGND.n13 4.65
R136 VGND.n15 VGND.n3 4.65
R137 VGND.n17 VGND.n16 4.65
R138 VGND.n18 VGND.n2 4.65
R139 VGND.n20 VGND.n19 4.65
R140 VGND.n21 VGND.n0 4.65
R141 VGND.n24 VGND.n23 3.932
R142 VGND.n8 VGND.n6 3.897
R143 VGND.n6 VGND.n5 0.224
R144 VGND.n24 VGND.n0 0.137
R145 VGND.n11 VGND.n5 0.119
R146 VGND.n12 VGND.n11 0.119
R147 VGND.n13 VGND.n12 0.119
R148 VGND.n13 VGND.n3 0.119
R149 VGND.n17 VGND.n3 0.119
R150 VGND.n18 VGND.n17 0.119
R151 VGND.n19 VGND.n18 0.119
R152 VGND.n19 VGND.n0 0.119
R153 VGND VGND.n24 0.101
R154 RESET_B.n0 RESET_B.t0 241.534
R155 RESET_B.n0 RESET_B.t1 169.234
R156 RESET_B RESET_B.n0 86.86
R157 a_193_47.n0 a_193_47.t3 462.718
R158 a_193_47.n0 a_193_47.t2 242.606
R159 a_193_47.n1 a_193_47.t0 230.004
R160 a_193_47.t1 a_193_47.n1 121.759
R161 a_193_47.n1 a_193_47.n0 99.063
R162 a_465_369.t1 a_465_369.t0 134.63
R163 GATE_N.n0 GATE_N.t0 269.919
R164 GATE_N.n0 GATE_N.t1 234.573
R165 GATE_N.n1 GATE_N.n0 76
R166 GATE_N GATE_N.n1 10.971
R167 GATE_N.n1 GATE_N 6.791
R168 Q Q.n2 300.796
R169 Q.n1 Q.n0 146.59
R170 Q.n2 Q.t2 30.535
R171 Q.n2 Q.t3 29.55
R172 Q.n0 Q.t0 24.923
R173 Q.n0 Q.t1 24.923
R174 Q.n1 Q 9.6
R175 Q.n3 Q 4.828
R176 Q Q.n3 2.807
R177 Q.n1 Q 2.188
R178 Q.n3 Q.n1 0.547
R179 a_658_47.t1 a_658_47.t0 93.059
R180 a_941_47.t0 a_941_47.t1 49.846
C0 VGND Q 0.19fF
C1 VPB VPWR 0.14fF
C2 Q VPWR 0.26fF
C3 VGND VPWR 0.10fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__dlrtn_4.ext - technology: sky130A

.subckt sky130_fd_sc_hd__dlrtn_4 Q D GATE_N RESET_B VPWR VGND VNB VPB
X0 VPWR.t7 RESET_B.t0 a_725_21.t2 VPB.t8 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_466_47.t0 a_300_47.t2 VGND.t1 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 a_562_413.t1 a_27_47.t2 a_466_47.t1 VNB.t10 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X3 Q.t7 a_725_21.t3 VPWR.t5 VPB.t7 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 VGND.t6 a_725_21.t4 a_660_47.t1 VNB.t8 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 VGND.t5 a_725_21.t5 Q.t3 VNB.t7 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 a_466_369.t1 a_300_47.t3 VPWR.t8 VPB.t9 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X7 VPWR.t10 GATE_N.t0 a_27_47.t0 VPB.t12 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X8 VPWR.t0 D.t0 a_300_47.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X9 VPWR.t4 a_725_21.t6 Q.t6 VPB.t6 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 VGND.t4 a_725_21.t7 Q.t2 VNB.t6 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 a_562_413.t2 a_193_47.t2 a_466_369.t0 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12 a_725_21.t0 a_562_413.t4 VPWR.t1 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13 a_193_47.t0 a_27_47.t3 VGND.t8 VNB.t11 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14 VPWR.t6 a_725_21.t8 a_683_413.t1 VPB.t5 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15 a_943_47.t0 a_562_413.t5 a_725_21.t1 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X16 Q.t1 a_725_21.t9 VGND.t3 VNB.t5 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X17 Q.t5 a_725_21.t10 VPWR.t3 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X18 a_683_413.t0 a_27_47.t4 a_562_413.t0 VPB.t10 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19 a_193_47.t1 a_27_47.t5 VPWR.t9 VPB.t11 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X20 a_660_47.t0 a_193_47.t3 a_562_413.t3 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X21 Q.t0 a_725_21.t11 VGND.t2 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X22 VGND.t0 D.t1 a_300_47.t1 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23 VGND.t7 RESET_B.t1 a_943_47.t1 VNB.t9 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X24 VPWR.t2 a_725_21.t12 Q.t4 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X25 VGND.t9 GATE_N.t1 a_27_47.t1 VNB.t12 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
R0 RESET_B.n0 RESET_B.t0 241.534
R1 RESET_B.n0 RESET_B.t1 169.234
R2 RESET_B RESET_B.n0 86.278
R3 a_725_21.n5 a_725_21.t4 368.328
R4 a_725_21.n3 a_725_21.t3 212.079
R5 a_725_21.n0 a_725_21.t12 212.079
R6 a_725_21.n1 a_725_21.t10 212.079
R7 a_725_21.n2 a_725_21.t6 212.079
R8 a_725_21.n4 a_725_21.t1 184.957
R9 a_725_21.n7 a_725_21.n6 152.768
R10 a_725_21.n5 a_725_21.t8 149.821
R11 a_725_21.n3 a_725_21.t9 139.779
R12 a_725_21.n0 a_725_21.t7 139.779
R13 a_725_21.n1 a_725_21.t11 139.779
R14 a_725_21.n2 a_725_21.t5 139.779
R15 a_725_21.n6 a_725_21.n5 111.684
R16 a_725_21.n6 a_725_21.n4 76.719
R17 a_725_21.n4 a_725_21.n3 76
R18 a_725_21.n1 a_725_21.n0 67.187
R19 a_725_21.n3 a_725_21.n2 66.457
R20 a_725_21.n2 a_725_21.n1 63.536
R21 a_725_21.n7 a_725_21.t2 26.595
R22 a_725_21.t0 a_725_21.n7 26.595
R23 VPWR.n15 VPWR.t1 578.851
R24 VPWR.n4 VPWR.t6 374.358
R25 VPWR.n28 VPWR.n27 311.893
R26 VPWR.n2 VPWR.n1 165.066
R27 VPWR.n13 VPWR.n12 161.588
R28 VPWR.n9 VPWR.t2 149.837
R29 VPWR.n8 VPWR.n7 124.033
R30 VPWR.n1 VPWR.t8 41.554
R31 VPWR.n1 VPWR.t0 41.554
R32 VPWR.n27 VPWR.t9 41.554
R33 VPWR.n27 VPWR.t10 41.554
R34 VPWR.n20 VPWR.n19 34.635
R35 VPWR.n21 VPWR.n20 34.635
R36 VPWR.n26 VPWR.n25 34.635
R37 VPWR.n12 VPWR.t5 32.505
R38 VPWR.n12 VPWR.t7 32.505
R39 VPWR.n7 VPWR.t4 29.55
R40 VPWR.n8 VPWR.n6 28.988
R41 VPWR.n19 VPWR.n4 28.235
R42 VPWR.n7 VPWR.t3 26.595
R43 VPWR.n25 VPWR.n2 26.352
R44 VPWR.n28 VPWR.n26 22.964
R45 VPWR.n14 VPWR.n13 21.458
R46 VPWR.n13 VPWR.n6 19.952
R47 VPWR.n21 VPWR.n2 19.2
R48 VPWR.n15 VPWR.n14 18.447
R49 VPWR.n15 VPWR.n4 14.305
R50 VPWR.n10 VPWR.n6 4.65
R51 VPWR.n13 VPWR.n11 4.65
R52 VPWR.n14 VPWR.n5 4.65
R53 VPWR.n16 VPWR.n15 4.65
R54 VPWR.n17 VPWR.n4 4.65
R55 VPWR.n19 VPWR.n18 4.65
R56 VPWR.n20 VPWR.n3 4.65
R57 VPWR.n22 VPWR.n21 4.65
R58 VPWR.n23 VPWR.n2 4.65
R59 VPWR.n25 VPWR.n24 4.65
R60 VPWR.n26 VPWR.n0 4.65
R61 VPWR.n29 VPWR.n28 3.932
R62 VPWR.n9 VPWR.n8 3.757
R63 VPWR.n10 VPWR.n9 0.258
R64 VPWR.n29 VPWR.n0 0.137
R65 VPWR.n11 VPWR.n10 0.119
R66 VPWR.n11 VPWR.n5 0.119
R67 VPWR.n16 VPWR.n5 0.119
R68 VPWR.n17 VPWR.n16 0.119
R69 VPWR.n18 VPWR.n17 0.119
R70 VPWR.n18 VPWR.n3 0.119
R71 VPWR.n22 VPWR.n3 0.119
R72 VPWR.n23 VPWR.n22 0.119
R73 VPWR.n24 VPWR.n23 0.119
R74 VPWR.n24 VPWR.n0 0.119
R75 VPWR VPWR.n29 0.101
R76 VPB.t11 VPB.t0 559.345
R77 VPB.t5 VPB.t1 556.386
R78 VPB.t2 VPB.t10 358.099
R79 VPB.t8 VPB.t7 284.112
R80 VPB.t9 VPB.t2 284.112
R81 VPB.t4 VPB.t3 272.274
R82 VPB.t7 VPB.t6 269.314
R83 VPB.t6 VPB.t4 257.476
R84 VPB.t1 VPB.t8 248.598
R85 VPB.t0 VPB.t9 248.598
R86 VPB.t12 VPB.t11 248.598
R87 VPB.t10 VPB.t5 213.084
R88 VPB VPB.t12 139.096
R89 a_300_47.n0 a_300_47.t3 373.281
R90 a_300_47.t0 a_300_47.n1 292.715
R91 a_300_47.n1 a_300_47.t1 182.645
R92 a_300_47.n0 a_300_47.t2 132.281
R93 a_300_47.n1 a_300_47.n0 80.46
R94 VGND.n2 VGND.t4 194.286
R95 VGND.n12 VGND.t6 148.331
R96 VGND.n1 VGND.n0 110.514
R97 VGND.n28 VGND.n27 107.239
R98 VGND.n21 VGND.n20 106.463
R99 VGND.n6 VGND.n5 106.052
R100 VGND.n20 VGND.t1 38.571
R101 VGND.n20 VGND.t0 38.571
R102 VGND.n27 VGND.t8 38.571
R103 VGND.n27 VGND.t9 38.571
R104 VGND.n5 VGND.t3 35.076
R105 VGND.n0 VGND.t5 27.692
R106 VGND.n5 VGND.t7 25.846
R107 VGND.n0 VGND.t2 24.923
R108 VGND.n4 VGND.n3 4.65
R109 VGND.n7 VGND.n6 4.65
R110 VGND.n9 VGND.n8 4.65
R111 VGND.n11 VGND.n10 4.65
R112 VGND.n13 VGND.n12 4.65
R113 VGND.n15 VGND.n14 4.65
R114 VGND.n17 VGND.n16 4.65
R115 VGND.n19 VGND.n18 4.65
R116 VGND.n22 VGND.n21 4.65
R117 VGND.n24 VGND.n23 4.65
R118 VGND.n26 VGND.n25 4.65
R119 VGND.n29 VGND.n28 3.932
R120 VGND.n2 VGND.n1 3.757
R121 VGND.n4 VGND.n2 0.258
R122 VGND.n29 VGND.n26 0.137
R123 VGND VGND.n29 0.121
R124 VGND.n7 VGND.n4 0.119
R125 VGND.n9 VGND.n7 0.119
R126 VGND.n11 VGND.n9 0.119
R127 VGND.n13 VGND.n11 0.119
R128 VGND.n15 VGND.n13 0.119
R129 VGND.n17 VGND.n15 0.119
R130 VGND.n19 VGND.n17 0.119
R131 VGND.n22 VGND.n19 0.119
R132 VGND.n24 VGND.n22 0.119
R133 VGND.n26 VGND.n24 0.119
R134 a_466_47.n0 a_466_47.t1 88.333
R135 a_466_47.n0 a_466_47.t0 26.393
R136 a_466_47.n1 a_466_47.n0 14.4
R137 VNB VNB.t12 6438.23
R138 VNB.t11 VNB.t0 6114.71
R139 VNB.t8 VNB.t1 5321.88
R140 VNB.t3 VNB.t10 3494.12
R141 VNB.t2 VNB.t8 3073.53
R142 VNB.t10 VNB.t2 2782.35
R143 VNB.t0 VNB.t3 2717.65
R144 VNB.t12 VNB.t11 2717.65
R145 VNB.t9 VNB.t5 2320.88
R146 VNB.t4 VNB.t6 2224.18
R147 VNB.t5 VNB.t7 2200
R148 VNB.t7 VNB.t4 2103.3
R149 VNB.t1 VNB.t9 2030.77
R150 a_27_47.t0 a_27_47.n3 269.575
R151 a_27_47.n1 a_27_47.t5 263.171
R152 a_27_47.n0 a_27_47.t4 240.108
R153 a_27_47.n0 a_27_47.t2 239.726
R154 a_27_47.n1 a_27_47.t3 227.825
R155 a_27_47.n2 a_27_47.t1 202.368
R156 a_27_47.n2 a_27_47.n1 76
R157 a_27_47.n3 a_27_47.n2 18.97
R158 a_27_47.n3 a_27_47.n0 11.272
R159 a_562_413.n3 a_562_413.n2 452.97
R160 a_562_413.n0 a_562_413.t4 221.719
R161 a_562_413.n2 a_562_413.n1 188.191
R162 a_562_413.n2 a_562_413.n0 178.019
R163 a_562_413.n0 a_562_413.t5 149.419
R164 a_562_413.n3 a_562_413.t2 121.952
R165 a_562_413.t0 a_562_413.n3 91.464
R166 a_562_413.n1 a_562_413.t3 46.666
R167 a_562_413.n1 a_562_413.t1 46.666
R168 Q Q.n3 300.359
R169 Q.n5 Q.n0 192.136
R170 Q.n4 Q.n2 118.089
R171 Q.n5 Q.n1 110.1
R172 Q.n4 Q 52.639
R173 Q.n3 Q.t6 30.535
R174 Q.n0 Q.t4 30.535
R175 Q.n0 Q.t5 30.535
R176 Q.n3 Q.t7 29.55
R177 Q.n2 Q.t1 29.538
R178 Q.n1 Q.t2 28.615
R179 Q.n1 Q.t0 28.615
R180 Q.n2 Q.t3 26.769
R181 Q Q.n5 9.6
R182 Q Q.n4 6.742
R183 Q.n5 Q 0.914
R184 a_660_47.t1 a_660_47.t0 93.059
R185 a_466_369.t1 a_466_369.t0 134.63
R186 GATE_N.n0 GATE_N.t0 269.919
R187 GATE_N.n0 GATE_N.t1 234.573
R188 GATE_N.n1 GATE_N.n0 76
R189 GATE_N GATE_N.n1 10.971
R190 GATE_N.n1 GATE_N 6.791
R191 D.n0 D.t0 327.642
R192 D.n0 D.t1 157.336
R193 D D.n0 78.594
R194 a_193_47.n0 a_193_47.t3 464.325
R195 a_193_47.n0 a_193_47.t2 242.606
R196 a_193_47.n1 a_193_47.t0 230.004
R197 a_193_47.t1 a_193_47.n1 121.759
R198 a_193_47.n1 a_193_47.n0 99.067
R199 a_683_413.t0 a_683_413.t1 98.5
R200 a_943_47.t0 a_943_47.t1 49.846
C0 VPB VPWR 0.16fF
C1 VGND Q 0.42fF
C2 VPWR Q 0.68fF
C3 VPWR VGND 0.13fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__dlrtp_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__dlrtp_1 RESET_B D GATE Q VGND VPWR VNB VPB
X0 a_929_47.t1 a_560_425.t4 a_711_21.t1 VNB.t6 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 VPWR.t1 D.t0 a_299_47.t0 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X2 Q.t1 a_711_21.t3 VPWR.t3 VPB.t6 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 a_465_47.t0 a_299_47.t2 VGND.t2 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 VGND.t4 a_711_21.t4 a_654_47.t1 VNB.t5 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 VPWR.t7 GATE.t0 a_27_47.t1 VPB.t9 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X6 Q.t0 a_711_21.t5 VGND.t3 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 a_560_425.t1 a_27_47.t2 a_465_369.t1 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X8 VPWR.t4 a_711_21.t6 a_664_425.t1 VPB.t5 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9 a_654_47.t0 a_27_47.t3 a_560_425.t2 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10 a_193_47.t0 a_27_47.t4 VGND.t5 VNB.t8 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11 a_711_21.t2 a_560_425.t5 VPWR.t5 VPB.t7 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 VPWR.t0 RESET_B.t0 a_711_21.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13 a_193_47.t1 a_27_47.t5 VPWR.t6 VPB.t8 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X14 a_560_425.t3 a_193_47.t2 a_465_47.t1 VNB.t7 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15 a_664_425.t0 a_193_47.t3 a_560_425.t0 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X16 VGND.t1 D.t1 a_299_47.t1 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17 VGND.t0 RESET_B.t1 a_929_47.t0 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X18 a_465_369.t0 a_299_47.t3 VPWR.t2 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X19 VGND.t6 GATE.t1 a_27_47.t0 VNB.t9 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
R0 a_560_425.n2 a_560_425.n0 427.064
R1 a_560_425.n1 a_560_425.t5 212.079
R2 a_560_425.n3 a_560_425.n2 190.004
R3 a_560_425.n2 a_560_425.n1 166.814
R4 a_560_425.n1 a_560_425.t4 139.779
R5 a_560_425.n0 a_560_425.t0 106.708
R6 a_560_425.n0 a_560_425.t1 95.763
R7 a_560_425.t2 a_560_425.n3 40
R8 a_560_425.n3 a_560_425.t3 40
R9 a_711_21.n1 a_711_21.t4 358.18
R10 a_711_21.n0 a_711_21.t3 241.534
R11 a_711_21.n0 a_711_21.t5 169.234
R12 a_711_21.n1 a_711_21.t6 149.821
R13 a_711_21.n4 a_711_21.n3 149.788
R14 a_711_21.n2 a_711_21.t1 129.861
R15 a_711_21.n3 a_711_21.n0 120.668
R16 a_711_21.n2 a_711_21.n1 97.348
R17 a_711_21.n4 a_711_21.t2 33.49
R18 a_711_21.t0 a_711_21.n4 31.52
R19 a_711_21.n3 a_711_21.n2 12.276
R20 a_929_47.t0 a_929_47.t1 60.923
R21 VNB.t8 VNB.t2 6082.35
R22 VNB.t5 VNB.t6 5321.88
R23 VNB VNB.t9 4270.59
R24 VNB.t1 VNB.t7 3332.35
R25 VNB.t3 VNB.t5 2814.71
R26 VNB.t7 VNB.t3 2782.35
R27 VNB.t2 VNB.t1 2717.65
R28 VNB.t9 VNB.t8 2717.65
R29 VNB.t6 VNB.t0 2320.88
R30 VNB.t0 VNB.t4 2224.18
R31 D.n0 D.t0 332.98
R32 D.n0 D.t1 156.248
R33 D D.n0 78.594
R34 a_299_47.n0 a_299_47.t3 373.281
R35 a_299_47.t0 a_299_47.n1 289.484
R36 a_299_47.n1 a_299_47.t1 178.929
R37 a_299_47.n0 a_299_47.t2 132.281
R38 a_299_47.n1 a_299_47.n0 81.236
R39 VPWR.n22 VPWR.n21 311.893
R40 VPWR.n5 VPWR.n4 292.5
R41 VPWR.n1 VPWR.n0 292.5
R42 VPWR.n3 VPWR.n2 167.784
R43 VPWR.n15 VPWR.n14 166.681
R44 VPWR.n4 VPWR.t4 63.321
R45 VPWR.n14 VPWR.t2 41.554
R46 VPWR.n14 VPWR.t1 41.554
R47 VPWR.n21 VPWR.t6 41.554
R48 VPWR.n21 VPWR.t7 41.554
R49 VPWR.n2 VPWR.t0 34.475
R50 VPWR.n0 VPWR.t5 29.315
R51 VPWR.n2 VPWR.t3 26.595
R52 VPWR.n7 VPWR.n6 4.65
R53 VPWR.n9 VPWR.n8 4.65
R54 VPWR.n11 VPWR.n10 4.65
R55 VPWR.n13 VPWR.n12 4.65
R56 VPWR.n16 VPWR.n15 4.65
R57 VPWR.n18 VPWR.n17 4.65
R58 VPWR.n20 VPWR.n19 4.65
R59 VPWR.n3 VPWR.n1 4.204
R60 VPWR.n23 VPWR.n22 3.932
R61 VPWR.n6 VPWR.n5 3.224
R62 VPWR.n7 VPWR.n3 0.205
R63 VPWR.n23 VPWR.n20 0.137
R64 VPWR VPWR.n23 0.123
R65 VPWR.n9 VPWR.n7 0.119
R66 VPWR.n11 VPWR.n9 0.119
R67 VPWR.n13 VPWR.n11 0.119
R68 VPWR.n16 VPWR.n13 0.119
R69 VPWR.n18 VPWR.n16 0.119
R70 VPWR.n20 VPWR.n18 0.119
R71 VPB.t8 VPB.t1 556.386
R72 VPB.t5 VPB.t7 449.844
R73 VPB.t2 VPB.t5 334.423
R74 VPB.t4 VPB.t2 307.788
R75 VPB.t7 VPB.t0 284.112
R76 VPB.t3 VPB.t4 281.152
R77 VPB.t0 VPB.t6 272.274
R78 VPB.t1 VPB.t3 248.598
R79 VPB.t9 VPB.t8 248.598
R80 VPB VPB.t9 142.056
R81 Q.n0 Q.t1 226.813
R82 Q.n1 Q.t0 117.423
R83 Q Q.n1 82.718
R84 Q Q.n0 8.551
R85 Q.n0 Q 7.973
R86 Q.n1 Q 6.961
R87 VGND.n1 VGND.t4 152.167
R88 VGND.n2 VGND.n0 121.005
R89 VGND.n17 VGND.n16 107.239
R90 VGND.n10 VGND.n9 106.463
R91 VGND.n9 VGND.t2 38.571
R92 VGND.n9 VGND.t1 38.571
R93 VGND.n16 VGND.t5 38.571
R94 VGND.n16 VGND.t6 38.571
R95 VGND.n0 VGND.t0 32.307
R96 VGND.n0 VGND.t3 24.923
R97 VGND.n4 VGND.n3 4.65
R98 VGND.n6 VGND.n5 4.65
R99 VGND.n8 VGND.n7 4.65
R100 VGND.n11 VGND.n10 4.65
R101 VGND.n13 VGND.n12 4.65
R102 VGND.n15 VGND.n14 4.65
R103 VGND.n2 VGND.n1 4.005
R104 VGND.n18 VGND.n17 3.932
R105 VGND.n4 VGND.n2 0.145
R106 VGND.n18 VGND.n15 0.137
R107 VGND VGND.n18 0.123
R108 VGND.n6 VGND.n4 0.119
R109 VGND.n8 VGND.n6 0.119
R110 VGND.n11 VGND.n8 0.119
R111 VGND.n13 VGND.n11 0.119
R112 VGND.n15 VGND.n13 0.119
R113 a_465_47.t0 a_465_47.t1 104.285
R114 a_654_47.t0 a_654_47.t1 81.428
R115 GATE.n0 GATE.t0 272.06
R116 GATE.n0 GATE.t1 236.714
R117 GATE.n1 GATE.n0 76
R118 GATE GATE.n1 11.2
R119 GATE.n1 GATE 6.933
R120 a_27_47.n0 a_27_47.t3 425.533
R121 a_27_47.t1 a_27_47.n3 264.681
R122 a_27_47.n1 a_27_47.t5 262.942
R123 a_27_47.n0 a_27_47.t2 228.464
R124 a_27_47.n1 a_27_47.t4 227.596
R125 a_27_47.n2 a_27_47.t0 201.541
R126 a_27_47.n2 a_27_47.n1 76
R127 a_27_47.n3 a_27_47.n2 18.97
R128 a_27_47.n3 a_27_47.n0 17.031
R129 a_465_369.t0 a_465_369.t1 147.92
R130 a_664_425.n0 a_664_425.t0 158.694
R131 a_664_425.n0 a_664_425.t1 43.328
R132 a_664_425.n1 a_664_425.n0 23.64
R133 a_193_47.n0 a_193_47.t2 258.779
R134 a_193_47.n1 a_193_47.t0 230.23
R135 a_193_47.n0 a_193_47.t3 214.611
R136 a_193_47.t1 a_193_47.n1 121.825
R137 a_193_47.n1 a_193_47.n0 11.187
R138 RESET_B.n0 RESET_B.t0 241.534
R139 RESET_B.n0 RESET_B.t1 169.234
R140 RESET_B.n1 RESET_B.n0 81.042
R141 RESET_B RESET_B.n1 12.8
R142 RESET_B.n1 RESET_B 4.46
C0 VPWR Q 0.11fF
C1 VPB VPWR 0.12fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__dlrtp_2.ext - technology: sky130A

.subckt sky130_fd_sc_hd__dlrtp_2 RESET_B Q D GATE VGND VPWR VNB VPB
X0 a_560_47.t0 a_193_47.t2 a_465_47.t0 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X1 VPWR.t6 D.t0 a_299_47.t1 VPB.t7 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X2 VPWR.t1 a_711_307.t3 a_644_413.t1 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3 a_465_47.t1 a_299_47.t2 VGND.t0 VNB.t10 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 VPWR.t8 GATE.t0 a_27_47.t1 VPB.t10 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X5 Q.t3 a_711_307.t4 VPWR.t2 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 VGND.t5 a_711_307.t5 a_657_47.t1 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7 a_657_47.t0 a_27_47.t2 a_560_47.t2 VNB.t5 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X8 VPWR.t3 a_711_307.t6 Q.t2 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 a_193_47.t0 a_27_47.t3 VGND.t3 VNB.t6 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10 Q.t1 a_711_307.t7 VGND.t7 VNB.t8 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 VPWR.t5 RESET_B.t0 a_711_307.t2 VPB.t6 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 a_940_47.t0 a_560_47.t4 a_711_307.t1 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 a_193_47.t1 a_27_47.t4 VPWR.t7 VPB.t8 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X14 VGND.t6 a_711_307.t8 Q.t0 VNB.t9 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X15 a_711_307.t0 a_560_47.t5 VPWR.t4 VPB.t5 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16 VGND.t2 D.t1 a_299_47.t0 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17 a_644_413.t0 a_193_47.t3 a_560_47.t1 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18 VGND.t1 RESET_B.t1 a_940_47.t1 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X19 a_465_369.t0 a_299_47.t3 VPWR.t0 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X20 a_560_47.t3 a_27_47.t5 a_465_369.t1 VPB.t9 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21 VGND.t4 GATE.t1 a_27_47.t0 VNB.t7 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
R0 a_193_47.n0 a_193_47.t2 267.083
R1 a_193_47.n1 a_193_47.t0 230.004
R2 a_193_47.n0 a_193_47.t3 222.644
R3 a_193_47.t1 a_193_47.n1 121.759
R4 a_193_47.n1 a_193_47.n0 12.512
R5 a_465_47.n0 a_465_47.t0 66.666
R6 a_465_47.n0 a_465_47.t1 26.393
R7 a_465_47.n1 a_465_47.n0 14.4
R8 a_560_47.n3 a_560_47.n2 415.873
R9 a_560_47.n0 a_560_47.t5 221.719
R10 a_560_47.n2 a_560_47.n0 187.328
R11 a_560_47.n2 a_560_47.n1 163.985
R12 a_560_47.n0 a_560_47.t4 149.419
R13 a_560_47.n1 a_560_47.t2 66.666
R14 a_560_47.t1 a_560_47.n3 63.321
R15 a_560_47.n3 a_560_47.t3 63.321
R16 a_560_47.n1 a_560_47.t0 45
R17 VNB VNB.t7 6438.23
R18 VNB.t6 VNB.t3 6082.35
R19 VNB.t1 VNB.t2 5321.88
R20 VNB.t0 VNB.t5 3138.24
R21 VNB.t5 VNB.t1 3073.53
R22 VNB.t10 VNB.t0 3073.53
R23 VNB.t3 VNB.t10 2717.65
R24 VNB.t7 VNB.t6 2717.65
R25 VNB.t2 VNB.t4 2272.53
R26 VNB.t4 VNB.t8 2200
R27 VNB.t8 VNB.t9 2030.77
R28 D.n0 D.t0 326.761
R29 D.n0 D.t1 156.455
R30 D D.n0 78.594
R31 a_299_47.n0 a_299_47.t3 373.281
R32 a_299_47.t1 a_299_47.n1 290.114
R33 a_299_47.n1 a_299_47.t0 179.635
R34 a_299_47.n0 a_299_47.t2 132.281
R35 a_299_47.n1 a_299_47.n0 81.042
R36 VPWR.n6 VPWR.t4 568.889
R37 VPWR.n8 VPWR.t1 370.126
R38 VPWR.n24 VPWR.n0 311.893
R39 VPWR.n3 VPWR.t3 260.943
R40 VPWR.n17 VPWR.n16 166.336
R41 VPWR.n2 VPWR.n1 162.694
R42 VPWR.n16 VPWR.t0 41.554
R43 VPWR.n16 VPWR.t6 41.554
R44 VPWR.n0 VPWR.t7 41.554
R45 VPWR.n0 VPWR.t8 41.554
R46 VPWR.n1 VPWR.t2 26.595
R47 VPWR.n1 VPWR.t5 26.595
R48 VPWR.n25 VPWR.n24 26.108
R49 VPWR.n24 VPWR.n23 4.65
R50 VPWR.n5 VPWR.n4 4.65
R51 VPWR.n7 VPWR.n6 4.65
R52 VPWR.n9 VPWR.n8 4.65
R53 VPWR.n11 VPWR.n10 4.65
R54 VPWR.n13 VPWR.n12 4.65
R55 VPWR.n15 VPWR.n14 4.65
R56 VPWR.n18 VPWR.n17 4.65
R57 VPWR.n20 VPWR.n19 4.65
R58 VPWR.n22 VPWR.n21 4.65
R59 VPWR.n3 VPWR.n2 3.778
R60 VPWR.n5 VPWR.n3 0.24
R61 VPWR.n7 VPWR.n5 0.119
R62 VPWR.n9 VPWR.n7 0.119
R63 VPWR.n11 VPWR.n9 0.119
R64 VPWR.n13 VPWR.n11 0.119
R65 VPWR.n15 VPWR.n13 0.119
R66 VPWR.n18 VPWR.n15 0.119
R67 VPWR.n20 VPWR.n18 0.119
R68 VPWR.n22 VPWR.n20 0.119
R69 VPWR.n23 VPWR.n22 0.119
R70 VPWR.n23 VPWR 0.118
R71 VPWR VPWR.n25 0.02
R72 VPWR.n25 VPWR 0.001
R73 VPB.t2 VPB.t5 588.94
R74 VPB.t8 VPB.t7 556.386
R75 VPB.t0 VPB.t2 287.071
R76 VPB.t1 VPB.t9 281.152
R77 VPB.t5 VPB.t6 278.193
R78 VPB.t3 VPB.t4 269.314
R79 VPB.t6 VPB.t3 248.598
R80 VPB.t9 VPB.t0 248.598
R81 VPB.t7 VPB.t1 248.598
R82 VPB.t10 VPB.t8 248.598
R83 VPB VPB.t10 139.096
R84 a_711_307.n4 a_711_307.t5 368.328
R85 a_711_307.n2 a_711_307.t4 214.269
R86 a_711_307.n0 a_711_307.t6 212.079
R87 a_711_307.n3 a_711_307.t1 176.282
R88 a_711_307.n6 a_711_307.n5 153.497
R89 a_711_307.n4 a_711_307.t3 149.821
R90 a_711_307.n0 a_711_307.t8 139.779
R91 a_711_307.n1 a_711_307.t7 139.779
R92 a_711_307.n5 a_711_307.n4 115.757
R93 a_711_307.n3 a_711_307.n2 76
R94 a_711_307.n5 a_711_307.n3 69.572
R95 a_711_307.n1 a_711_307.n0 61.345
R96 a_711_307.t0 a_711_307.n6 36.445
R97 a_711_307.n6 a_711_307.t2 26.595
R98 a_711_307.n2 a_711_307.n1 2.921
R99 a_644_413.t0 a_644_413.t1 157.13
R100 VGND.n0 VGND.t6 197.784
R101 VGND.n9 VGND.t5 147.823
R102 VGND.n2 VGND.n1 113.205
R103 VGND.n25 VGND.n24 107.239
R104 VGND.n18 VGND.n17 106.463
R105 VGND.n17 VGND.t0 38.571
R106 VGND.n17 VGND.t2 38.571
R107 VGND.n24 VGND.t3 38.571
R108 VGND.n24 VGND.t4 38.571
R109 VGND.n1 VGND.t1 31.384
R110 VGND.n1 VGND.t7 24.923
R111 VGND.n4 VGND.n3 4.65
R112 VGND.n6 VGND.n5 4.65
R113 VGND.n8 VGND.n7 4.65
R114 VGND.n10 VGND.n9 4.65
R115 VGND.n12 VGND.n11 4.65
R116 VGND.n14 VGND.n13 4.65
R117 VGND.n16 VGND.n15 4.65
R118 VGND.n19 VGND.n18 4.65
R119 VGND.n21 VGND.n20 4.65
R120 VGND.n23 VGND.n22 4.65
R121 VGND.n26 VGND.n25 3.932
R122 VGND.n3 VGND.n2 3.764
R123 VGND.n4 VGND.n0 0.746
R124 VGND.n26 VGND.n23 0.137
R125 VGND VGND.n26 0.121
R126 VGND.n6 VGND.n4 0.119
R127 VGND.n8 VGND.n6 0.119
R128 VGND.n10 VGND.n8 0.119
R129 VGND.n12 VGND.n10 0.119
R130 VGND.n14 VGND.n12 0.119
R131 VGND.n16 VGND.n14 0.119
R132 VGND.n19 VGND.n16 0.119
R133 VGND.n21 VGND.n19 0.119
R134 VGND.n23 VGND.n21 0.119
R135 GATE.n0 GATE.t0 270.454
R136 GATE.n0 GATE.t1 235.108
R137 GATE.n1 GATE.n0 76
R138 GATE GATE.n1 11.2
R139 GATE.n1 GATE 6.933
R140 a_27_47.n2 a_27_47.t2 441.612
R141 a_27_47.t1 a_27_47.n7 269.575
R142 a_27_47.n5 a_27_47.t4 263.171
R143 a_27_47.n1 a_27_47.t5 234.95
R144 a_27_47.n5 a_27_47.t3 227.825
R145 a_27_47.n6 a_27_47.t0 196.895
R146 a_27_47.n6 a_27_47.n5 76
R147 a_27_47.n7 a_27_47.n6 18.97
R148 a_27_47.n4 a_27_47.n3 14.412
R149 a_27_47.n3 a_27_47.n2 10.554
R150 a_27_47.n7 a_27_47.n4 9.726
R151 a_27_47.n4 a_27_47.n0 2.715
R152 a_27_47.n3 a_27_47.n1 1.417
R153 Q Q.n2 300.796
R154 Q.n1 Q.n0 146.59
R155 Q.n2 Q.t2 30.535
R156 Q.n2 Q.t3 29.55
R157 Q.n0 Q.t0 24.923
R158 Q.n0 Q.t1 24.923
R159 Q.n1 Q 11.52
R160 Q.n3 Q 4.828
R161 Q Q.n3 2.807
R162 Q.n1 Q 2.188
R163 Q.n3 Q.n1 0.547
R164 a_657_47.t1 a_657_47.t0 93.059
R165 RESET_B.n0 RESET_B.t0 240.999
R166 RESET_B.n0 RESET_B.t1 168.699
R167 RESET_B.n1 RESET_B.n0 86.372
R168 RESET_B.n1 RESET_B 2.865
R169 RESET_B RESET_B.n1 1.986
R170 a_940_47.t0 a_940_47.t1 59.076
R171 a_465_369.t0 a_465_369.t1 132.285
C0 VPB VPWR 0.14fF
C1 VPWR Q 0.27fF
C2 VPWR VGND 0.10fF
C3 VGND Q 0.20fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__dlrtp_4.ext - technology: sky130A

.subckt sky130_fd_sc_hd__dlrtp_4 GATE Q RESET_B D VGND VPWR VNB VPB
X0 VPWR.t9 RESET_B.t0 a_725_21.t0 VPB.t11 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_466_47.t0 a_300_47.t2 VGND.t0 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 a_562_413.t3 a_193_47.t2 a_466_47.t1 VNB.t9 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X3 Q.t3 a_725_21.t3 VPWR.t0 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 VGND.t1 a_725_21.t4 a_660_47.t0 VNB.t5 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 VGND.t5 a_725_21.t5 Q.t7 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 a_466_369.t0 a_300_47.t3 VPWR.t5 VPB.t5 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X7 VPWR.t7 GATE.t0 a_27_47.t0 VPB.t7 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X8 VPWR.t8 D.t0 a_300_47.t0 VPB.t10 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X9 VPWR.t4 a_725_21.t6 Q.t2 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 VGND.t4 a_725_21.t7 Q.t6 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 a_562_413.t1 a_27_47.t2 a_466_369.t1 VPB.t8 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12 a_725_21.t1 a_562_413.t4 VPWR.t10 VPB.t12 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13 a_193_47.t1 a_27_47.t3 VGND.t7 VNB.t8 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14 VPWR.t1 a_725_21.t8 a_683_413.t0 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15 a_943_47.t0 a_562_413.t5 a_725_21.t2 VNB.t12 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X16 Q.t5 a_725_21.t9 VGND.t3 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X17 Q.t1 a_725_21.t10 VPWR.t3 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X18 a_683_413.t1 a_193_47.t3 a_562_413.t2 VPB.t9 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19 a_193_47.t0 a_27_47.t4 VPWR.t6 VPB.t6 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X20 a_660_47.t1 a_27_47.t5 a_562_413.t0 VNB.t6 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X21 Q.t4 a_725_21.t11 VGND.t2 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X22 VGND.t8 D.t1 a_300_47.t1 VNB.t10 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23 VGND.t9 RESET_B.t1 a_943_47.t1 VNB.t11 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X24 VPWR.t2 a_725_21.t12 Q.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X25 VGND.t6 GATE.t1 a_27_47.t1 VNB.t7 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
R0 RESET_B.n0 RESET_B.t0 241.534
R1 RESET_B.n0 RESET_B.t1 169.234
R2 RESET_B RESET_B.n0 86.278
R3 a_725_21.n5 a_725_21.t4 368.328
R4 a_725_21.n3 a_725_21.t3 212.079
R5 a_725_21.n0 a_725_21.t12 212.079
R6 a_725_21.n1 a_725_21.t10 212.079
R7 a_725_21.n2 a_725_21.t6 212.079
R8 a_725_21.n4 a_725_21.t2 185.141
R9 a_725_21.n7 a_725_21.n6 152.768
R10 a_725_21.n5 a_725_21.t8 149.821
R11 a_725_21.n3 a_725_21.t9 139.779
R12 a_725_21.n0 a_725_21.t7 139.779
R13 a_725_21.n1 a_725_21.t11 139.779
R14 a_725_21.n2 a_725_21.t5 139.779
R15 a_725_21.n6 a_725_21.n5 111.684
R16 a_725_21.n6 a_725_21.n4 76.719
R17 a_725_21.n4 a_725_21.n3 76
R18 a_725_21.n1 a_725_21.n0 67.187
R19 a_725_21.n3 a_725_21.n2 66.457
R20 a_725_21.n2 a_725_21.n1 63.536
R21 a_725_21.t0 a_725_21.n7 26.595
R22 a_725_21.n7 a_725_21.t1 26.595
R23 VPWR.n15 VPWR.t10 578.851
R24 VPWR.n4 VPWR.t1 374.358
R25 VPWR.n28 VPWR.n27 311.893
R26 VPWR.n2 VPWR.n1 165.066
R27 VPWR.n13 VPWR.n12 161.588
R28 VPWR.n9 VPWR.t2 149.837
R29 VPWR.n8 VPWR.n7 124.033
R30 VPWR.n1 VPWR.t5 41.554
R31 VPWR.n1 VPWR.t8 41.554
R32 VPWR.n27 VPWR.t6 41.554
R33 VPWR.n27 VPWR.t7 41.554
R34 VPWR.n20 VPWR.n19 34.635
R35 VPWR.n21 VPWR.n20 34.635
R36 VPWR.n26 VPWR.n25 34.635
R37 VPWR.n12 VPWR.t0 32.505
R38 VPWR.n12 VPWR.t9 32.505
R39 VPWR.n7 VPWR.t4 29.55
R40 VPWR.n8 VPWR.n6 28.988
R41 VPWR.n19 VPWR.n4 28.235
R42 VPWR.n7 VPWR.t3 26.595
R43 VPWR.n25 VPWR.n2 26.352
R44 VPWR.n28 VPWR.n26 22.964
R45 VPWR.n14 VPWR.n13 21.458
R46 VPWR.n13 VPWR.n6 19.952
R47 VPWR.n21 VPWR.n2 19.2
R48 VPWR.n15 VPWR.n14 18.447
R49 VPWR.n15 VPWR.n4 14.305
R50 VPWR.n10 VPWR.n6 4.65
R51 VPWR.n13 VPWR.n11 4.65
R52 VPWR.n14 VPWR.n5 4.65
R53 VPWR.n16 VPWR.n15 4.65
R54 VPWR.n17 VPWR.n4 4.65
R55 VPWR.n19 VPWR.n18 4.65
R56 VPWR.n20 VPWR.n3 4.65
R57 VPWR.n22 VPWR.n21 4.65
R58 VPWR.n23 VPWR.n2 4.65
R59 VPWR.n25 VPWR.n24 4.65
R60 VPWR.n26 VPWR.n0 4.65
R61 VPWR.n29 VPWR.n28 3.932
R62 VPWR.n9 VPWR.n8 3.757
R63 VPWR.n10 VPWR.n9 0.258
R64 VPWR.n29 VPWR.n0 0.137
R65 VPWR.n11 VPWR.n10 0.119
R66 VPWR.n11 VPWR.n5 0.119
R67 VPWR.n16 VPWR.n5 0.119
R68 VPWR.n17 VPWR.n16 0.119
R69 VPWR.n18 VPWR.n17 0.119
R70 VPWR.n18 VPWR.n3 0.119
R71 VPWR.n22 VPWR.n3 0.119
R72 VPWR.n23 VPWR.n22 0.119
R73 VPWR.n24 VPWR.n23 0.119
R74 VPWR.n24 VPWR.n0 0.119
R75 VPWR VPWR.n29 0.101
R76 VPB.t6 VPB.t10 559.345
R77 VPB.t2 VPB.t12 556.386
R78 VPB.t8 VPB.t9 358.099
R79 VPB.t11 VPB.t4 284.112
R80 VPB.t5 VPB.t8 284.112
R81 VPB.t1 VPB.t0 272.274
R82 VPB.t4 VPB.t3 269.314
R83 VPB.t3 VPB.t1 257.476
R84 VPB.t12 VPB.t11 248.598
R85 VPB.t10 VPB.t5 248.598
R86 VPB.t7 VPB.t6 248.598
R87 VPB.t9 VPB.t2 213.084
R88 VPB VPB.t7 139.096
R89 a_300_47.n0 a_300_47.t3 373.281
R90 a_300_47.t0 a_300_47.n1 292.715
R91 a_300_47.n1 a_300_47.t1 182.645
R92 a_300_47.n0 a_300_47.t2 132.281
R93 a_300_47.n1 a_300_47.n0 80.46
R94 VGND.n2 VGND.t4 194.286
R95 VGND.n12 VGND.t1 148.331
R96 VGND.n1 VGND.n0 110.514
R97 VGND.n28 VGND.n27 107.239
R98 VGND.n21 VGND.n20 106.463
R99 VGND.n6 VGND.n5 106.052
R100 VGND.n20 VGND.t0 38.571
R101 VGND.n20 VGND.t8 38.571
R102 VGND.n27 VGND.t7 38.571
R103 VGND.n27 VGND.t6 38.571
R104 VGND.n5 VGND.t3 35.076
R105 VGND.n0 VGND.t5 27.692
R106 VGND.n5 VGND.t9 25.846
R107 VGND.n0 VGND.t2 24.923
R108 VGND.n4 VGND.n3 4.65
R109 VGND.n7 VGND.n6 4.65
R110 VGND.n9 VGND.n8 4.65
R111 VGND.n11 VGND.n10 4.65
R112 VGND.n13 VGND.n12 4.65
R113 VGND.n15 VGND.n14 4.65
R114 VGND.n17 VGND.n16 4.65
R115 VGND.n19 VGND.n18 4.65
R116 VGND.n22 VGND.n21 4.65
R117 VGND.n24 VGND.n23 4.65
R118 VGND.n26 VGND.n25 4.65
R119 VGND.n29 VGND.n28 3.932
R120 VGND.n2 VGND.n1 3.757
R121 VGND.n4 VGND.n2 0.258
R122 VGND.n29 VGND.n26 0.137
R123 VGND VGND.n29 0.121
R124 VGND.n7 VGND.n4 0.119
R125 VGND.n9 VGND.n7 0.119
R126 VGND.n11 VGND.n9 0.119
R127 VGND.n13 VGND.n11 0.119
R128 VGND.n15 VGND.n13 0.119
R129 VGND.n17 VGND.n15 0.119
R130 VGND.n19 VGND.n17 0.119
R131 VGND.n22 VGND.n19 0.119
R132 VGND.n24 VGND.n22 0.119
R133 VGND.n26 VGND.n24 0.119
R134 a_466_47.n0 a_466_47.t1 88.333
R135 a_466_47.n0 a_466_47.t0 26.393
R136 a_466_47.n1 a_466_47.n0 14.4
R137 VNB VNB.t7 6438.23
R138 VNB.t8 VNB.t10 6114.71
R139 VNB.t5 VNB.t12 5321.88
R140 VNB.t0 VNB.t9 3494.12
R141 VNB.t6 VNB.t5 3073.53
R142 VNB.t9 VNB.t6 2782.35
R143 VNB.t10 VNB.t0 2717.65
R144 VNB.t7 VNB.t8 2717.65
R145 VNB.t11 VNB.t2 2320.88
R146 VNB.t1 VNB.t3 2224.18
R147 VNB.t2 VNB.t4 2200
R148 VNB.t4 VNB.t1 2103.3
R149 VNB.t12 VNB.t11 2030.77
R150 a_193_47.n0 a_193_47.t2 255.425
R151 a_193_47.n1 a_193_47.t1 230.004
R152 a_193_47.n0 a_193_47.t3 172.23
R153 a_193_47.t0 a_193_47.n1 121.759
R154 a_193_47.n1 a_193_47.n0 6.548
R155 a_562_413.n3 a_562_413.n2 423.37
R156 a_562_413.n0 a_562_413.t4 221.719
R157 a_562_413.n2 a_562_413.n1 191.134
R158 a_562_413.n2 a_562_413.n0 185.309
R159 a_562_413.n0 a_562_413.t5 149.419
R160 a_562_413.t1 a_562_413.n3 121.952
R161 a_562_413.n3 a_562_413.t2 91.464
R162 a_562_413.n1 a_562_413.t0 46.666
R163 a_562_413.n1 a_562_413.t3 46.666
R164 Q Q.n3 300.359
R165 Q.n2 Q.n0 192.136
R166 Q.n5 Q.n4 118.089
R167 Q.n2 Q.n1 110.1
R168 Q.n5 Q 52.639
R169 Q.n0 Q.t0 30.535
R170 Q.n0 Q.t1 30.535
R171 Q.n3 Q.t2 30.535
R172 Q.n3 Q.t3 29.55
R173 Q.n4 Q.t5 29.538
R174 Q.n1 Q.t6 28.615
R175 Q.n1 Q.t4 28.615
R176 Q.n4 Q.t7 26.769
R177 Q.n2 Q 9.6
R178 Q Q.n5 6.742
R179 Q Q.n2 0.914
R180 a_660_47.t0 a_660_47.t1 93.059
R181 a_466_369.t0 a_466_369.t1 134.63
R182 GATE.n0 GATE.t0 269.919
R183 GATE.n0 GATE.t1 234.573
R184 GATE.n1 GATE.n0 76
R185 GATE GATE.n1 10.971
R186 GATE.n1 GATE 6.791
R187 a_27_47.n2 a_27_47.t5 450.47
R188 a_27_47.t0 a_27_47.n7 269.575
R189 a_27_47.n5 a_27_47.t4 263.171
R190 a_27_47.n1 a_27_47.t2 241
R191 a_27_47.n5 a_27_47.t3 227.825
R192 a_27_47.n6 a_27_47.t1 202.368
R193 a_27_47.n6 a_27_47.n5 76
R194 a_27_47.n7 a_27_47.n6 18.97
R195 a_27_47.n4 a_27_47.n3 15.872
R196 a_27_47.n3 a_27_47.n2 11.851
R197 a_27_47.n7 a_27_47.n4 9.609
R198 a_27_47.n4 a_27_47.n0 2.327
R199 a_27_47.n3 a_27_47.n1 1.606
R200 D.n0 D.t0 327.642
R201 D.n0 D.t1 157.336
R202 D D.n0 78.594
R203 a_683_413.t0 a_683_413.t1 98.5
R204 a_943_47.t0 a_943_47.t1 49.846
C0 VPB VPWR 0.16fF
C1 VGND Q 0.42fF
C2 VPWR Q 0.68fF
C3 VPWR VGND 0.13fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__dlxbn_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__dlxbn_1 Q_N D GATE_N Q VGND VPWR VNB VPB
X0 a_560_47.t0 a_27_47.t2 a_465_47.t0 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X1 a_560_47.t2 a_193_47.t2 a_470_369.t0 VPB.t8 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 a_465_47.t1 a_299_47.t2 VGND.t2 VNB.t10 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3 a_674_413.t0 a_27_47.t3 a_560_47.t1 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 VPWR.t6 a_716_21.t2 a_1124_47.t0 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X5 VPWR.t3 GATE_N.t0 a_27_47.t0 VPB.t6 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X6 VGND.t0 a_560_47.t4 a_716_21.t1 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 Q.t0 a_716_21.t3 VPWR.t7 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 a_193_47.t1 a_27_47.t4 VGND.t1 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9 a_651_47.t0 a_193_47.t3 a_560_47.t3 VNB.t9 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X10 Q.t1 a_716_21.t4 VGND.t3 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 Q_N.t0 a_1124_47.t2 VPWR.t4 VPB.t7 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 a_193_47.t0 a_27_47.t5 VPWR.t1 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X13 VPWR.t0 a_560_47.t5 a_716_21.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14 Q_N.t1 a_1124_47.t3 VGND.t8 VNB.t8 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X15 a_470_369.t1 a_299_47.t3 VPWR.t2 VPB.t10 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X16 VGND.t7 D.t0 a_299_47.t0 VNB.t7 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17 VGND.t4 a_716_21.t5 a_1124_47.t1 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18 VPWR.t5 D.t1 a_299_47.t1 VPB.t9 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X19 VPWR.t8 a_716_21.t6 a_674_413.t1 VPB.t5 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20 VGND.t5 a_716_21.t7 a_651_47.t1 VNB.t5 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21 VGND.t6 GATE_N.t1 a_27_47.t1 VNB.t6 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
R0 a_27_47.n0 a_27_47.t2 295.235
R1 a_27_47.t0 a_27_47.n3 269.575
R2 a_27_47.n1 a_27_47.t5 263.171
R3 a_27_47.n1 a_27_47.t4 227.825
R4 a_27_47.n0 a_27_47.t3 227.086
R5 a_27_47.n2 a_27_47.t1 202.368
R6 a_27_47.n2 a_27_47.n1 76
R7 a_27_47.n3 a_27_47.n2 18.97
R8 a_27_47.n3 a_27_47.n0 11.29
R9 a_465_47.n0 a_465_47.t0 66.666
R10 a_465_47.n0 a_465_47.t1 26.393
R11 a_465_47.n1 a_465_47.n0 14.4
R12 a_560_47.n3 a_560_47.n2 436.334
R13 a_560_47.n0 a_560_47.t5 212.079
R14 a_560_47.n2 a_560_47.n1 193.769
R15 a_560_47.n2 a_560_47.n0 165.045
R16 a_560_47.n0 a_560_47.t4 139.779
R17 a_560_47.n3 a_560_47.t2 119.607
R18 a_560_47.t1 a_560_47.n3 63.321
R19 a_560_47.n1 a_560_47.t0 51.666
R20 a_560_47.n1 a_560_47.t3 50
R21 VNB.t1 VNB.t7 6082.35
R22 VNB.t5 VNB.t0 5321.88
R23 VNB.t3 VNB.t4 4545.05
R24 VNB VNB.t6 4238.23
R25 VNB.t9 VNB.t5 3073.53
R26 VNB.t10 VNB.t2 3073.53
R27 VNB.t2 VNB.t9 2944.12
R28 VNB.t7 VNB.t10 2717.65
R29 VNB.t6 VNB.t1 2717.65
R30 VNB.t4 VNB.t8 2296.7
R31 VNB.t0 VNB.t3 2030.77
R32 a_193_47.n0 a_193_47.t3 562.709
R33 a_193_47.n1 a_193_47.t1 230.004
R34 a_193_47.n0 a_193_47.t2 219.041
R35 a_193_47.t0 a_193_47.n1 121.759
R36 a_193_47.n1 a_193_47.n0 99.085
R37 a_470_369.t1 a_470_369.t0 134.63
R38 VPB.t1 VPB.t9 571.183
R39 VPB.t4 VPB.t3 556.386
R40 VPB.t5 VPB.t0 556.386
R41 VPB.t8 VPB.t2 319.626
R42 VPB.t10 VPB.t8 284.112
R43 VPB.t3 VPB.t7 281.152
R44 VPB.t0 VPB.t4 248.598
R45 VPB.t9 VPB.t10 248.598
R46 VPB.t6 VPB.t1 248.598
R47 VPB.t2 VPB.t5 213.084
R48 VPB VPB.t6 139.096
R49 a_299_47.n0 a_299_47.t2 464.683
R50 a_299_47.n0 a_299_47.t3 328.294
R51 a_299_47.t1 a_299_47.n1 275.458
R52 a_299_47.n1 a_299_47.t0 188.354
R53 a_299_47.n1 a_299_47.n0 76
R54 VGND.n7 VGND.t5 148.331
R55 VGND.n4 VGND.n1 112.777
R56 VGND.n3 VGND.n2 107.239
R57 VGND.n23 VGND.n0 107.239
R58 VGND.n16 VGND.n15 105.48
R59 VGND.n1 VGND.t4 54.285
R60 VGND.n15 VGND.t2 38.571
R61 VGND.n15 VGND.t7 38.571
R62 VGND.n0 VGND.t1 38.571
R63 VGND.n0 VGND.t6 38.571
R64 VGND.n24 VGND.n23 26.108
R65 VGND.n1 VGND.t8 25.934
R66 VGND.n2 VGND.t3 24.923
R67 VGND.n2 VGND.t0 24.923
R68 VGND.n23 VGND.n22 4.65
R69 VGND.n6 VGND.n5 4.65
R70 VGND.n8 VGND.n7 4.65
R71 VGND.n10 VGND.n9 4.65
R72 VGND.n12 VGND.n11 4.65
R73 VGND.n14 VGND.n13 4.65
R74 VGND.n17 VGND.n16 4.65
R75 VGND.n19 VGND.n18 4.65
R76 VGND.n21 VGND.n20 4.65
R77 VGND.n4 VGND.n3 3.969
R78 VGND.n6 VGND.n4 0.146
R79 VGND.n8 VGND.n6 0.119
R80 VGND.n10 VGND.n8 0.119
R81 VGND.n12 VGND.n10 0.119
R82 VGND.n14 VGND.n12 0.119
R83 VGND.n17 VGND.n14 0.119
R84 VGND.n19 VGND.n17 0.119
R85 VGND.n21 VGND.n19 0.119
R86 VGND.n22 VGND.n21 0.119
R87 VGND.n22 VGND 0.118
R88 VGND VGND.n24 0.02
R89 VGND.n24 VGND 0.001
R90 a_674_413.t0 a_674_413.t1 98.5
R91 a_716_21.n4 a_716_21.t7 368.328
R92 a_716_21.n0 a_716_21.t2 268.364
R93 a_716_21.t0 a_716_21.n5 259.439
R94 a_716_21.n1 a_716_21.t3 212.079
R95 a_716_21.n0 a_716_21.t5 175.178
R96 a_716_21.n4 a_716_21.t6 149.821
R97 a_716_21.n3 a_716_21.t1 142.398
R98 a_716_21.n1 a_716_21.t4 139.779
R99 a_716_21.n2 a_716_21.n0 130.724
R100 a_716_21.n3 a_716_21.n2 98.109
R101 a_716_21.n5 a_716_21.n4 91.151
R102 a_716_21.n5 a_716_21.n3 61.211
R103 a_716_21.n2 a_716_21.n1 5.842
R104 a_1124_47.t0 a_1124_47.n1 377.062
R105 a_1124_47.n0 a_1124_47.t2 241.534
R106 a_1124_47.n0 a_1124_47.t3 169.234
R107 a_1124_47.n1 a_1124_47.t1 155.903
R108 a_1124_47.n1 a_1124_47.n0 98.69
R109 VPWR.n7 VPWR.t8 378.032
R110 VPWR.n24 VPWR.n0 311.893
R111 VPWR.n2 VPWR.n1 170.189
R112 VPWR.n4 VPWR.n3 170.127
R113 VPWR.n17 VPWR.n16 165.066
R114 VPWR.n3 VPWR.t6 58.484
R115 VPWR.n16 VPWR.t2 41.554
R116 VPWR.n16 VPWR.t5 41.554
R117 VPWR.n0 VPWR.t1 41.554
R118 VPWR.n0 VPWR.t3 41.554
R119 VPWR.n3 VPWR.t4 31.605
R120 VPWR.n1 VPWR.t7 26.595
R121 VPWR.n1 VPWR.t0 26.595
R122 VPWR.n25 VPWR.n24 26.108
R123 VPWR.n24 VPWR.n23 4.65
R124 VPWR.n6 VPWR.n5 4.65
R125 VPWR.n9 VPWR.n8 4.65
R126 VPWR.n11 VPWR.n10 4.65
R127 VPWR.n13 VPWR.n12 4.65
R128 VPWR.n15 VPWR.n14 4.65
R129 VPWR.n18 VPWR.n17 4.65
R130 VPWR.n20 VPWR.n19 4.65
R131 VPWR.n22 VPWR.n21 4.65
R132 VPWR.n4 VPWR.n2 3.969
R133 VPWR.n8 VPWR.n7 3.388
R134 VPWR.n6 VPWR.n4 0.146
R135 VPWR.n9 VPWR.n6 0.119
R136 VPWR.n11 VPWR.n9 0.119
R137 VPWR.n13 VPWR.n11 0.119
R138 VPWR.n15 VPWR.n13 0.119
R139 VPWR.n18 VPWR.n15 0.119
R140 VPWR.n20 VPWR.n18 0.119
R141 VPWR.n22 VPWR.n20 0.119
R142 VPWR.n23 VPWR.n22 0.119
R143 VPWR.n23 VPWR 0.118
R144 VPWR VPWR.n25 0.02
R145 VPWR.n25 VPWR 0.001
R146 GATE_N.n0 GATE_N.t0 270.454
R147 GATE_N.n0 GATE_N.t1 235.108
R148 GATE_N.n1 GATE_N.n0 76
R149 GATE_N GATE_N.n1 11.2
R150 GATE_N.n1 GATE_N 6.933
R151 Q.n0 Q.t0 227.256
R152 Q.n1 Q.t1 117.423
R153 Q Q.n1 80.187
R154 Q Q.n0 6.565
R155 Q.n0 Q 6.109
R156 Q.n1 Q 5.835
R157 a_651_47.t1 a_651_47.t0 93.059
R158 Q_N.n1 Q_N.t0 207.372
R159 Q_N.n0 Q_N.t1 117.423
R160 Q_N Q_N.n0 72.64
R161 Q_N.n1 Q_N 9.019
R162 Q_N Q_N.n1 7.458
R163 Q_N.n0 Q_N 6.646
R164 D.n0 D.t1 314.298
R165 D.n0 D.t0 157.542
R166 D D.n0 78.447
C0 VPWR Q_N 0.11fF
C1 VPWR Q 0.14fF
C2 VPWR VGND 0.11fF
C3 VPB VPWR 0.15fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__dlxbn_2.ext - technology: sky130A

.subckt sky130_fd_sc_hd__dlxbn_2 D GATE_N Q Q_N VPWR VGND VNB VPB
X0 VPWR.t8 a_728_21.t2 Q.t3 VPB.t9 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 VGND.t8 a_728_21.t3 a_663_47.t0 VNB.t9 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 VPWR.t5 a_728_21.t4 a_686_413.t1 VPB.t8 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3 Q_N.t1 a_1223_47.t2 VPWR.t3 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 VPWR.t0 GATE_N.t0 a_27_47.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X5 a_686_413.t0 a_27_47.t2 a_565_413.t0 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 VPWR.t4 a_1223_47.t3 Q_N.t0 VPB.t5 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 VGND.t7 a_728_21.t5 Q.t1 VNB.t8 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 Q.t2 a_728_21.t6 VPWR.t7 VPB.t7 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 VGND.t3 a_565_413.t4 a_728_21.t0 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 a_193_47.t1 a_27_47.t3 VGND.t4 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11 Q_N.t3 a_1223_47.t4 VGND.t1 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 VPWR.t6 a_728_21.t7 a_1223_47.t0 VPB.t6 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X13 a_663_47.t1 a_193_47.t2 a_565_413.t2 VNB.t12 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X14 VGND.t5 a_728_21.t8 a_1223_47.t1 VNB.t7 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15 a_469_369.t0 a_303_47.t2 VPWR.t10 VPB.t11 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X16 VGND.t10 D.t0 a_303_47.t0 VNB.t11 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17 a_193_47.t0 a_27_47.t4 VPWR.t2 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X18 VPWR.t9 D.t1 a_303_47.t1 VPB.t10 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X19 VGND.t2 a_1223_47.t5 Q_N.t2 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X20 a_565_413.t3 a_193_47.t3 a_469_369.t1 VPB.t12 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21 VPWR.t1 a_565_413.t5 a_728_21.t1 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X22 a_469_47.t1 a_303_47.t3 VGND.t9 VNB.t10 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23 a_565_413.t1 a_27_47.t5 a_469_47.t0 VNB.t5 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X24 VGND.t0 GATE_N.t1 a_27_47.t1 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X25 Q.t0 a_728_21.t9 VGND.t6 VNB.t6 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
R0 a_728_21.t1 a_728_21.n6 466.769
R1 a_728_21.n5 a_728_21.t3 368.328
R2 a_728_21.n0 a_728_21.t7 247.54
R3 a_728_21.n1 a_728_21.t2 212.079
R4 a_728_21.n2 a_728_21.t6 212.079
R5 a_728_21.n0 a_728_21.t8 154.354
R6 a_728_21.n5 a_728_21.t4 149.821
R7 a_728_21.n3 a_728_21.t0 144.477
R8 a_728_21.n1 a_728_21.t5 139.779
R9 a_728_21.n2 a_728_21.t9 139.779
R10 a_728_21.n1 a_728_21.n0 118.309
R11 a_728_21.n3 a_728_21.n2 100.686
R12 a_728_21.n6 a_728_21.n5 95.393
R13 a_728_21.n2 a_728_21.n1 61.345
R14 a_728_21.n4 a_728_21.n3 16.78
R15 a_728_21.n6 a_728_21.n4 0.969
R16 Q.n1 Q.n0 144.712
R17 Q.n3 Q.n2 92.5
R18 Q Q.n3 26.754
R19 Q.n0 Q.t3 26.595
R20 Q.n0 Q.t2 26.595
R21 Q.n2 Q.t1 24.923
R22 Q.n2 Q.t0 24.923
R23 Q Q.n1 9.7
R24 Q.n3 Q 7.936
R25 Q.n1 Q 7.346
R26 VPWR.n14 VPWR.t5 373.741
R27 VPWR.n30 VPWR.n29 311.893
R28 VPWR.n5 VPWR.t8 194.781
R29 VPWR.n10 VPWR.n9 169.982
R30 VPWR.n1 VPWR.n0 166.336
R31 VPWR.n23 VPWR.n22 165.066
R32 VPWR.n2 VPWR.t4 155.734
R33 VPWR.n0 VPWR.t6 58.484
R34 VPWR.n22 VPWR.t10 41.554
R35 VPWR.n22 VPWR.t9 41.554
R36 VPWR.n29 VPWR.t2 41.554
R37 VPWR.n29 VPWR.t0 41.554
R38 VPWR.n0 VPWR.t3 31.605
R39 VPWR.n9 VPWR.t1 29.55
R40 VPWR.n9 VPWR.t7 26.595
R41 VPWR.n4 VPWR.n3 4.65
R42 VPWR.n6 VPWR.n5 4.65
R43 VPWR.n8 VPWR.n7 4.65
R44 VPWR.n11 VPWR.n10 4.65
R45 VPWR.n13 VPWR.n12 4.65
R46 VPWR.n15 VPWR.n14 4.65
R47 VPWR.n17 VPWR.n16 4.65
R48 VPWR.n19 VPWR.n18 4.65
R49 VPWR.n21 VPWR.n20 4.65
R50 VPWR.n24 VPWR.n23 4.65
R51 VPWR.n26 VPWR.n25 4.65
R52 VPWR.n28 VPWR.n27 4.65
R53 VPWR.n31 VPWR.n30 3.932
R54 VPWR.n2 VPWR.n1 3.742
R55 VPWR.n4 VPWR.n2 0.245
R56 VPWR.n31 VPWR.n28 0.137
R57 VPWR VPWR.n31 0.123
R58 VPWR.n6 VPWR.n4 0.119
R59 VPWR.n8 VPWR.n6 0.119
R60 VPWR.n11 VPWR.n8 0.119
R61 VPWR.n13 VPWR.n11 0.119
R62 VPWR.n15 VPWR.n13 0.119
R63 VPWR.n17 VPWR.n15 0.119
R64 VPWR.n19 VPWR.n17 0.119
R65 VPWR.n21 VPWR.n19 0.119
R66 VPWR.n24 VPWR.n21 0.119
R67 VPWR.n26 VPWR.n24 0.119
R68 VPWR.n28 VPWR.n26 0.119
R69 VPB.t3 VPB.t10 568.224
R70 VPB.t9 VPB.t6 556.386
R71 VPB.t8 VPB.t1 556.386
R72 VPB.t12 VPB.t2 358.099
R73 VPB.t11 VPB.t12 284.112
R74 VPB.t6 VPB.t4 281.152
R75 VPB.t1 VPB.t7 257.476
R76 VPB.t4 VPB.t5 251.557
R77 VPB.t7 VPB.t9 248.598
R78 VPB.t10 VPB.t11 248.598
R79 VPB.t0 VPB.t3 248.598
R80 VPB.t2 VPB.t8 213.084
R81 VPB VPB.t0 192.367
R82 a_663_47.t0 a_663_47.t1 93.059
R83 VGND.n5 VGND.t7 193.59
R84 VGND.n14 VGND.t8 148.331
R85 VGND.n10 VGND.n9 117.201
R86 VGND.n2 VGND.t2 112.437
R87 VGND.n1 VGND.n0 108.988
R88 VGND.n30 VGND.n29 107.239
R89 VGND.n23 VGND.n22 106.463
R90 VGND.n0 VGND.t5 54.285
R91 VGND.n22 VGND.t9 38.571
R92 VGND.n22 VGND.t10 38.571
R93 VGND.n29 VGND.t4 38.571
R94 VGND.n29 VGND.t0 38.571
R95 VGND.n9 VGND.t3 27.692
R96 VGND.n0 VGND.t1 25.934
R97 VGND.n9 VGND.t6 24.923
R98 VGND.n4 VGND.n3 4.65
R99 VGND.n6 VGND.n5 4.65
R100 VGND.n8 VGND.n7 4.65
R101 VGND.n11 VGND.n10 4.65
R102 VGND.n13 VGND.n12 4.65
R103 VGND.n15 VGND.n14 4.65
R104 VGND.n17 VGND.n16 4.65
R105 VGND.n19 VGND.n18 4.65
R106 VGND.n21 VGND.n20 4.65
R107 VGND.n24 VGND.n23 4.65
R108 VGND.n26 VGND.n25 4.65
R109 VGND.n28 VGND.n27 4.65
R110 VGND.n31 VGND.n30 3.932
R111 VGND.n2 VGND.n1 3.742
R112 VGND.n4 VGND.n2 0.245
R113 VGND.n31 VGND.n28 0.137
R114 VGND VGND.n31 0.123
R115 VGND.n6 VGND.n4 0.119
R116 VGND.n8 VGND.n6 0.119
R117 VGND.n11 VGND.n8 0.119
R118 VGND.n13 VGND.n11 0.119
R119 VGND.n15 VGND.n13 0.119
R120 VGND.n17 VGND.n15 0.119
R121 VGND.n19 VGND.n17 0.119
R122 VGND.n21 VGND.n19 0.119
R123 VGND.n24 VGND.n21 0.119
R124 VGND.n26 VGND.n24 0.119
R125 VGND.n28 VGND.n26 0.119
R126 VNB VNB.t0 6470.59
R127 VNB.t4 VNB.t11 6211.76
R128 VNB.t9 VNB.t3 5321.88
R129 VNB.t8 VNB.t7 4545.05
R130 VNB.t10 VNB.t5 3494.12
R131 VNB.t12 VNB.t9 3073.53
R132 VNB.t5 VNB.t12 2782.35
R133 VNB.t11 VNB.t10 2717.65
R134 VNB.t0 VNB.t4 2717.65
R135 VNB.t7 VNB.t1 2296.7
R136 VNB.t3 VNB.t6 2103.3
R137 VNB.t1 VNB.t2 2054.95
R138 VNB.t6 VNB.t8 2030.77
R139 a_686_413.t0 a_686_413.t1 98.5
R140 a_1223_47.t0 a_1223_47.n2 240.007
R141 a_1223_47.n1 a_1223_47.t2 239.038
R142 a_1223_47.n0 a_1223_47.t3 221.719
R143 a_1223_47.n1 a_1223_47.t4 166.738
R144 a_1223_47.n2 a_1223_47.t1 149.883
R145 a_1223_47.n0 a_1223_47.t5 149.419
R146 a_1223_47.n2 a_1223_47.n1 99.272
R147 a_1223_47.n1 a_1223_47.n0 62.481
R148 Q_N.n4 Q_N.n3 142.958
R149 Q_N.n1 Q_N.n0 92.5
R150 Q_N.n3 Q_N.t0 27.58
R151 Q_N.n2 Q_N.n1 27.32
R152 Q_N.n3 Q_N.t1 26.595
R153 Q_N.n0 Q_N.t2 25.846
R154 Q_N.n0 Q_N.t3 24.923
R155 Q_N Q_N.n2 24.38
R156 Q_N.n2 Q_N 16.829
R157 Q_N.n4 Q_N 9.194
R158 Q_N Q_N.n4 7.483
R159 Q_N.n1 Q_N 6.776
R160 GATE_N.n0 GATE_N.t0 270.454
R161 GATE_N.n0 GATE_N.t1 235.108
R162 GATE_N.n1 GATE_N.n0 76
R163 GATE_N GATE_N.n1 10.971
R164 GATE_N.n1 GATE_N 6.791
R165 a_27_47.t0 a_27_47.n3 269.575
R166 a_27_47.n1 a_27_47.t4 263.171
R167 a_27_47.n0 a_27_47.t2 240.108
R168 a_27_47.n0 a_27_47.t5 239.726
R169 a_27_47.n1 a_27_47.t3 227.825
R170 a_27_47.n2 a_27_47.t1 202.368
R171 a_27_47.n2 a_27_47.n1 76
R172 a_27_47.n3 a_27_47.n2 18.97
R173 a_27_47.n3 a_27_47.n0 11.286
R174 a_565_413.n3 a_565_413.n2 422.17
R175 a_565_413.n0 a_565_413.t5 212.079
R176 a_565_413.n2 a_565_413.n1 190.005
R177 a_565_413.n2 a_565_413.n0 172.656
R178 a_565_413.n0 a_565_413.t4 139.779
R179 a_565_413.n3 a_565_413.t3 121.952
R180 a_565_413.t0 a_565_413.n3 91.464
R181 a_565_413.n1 a_565_413.t2 46.666
R182 a_565_413.n1 a_565_413.t1 46.666
R183 a_193_47.n0 a_193_47.t2 464.325
R184 a_193_47.n0 a_193_47.t3 242.606
R185 a_193_47.n1 a_193_47.t1 230.004
R186 a_193_47.t0 a_193_47.n1 121.759
R187 a_193_47.n1 a_193_47.n0 99.08
R188 a_303_47.n0 a_303_47.t2 373.281
R189 a_303_47.t1 a_303_47.n1 292.715
R190 a_303_47.n1 a_303_47.t0 182.645
R191 a_303_47.n0 a_303_47.t3 132.281
R192 a_303_47.n1 a_303_47.n0 80.46
R193 a_469_369.t0 a_469_369.t1 134.63
R194 D.n0 D.t1 327.642
R195 D.n0 D.t0 157.336
R196 D D.n0 78.594
R197 a_469_47.n0 a_469_47.t0 88.333
R198 a_469_47.n0 a_469_47.t1 26.393
R199 a_469_47.n1 a_469_47.n0 14.4
C0 VGND Q_N 0.20fF
C1 VGND Q 0.13fF
C2 VPWR Q_N 0.31fF
C3 VPWR Q 0.28fF
C4 VPWR VGND 0.14fF
C5 VPB VPWR 0.17fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__dlxbp_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__dlxbp_1 D GATE Q Q_N VGND VPWR VNB VPB
X0 a_560_47.t3 a_193_47.t2 a_465_47.t1 VNB.t8 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X1 a_465_47.t0 a_299_47.t2 VGND.t8 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 VPWR.t1 a_716_21.t2 a_1124_47.t0 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X3 VPWR.t3 GATE.t0 a_27_47.t0 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X4 a_467_369.t1 a_299_47.t3 VPWR.t8 VPB.t10 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X5 a_560_47.t0 a_27_47.t2 a_467_369.t0 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 VGND.t7 a_560_47.t4 a_716_21.t1 VNB.t10 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 VPWR.t5 D.t0 a_299_47.t0 VPB.t6 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X8 Q.t0 a_716_21.t3 VPWR.t0 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 a_193_47.t0 a_27_47.t3 VGND.t4 VNB.t5 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10 a_651_47.t0 a_27_47.t4 a_560_47.t1 VNB.t6 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X11 a_648_413.t1 a_193_47.t3 a_560_47.t2 VPB.t7 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12 Q.t1 a_716_21.t4 VGND.t1 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 Q_N.t0 a_1124_47.t2 VPWR.t6 VPB.t8 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14 a_193_47.t1 a_27_47.t5 VPWR.t4 VPB.t5 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X15 VPWR.t7 a_560_47.t5 a_716_21.t0 VPB.t9 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16 Q_N.t1 a_1124_47.t3 VGND.t6 VNB.t9 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X17 VGND.t5 D.t1 a_299_47.t1 VNB.t7 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18 VGND.t2 a_716_21.t5 a_1124_47.t1 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19 VPWR.t2 a_716_21.t6 a_648_413.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20 VGND.t3 a_716_21.t7 a_651_47.t1 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21 VGND.t0 GATE.t1 a_27_47.t1 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
R0 a_193_47.n0 a_193_47.t2 308.87
R1 a_193_47.n1 a_193_47.t0 230.004
R2 a_193_47.n0 a_193_47.t3 139.377
R3 a_193_47.t1 a_193_47.n1 121.759
R4 a_193_47.n1 a_193_47.n0 6.405
R5 a_465_47.n0 a_465_47.t1 66.666
R6 a_465_47.n0 a_465_47.t0 26.393
R7 a_465_47.n1 a_465_47.n0 14.4
R8 a_560_47.n3 a_560_47.n2 417.144
R9 a_560_47.n0 a_560_47.t5 212.079
R10 a_560_47.n2 a_560_47.n1 190.758
R11 a_560_47.n2 a_560_47.n0 170.465
R12 a_560_47.n0 a_560_47.t4 139.779
R13 a_560_47.n3 a_560_47.t2 65.666
R14 a_560_47.t0 a_560_47.n3 65.666
R15 a_560_47.n1 a_560_47.t3 56.666
R16 a_560_47.n1 a_560_47.t1 45
R17 VNB.t5 VNB.t7 6082.35
R18 VNB.t3 VNB.t10 5321.88
R19 VNB.t1 VNB.t2 4545.05
R20 VNB VNB.t0 4238.23
R21 VNB.t6 VNB.t3 3073.53
R22 VNB.t4 VNB.t8 3073.53
R23 VNB.t8 VNB.t6 2944.12
R24 VNB.t7 VNB.t4 2717.65
R25 VNB.t0 VNB.t5 2717.65
R26 VNB.t2 VNB.t9 2296.7
R27 VNB.t10 VNB.t1 2030.77
R28 a_299_47.n0 a_299_47.t3 328.294
R29 a_299_47.t0 a_299_47.n1 253.909
R30 a_299_47.n0 a_299_47.t2 177.268
R31 a_299_47.n1 a_299_47.t1 168.036
R32 a_299_47.n1 a_299_47.n0 76
R33 VGND.n6 VGND.t3 147.581
R34 VGND.n2 VGND.n1 120.66
R35 VGND.n3 VGND.n0 112.777
R36 VGND.n22 VGND.n21 107.239
R37 VGND.n15 VGND.n14 106.463
R38 VGND.n0 VGND.t2 54.285
R39 VGND.n14 VGND.t8 38.571
R40 VGND.n14 VGND.t5 38.571
R41 VGND.n21 VGND.t4 38.571
R42 VGND.n21 VGND.t0 38.571
R43 VGND.n0 VGND.t6 25.934
R44 VGND.n1 VGND.t1 24.923
R45 VGND.n1 VGND.t7 24.923
R46 VGND.n5 VGND.n4 4.65
R47 VGND.n7 VGND.n6 4.65
R48 VGND.n9 VGND.n8 4.65
R49 VGND.n11 VGND.n10 4.65
R50 VGND.n13 VGND.n12 4.65
R51 VGND.n16 VGND.n15 4.65
R52 VGND.n18 VGND.n17 4.65
R53 VGND.n20 VGND.n19 4.65
R54 VGND.n3 VGND.n2 3.969
R55 VGND.n23 VGND.n22 3.932
R56 VGND.n5 VGND.n3 0.146
R57 VGND.n23 VGND.n20 0.137
R58 VGND VGND.n23 0.121
R59 VGND.n7 VGND.n5 0.119
R60 VGND.n9 VGND.n7 0.119
R61 VGND.n11 VGND.n9 0.119
R62 VGND.n13 VGND.n11 0.119
R63 VGND.n16 VGND.n13 0.119
R64 VGND.n18 VGND.n16 0.119
R65 VGND.n20 VGND.n18 0.119
R66 a_716_21.t0 a_716_21.n6 466.769
R67 a_716_21.n5 a_716_21.t7 367.542
R68 a_716_21.n0 a_716_21.t2 261.885
R69 a_716_21.n1 a_716_21.t3 212.079
R70 a_716_21.n0 a_716_21.t5 168.699
R71 a_716_21.n5 a_716_21.t6 149.035
R72 a_716_21.n3 a_716_21.t1 141.001
R73 a_716_21.n1 a_716_21.t4 139.779
R74 a_716_21.n2 a_716_21.n0 125.612
R75 a_716_21.n3 a_716_21.n2 100.048
R76 a_716_21.n6 a_716_21.n5 94.618
R77 a_716_21.n4 a_716_21.n3 17.555
R78 a_716_21.n2 a_716_21.n1 7.303
R79 a_716_21.n6 a_716_21.n4 0.581
R80 a_1124_47.t0 a_1124_47.n1 377.062
R81 a_1124_47.n0 a_1124_47.t2 239.038
R82 a_1124_47.n0 a_1124_47.t3 166.738
R83 a_1124_47.n1 a_1124_47.t1 155.903
R84 a_1124_47.n1 a_1124_47.n0 97.721
R85 VPWR.n6 VPWR.t2 380.141
R86 VPWR.n22 VPWR.n21 311.893
R87 VPWR.n3 VPWR.n2 170.127
R88 VPWR.n1 VPWR.n0 169.982
R89 VPWR.n15 VPWR.n14 167.407
R90 VPWR.n2 VPWR.t1 58.484
R91 VPWR.n14 VPWR.t8 41.554
R92 VPWR.n14 VPWR.t5 41.554
R93 VPWR.n21 VPWR.t4 41.554
R94 VPWR.n21 VPWR.t3 41.554
R95 VPWR.n2 VPWR.t6 31.605
R96 VPWR.n0 VPWR.t0 26.595
R97 VPWR.n0 VPWR.t7 26.595
R98 VPWR.n5 VPWR.n4 4.65
R99 VPWR.n7 VPWR.n6 4.65
R100 VPWR.n9 VPWR.n8 4.65
R101 VPWR.n11 VPWR.n10 4.65
R102 VPWR.n13 VPWR.n12 4.65
R103 VPWR.n16 VPWR.n15 4.65
R104 VPWR.n18 VPWR.n17 4.65
R105 VPWR.n20 VPWR.n19 4.65
R106 VPWR.n3 VPWR.n1 3.969
R107 VPWR.n23 VPWR.n22 3.932
R108 VPWR.n5 VPWR.n3 0.146
R109 VPWR.n23 VPWR.n20 0.137
R110 VPWR VPWR.n23 0.121
R111 VPWR.n7 VPWR.n5 0.119
R112 VPWR.n9 VPWR.n7 0.119
R113 VPWR.n11 VPWR.n9 0.119
R114 VPWR.n13 VPWR.n11 0.119
R115 VPWR.n16 VPWR.n13 0.119
R116 VPWR.n18 VPWR.n16 0.119
R117 VPWR.n20 VPWR.n18 0.119
R118 VPB.t5 VPB.t6 562.305
R119 VPB.t1 VPB.t2 556.386
R120 VPB.t0 VPB.t9 556.386
R121 VPB.t7 VPB.t0 290.031
R122 VPB.t2 VPB.t8 281.152
R123 VPB.t10 VPB.t4 281.152
R124 VPB.t4 VPB.t7 254.517
R125 VPB.t9 VPB.t1 248.598
R126 VPB.t6 VPB.t10 248.598
R127 VPB.t3 VPB.t5 248.598
R128 VPB VPB.t3 139.096
R129 GATE.n0 GATE.t0 269.919
R130 GATE.n0 GATE.t1 234.573
R131 GATE.n1 GATE.n0 76
R132 GATE GATE.n1 10.971
R133 GATE.n1 GATE 6.791
R134 a_27_47.n0 a_27_47.t4 520.863
R135 a_27_47.t0 a_27_47.n3 269.575
R136 a_27_47.n1 a_27_47.t5 263.171
R137 a_27_47.n1 a_27_47.t3 227.825
R138 a_27_47.n0 a_27_47.t2 218.899
R139 a_27_47.n2 a_27_47.t1 202.368
R140 a_27_47.n2 a_27_47.n1 76
R141 a_27_47.n3 a_27_47.n2 18.97
R142 a_27_47.n3 a_27_47.n0 16.301
R143 a_467_369.t1 a_467_369.t0 132.285
R144 D.n0 D.t0 393.53
R145 D.n0 D.t1 215.79
R146 D D.n0 78.594
R147 Q.n0 Q.t0 227.297
R148 Q Q.t1 157.297
R149 Q Q.n0 6.38
R150 Q.n0 Q 5.935
R151 a_651_47.t1 a_651_47.t0 93.059
R152 a_648_413.t0 a_648_413.t1 159.476
R153 Q_N.n1 Q_N.t0 207.372
R154 Q_N.n0 Q_N.t1 117.423
R155 Q_N Q_N.n0 66.695
R156 Q_N.n1 Q_N 9.019
R157 Q_N Q_N.n1 7.458
R158 Q_N.n0 Q_N 6.646
C0 VPWR Q_N 0.11fF
C1 VGND Q 0.13fF
C2 VPWR Q 0.18fF
C3 VPWR VGND 0.11fF
C4 VPB VPWR 0.14fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__dlxtn_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__dlxtn_1 D GATE_N Q VGND VPWR VNB VPB
X0 a_560_47.t3 a_27_47.t2 a_465_47.t0 VNB.t7 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X1 VPWR.t6 D.t0 a_299_47.t1 VPB.t8 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X2 a_465_47.t1 a_299_47.t2 VGND.t1 VNB.t8 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3 VPWR.t4 GATE_N.t0 a_27_47.t0 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X4 VGND.t0 a_560_47.t4 a_715_21.t1 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 a_193_47.t1 a_27_47.t3 VGND.t5 VNB.t6 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 a_650_47.t0 a_193_47.t2 a_560_47.t0 VNB.t5 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X7 VPWR.t0 a_560_47.t5 a_715_21.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 Q.t0 a_715_21.t2 VPWR.t2 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 a_193_47.t0 a_27_47.t4 VPWR.t5 VPB.t7 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X10 VPWR.t3 a_715_21.t3 a_644_413.t0 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11 VGND.t6 D.t1 a_299_47.t0 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12 Q.t1 a_715_21.t4 VGND.t2 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 a_644_413.t1 a_27_47.t5 a_560_47.t2 VPB.t6 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14 a_465_369.t1 a_299_47.t3 VPWR.t1 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X15 a_560_47.t1 a_193_47.t3 a_465_369.t0 VPB.t5 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16 VGND.t4 GATE_N.t1 a_27_47.t1 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17 VGND.t3 a_715_21.t5 a_650_47.t1 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
R0 a_27_47.n0 a_27_47.t2 285.192
R1 a_27_47.t0 a_27_47.n3 269.575
R2 a_27_47.n1 a_27_47.t4 263.171
R3 a_27_47.n1 a_27_47.t3 227.825
R4 a_27_47.n0 a_27_47.t5 221.031
R5 a_27_47.n2 a_27_47.t1 202.368
R6 a_27_47.n2 a_27_47.n1 76
R7 a_27_47.n3 a_27_47.n2 18.97
R8 a_27_47.n3 a_27_47.n0 11.286
R9 a_465_47.n0 a_465_47.t0 66.666
R10 a_465_47.n0 a_465_47.t1 26.393
R11 a_465_47.n1 a_465_47.n0 14.4
R12 a_560_47.n3 a_560_47.n2 438.221
R13 a_560_47.n0 a_560_47.t5 212.079
R14 a_560_47.n2 a_560_47.n1 171.957
R15 a_560_47.n2 a_560_47.n0 167.681
R16 a_560_47.n0 a_560_47.t4 139.779
R17 a_560_47.n3 a_560_47.t2 63.321
R18 a_560_47.t1 a_560_47.n3 63.321
R19 a_560_47.n1 a_560_47.t0 55
R20 a_560_47.n1 a_560_47.t3 45
R21 VNB.t6 VNB.t1 6082.35
R22 VNB.t3 VNB.t0 5321.88
R23 VNB VNB.t4 4238.23
R24 VNB.t5 VNB.t3 3073.53
R25 VNB.t8 VNB.t7 3073.53
R26 VNB.t7 VNB.t5 2911.76
R27 VNB.t1 VNB.t8 2717.65
R28 VNB.t4 VNB.t6 2717.65
R29 VNB.t0 VNB.t2 2224.18
R30 D.n0 D.t0 344.36
R31 D.n0 D.t1 161.579
R32 D D.n0 78.594
R33 a_299_47.n0 a_299_47.t2 464.683
R34 a_299_47.n0 a_299_47.t3 328.294
R35 a_299_47.t1 a_299_47.n1 284.213
R36 a_299_47.n1 a_299_47.t0 184.2
R37 a_299_47.n1 a_299_47.n0 78.723
R38 VPWR.n0 VPWR.t3 371.021
R39 VPWR.n17 VPWR.n16 311.893
R40 VPWR.n2 VPWR.n1 173.582
R41 VPWR.n10 VPWR.n9 166.681
R42 VPWR.n9 VPWR.t1 41.554
R43 VPWR.n9 VPWR.t6 41.554
R44 VPWR.n16 VPWR.t5 41.554
R45 VPWR.n16 VPWR.t4 41.554
R46 VPWR.n1 VPWR.t0 34.475
R47 VPWR.n1 VPWR.t2 26.595
R48 VPWR.n4 VPWR.n3 4.65
R49 VPWR.n6 VPWR.n5 4.65
R50 VPWR.n8 VPWR.n7 4.65
R51 VPWR.n11 VPWR.n10 4.65
R52 VPWR.n13 VPWR.n12 4.65
R53 VPWR.n15 VPWR.n14 4.65
R54 VPWR.n18 VPWR.n17 3.932
R55 VPWR.n2 VPWR.n0 3.814
R56 VPWR.n4 VPWR.n2 0.223
R57 VPWR.n18 VPWR.n15 0.137
R58 VPWR VPWR.n18 0.121
R59 VPWR.n6 VPWR.n4 0.119
R60 VPWR.n8 VPWR.n6 0.119
R61 VPWR.n11 VPWR.n8 0.119
R62 VPWR.n13 VPWR.n11 0.119
R63 VPWR.n15 VPWR.n13 0.119
R64 VPB.t3 VPB.t0 556.386
R65 VPB.t7 VPB.t8 556.386
R66 VPB.t6 VPB.t3 298.909
R67 VPB.t1 VPB.t5 281.152
R68 VPB.t0 VPB.t2 272.274
R69 VPB.t5 VPB.t6 248.598
R70 VPB.t8 VPB.t1 248.598
R71 VPB.t4 VPB.t7 248.598
R72 VPB VPB.t4 139.096
R73 VGND.n1 VGND.t3 149.085
R74 VGND.n2 VGND.n0 127.472
R75 VGND.n17 VGND.n16 107.239
R76 VGND.n10 VGND.n9 106.463
R77 VGND.n9 VGND.t1 38.571
R78 VGND.n9 VGND.t6 38.571
R79 VGND.n16 VGND.t5 38.571
R80 VGND.n16 VGND.t4 38.571
R81 VGND.n0 VGND.t0 32.307
R82 VGND.n0 VGND.t2 24.923
R83 VGND.n4 VGND.n3 4.65
R84 VGND.n6 VGND.n5 4.65
R85 VGND.n8 VGND.n7 4.65
R86 VGND.n11 VGND.n10 4.65
R87 VGND.n13 VGND.n12 4.65
R88 VGND.n15 VGND.n14 4.65
R89 VGND.n18 VGND.n17 3.932
R90 VGND.n2 VGND.n1 3.914
R91 VGND.n4 VGND.n2 0.207
R92 VGND.n18 VGND.n15 0.137
R93 VGND VGND.n18 0.121
R94 VGND.n6 VGND.n4 0.119
R95 VGND.n8 VGND.n6 0.119
R96 VGND.n11 VGND.n8 0.119
R97 VGND.n13 VGND.n11 0.119
R98 VGND.n15 VGND.n13 0.119
R99 GATE_N.n0 GATE_N.t0 269.919
R100 GATE_N.n0 GATE_N.t1 234.573
R101 GATE_N.n1 GATE_N.n0 76
R102 GATE_N GATE_N.n1 10.971
R103 GATE_N.n1 GATE_N 6.791
R104 a_715_21.t0 a_715_21.n4 466.769
R105 a_715_21.n3 a_715_21.t5 367.542
R106 a_715_21.n0 a_715_21.t2 239.038
R107 a_715_21.n0 a_715_21.t4 166.738
R108 a_715_21.n1 a_715_21.t1 153.54
R109 a_715_21.n3 a_715_21.t3 149.035
R110 a_715_21.n1 a_715_21.n0 97.527
R111 a_715_21.n4 a_715_21.n3 94.618
R112 a_715_21.n2 a_715_21.n1 17.362
R113 a_715_21.n4 a_715_21.n2 1.357
R114 a_193_47.n0 a_193_47.t2 562.709
R115 a_193_47.n1 a_193_47.t1 230.004
R116 a_193_47.n0 a_193_47.t3 219.041
R117 a_193_47.t0 a_193_47.n1 121.759
R118 a_193_47.n1 a_193_47.n0 96.694
R119 a_650_47.t1 a_650_47.t0 93.059
R120 Q.n0 Q.t0 226.813
R121 Q.n1 Q.t1 117.423
R122 Q Q.n1 83.431
R123 Q Q.n0 8.551
R124 Q.n0 Q 7.973
R125 Q.n1 Q 7.63
R126 a_644_413.t0 a_644_413.t1 166.511
R127 a_465_369.t1 a_465_369.t0 132.285
C0 VPB VPWR 0.12fF
C1 Q VPWR 0.16fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__dlxtn_2.ext - technology: sky130A

.subckt sky130_fd_sc_hd__dlxtn_2 D GATE_N Q VPWR VGND VNB VPB
X0 VPWR.t1 a_728_21.t2 Q.t3 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 VGND.t0 a_728_21.t3 a_663_47.t0 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 VPWR.t2 a_728_21.t4 a_686_413.t0 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3 VPWR.t5 GATE_N.t0 a_27_47.t1 VPB.t5 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X4 a_686_413.t1 a_27_47.t2 a_565_413.t0 VPB.t6 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 VGND.t2 a_728_21.t5 Q.t1 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 Q.t2 a_728_21.t6 VPWR.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 VGND.t4 a_565_413.t4 a_728_21.t0 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 a_193_47.t0 a_27_47.t3 VGND.t5 VNB.t5 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9 a_663_47.t1 a_193_47.t2 a_565_413.t2 VNB.t9 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X10 a_469_369.t1 a_303_47.t2 VPWR.t7 VPB.t8 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X11 VGND.t3 D.t0 a_303_47.t0 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12 a_193_47.t1 a_27_47.t4 VPWR.t6 VPB.t7 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X13 VPWR.t3 D.t1 a_303_47.t1 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X14 a_565_413.t3 a_193_47.t3 a_469_369.t0 VPB.t9 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15 VPWR.t4 a_565_413.t5 a_728_21.t1 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16 a_469_47.t1 a_303_47.t3 VGND.t6 VNB.t7 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17 a_565_413.t1 a_27_47.t5 a_469_47.t0 VNB.t6 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X18 VGND.t7 GATE_N.t1 a_27_47.t0 VNB.t8 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19 Q.t0 a_728_21.t7 VGND.t1 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
R0 a_728_21.t1 a_728_21.n5 466.769
R1 a_728_21.n4 a_728_21.t3 368.328
R2 a_728_21.n0 a_728_21.t2 212.079
R3 a_728_21.n1 a_728_21.t6 212.079
R4 a_728_21.n4 a_728_21.t4 149.821
R5 a_728_21.n2 a_728_21.t0 144.477
R6 a_728_21.n0 a_728_21.t5 139.779
R7 a_728_21.n1 a_728_21.t7 139.779
R8 a_728_21.n2 a_728_21.n1 100.686
R9 a_728_21.n5 a_728_21.n4 95.393
R10 a_728_21.n1 a_728_21.n0 61.345
R11 a_728_21.n3 a_728_21.n2 16.78
R12 a_728_21.n5 a_728_21.n3 0.969
R13 Q.n1 Q.n0 144.712
R14 Q.n3 Q.n2 92.5
R15 Q Q.n3 26.955
R16 Q.n0 Q.t3 26.595
R17 Q.n0 Q.t2 26.595
R18 Q.n2 Q.t1 24.923
R19 Q.n2 Q.t0 24.923
R20 Q Q.n1 9.7
R21 Q.n3 Q 7.936
R22 Q.n1 Q 7.346
R23 VPWR.n5 VPWR.t2 373.741
R24 VPWR.n21 VPWR.n20 311.893
R25 VPWR.n2 VPWR.t1 199.721
R26 VPWR.n1 VPWR.n0 169.982
R27 VPWR.n14 VPWR.n13 165.066
R28 VPWR.n13 VPWR.t7 41.554
R29 VPWR.n13 VPWR.t3 41.554
R30 VPWR.n20 VPWR.t6 41.554
R31 VPWR.n20 VPWR.t5 41.554
R32 VPWR.n0 VPWR.t4 29.55
R33 VPWR.n0 VPWR.t0 26.595
R34 VPWR.n4 VPWR.n3 4.65
R35 VPWR.n6 VPWR.n5 4.65
R36 VPWR.n8 VPWR.n7 4.65
R37 VPWR.n10 VPWR.n9 4.65
R38 VPWR.n12 VPWR.n11 4.65
R39 VPWR.n15 VPWR.n14 4.65
R40 VPWR.n17 VPWR.n16 4.65
R41 VPWR.n19 VPWR.n18 4.65
R42 VPWR.n22 VPWR.n21 3.932
R43 VPWR.n2 VPWR.n1 3.73
R44 VPWR.n4 VPWR.n2 0.247
R45 VPWR.n22 VPWR.n19 0.137
R46 VPWR VPWR.n22 0.121
R47 VPWR.n6 VPWR.n4 0.119
R48 VPWR.n8 VPWR.n6 0.119
R49 VPWR.n10 VPWR.n8 0.119
R50 VPWR.n12 VPWR.n10 0.119
R51 VPWR.n15 VPWR.n12 0.119
R52 VPWR.n17 VPWR.n15 0.119
R53 VPWR.n19 VPWR.n17 0.119
R54 VPB.t7 VPB.t3 568.224
R55 VPB.t1 VPB.t4 556.386
R56 VPB.t9 VPB.t6 358.099
R57 VPB.t8 VPB.t9 284.112
R58 VPB.t4 VPB.t0 257.476
R59 VPB.t0 VPB.t2 248.598
R60 VPB.t3 VPB.t8 248.598
R61 VPB.t5 VPB.t7 248.598
R62 VPB.t6 VPB.t1 213.084
R63 VPB VPB.t5 189.408
R64 a_663_47.t0 a_663_47.t1 93.059
R65 VGND.n2 VGND.t2 198.383
R66 VGND.n5 VGND.t0 148.331
R67 VGND.n1 VGND.n0 117.201
R68 VGND.n21 VGND.n20 107.239
R69 VGND.n14 VGND.n13 106.463
R70 VGND.n13 VGND.t6 38.571
R71 VGND.n13 VGND.t3 38.571
R72 VGND.n20 VGND.t5 38.571
R73 VGND.n20 VGND.t7 38.571
R74 VGND.n0 VGND.t4 27.692
R75 VGND.n0 VGND.t1 24.923
R76 VGND.n4 VGND.n3 4.65
R77 VGND.n6 VGND.n5 4.65
R78 VGND.n8 VGND.n7 4.65
R79 VGND.n10 VGND.n9 4.65
R80 VGND.n12 VGND.n11 4.65
R81 VGND.n15 VGND.n14 4.65
R82 VGND.n17 VGND.n16 4.65
R83 VGND.n19 VGND.n18 4.65
R84 VGND.n22 VGND.n21 3.932
R85 VGND.n2 VGND.n1 3.73
R86 VGND.n4 VGND.n2 0.247
R87 VGND.n22 VGND.n19 0.137
R88 VGND VGND.n22 0.121
R89 VGND.n6 VGND.n4 0.119
R90 VGND.n8 VGND.n6 0.119
R91 VGND.n10 VGND.n8 0.119
R92 VGND.n12 VGND.n10 0.119
R93 VGND.n15 VGND.n12 0.119
R94 VGND.n17 VGND.n15 0.119
R95 VGND.n19 VGND.n17 0.119
R96 VNB VNB.t8 6438.23
R97 VNB.t5 VNB.t3 6211.76
R98 VNB.t2 VNB.t4 5321.88
R99 VNB.t7 VNB.t6 3494.12
R100 VNB.t9 VNB.t2 3073.53
R101 VNB.t6 VNB.t9 2782.35
R102 VNB.t3 VNB.t7 2717.65
R103 VNB.t8 VNB.t5 2717.65
R104 VNB.t4 VNB.t0 2103.3
R105 VNB.t0 VNB.t1 2030.77
R106 a_686_413.t0 a_686_413.t1 98.5
R107 GATE_N.n0 GATE_N.t0 269.919
R108 GATE_N.n0 GATE_N.t1 234.573
R109 GATE_N.n1 GATE_N.n0 76
R110 GATE_N GATE_N.n1 10.971
R111 GATE_N.n1 GATE_N 6.791
R112 a_27_47.t1 a_27_47.n3 269.575
R113 a_27_47.n1 a_27_47.t4 263.171
R114 a_27_47.n0 a_27_47.t2 240.108
R115 a_27_47.n0 a_27_47.t5 239.726
R116 a_27_47.n1 a_27_47.t3 227.825
R117 a_27_47.n2 a_27_47.t0 202.368
R118 a_27_47.n2 a_27_47.n1 76
R119 a_27_47.n3 a_27_47.n2 18.97
R120 a_27_47.n3 a_27_47.n0 11.286
R121 a_565_413.n3 a_565_413.n2 422.17
R122 a_565_413.n0 a_565_413.t5 212.079
R123 a_565_413.n2 a_565_413.n1 190.005
R124 a_565_413.n2 a_565_413.n0 172.656
R125 a_565_413.n0 a_565_413.t4 139.779
R126 a_565_413.n3 a_565_413.t3 121.952
R127 a_565_413.t0 a_565_413.n3 91.464
R128 a_565_413.n1 a_565_413.t2 46.666
R129 a_565_413.n1 a_565_413.t1 46.666
R130 a_193_47.n0 a_193_47.t2 464.325
R131 a_193_47.n0 a_193_47.t3 242.606
R132 a_193_47.n1 a_193_47.t0 230.004
R133 a_193_47.t1 a_193_47.n1 121.759
R134 a_193_47.n1 a_193_47.n0 99.08
R135 a_303_47.n0 a_303_47.t2 373.281
R136 a_303_47.t1 a_303_47.n1 292.715
R137 a_303_47.n1 a_303_47.t0 182.645
R138 a_303_47.n0 a_303_47.t3 132.281
R139 a_303_47.n1 a_303_47.n0 80.46
R140 a_469_369.t1 a_469_369.t0 134.63
R141 D.n0 D.t1 327.642
R142 D.n0 D.t0 157.336
R143 D D.n0 78.594
R144 a_469_47.n0 a_469_47.t0 88.333
R145 a_469_47.n0 a_469_47.t1 26.393
R146 a_469_47.n1 a_469_47.n0 14.4
C0 VGND Q 0.13fF
C1 VPWR Q 0.29fF
C2 VPB VPWR 0.13fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__dlxtn_4.ext - technology: sky130A

.subckt sky130_fd_sc_hd__dlxtn_4 D GATE_N Q VPWR VGND VNB VPB
X0 VPWR.t0 D.t0 a_299_47.t0 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1 Q.t4 a_724_21.t2 VPWR.t5 VPB.t7 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 a_561_413.t2 a_27_47.t2 a_465_47.t0 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X3 a_465_47.t1 a_299_47.t2 VGND.t3 VNB.t5 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 a_561_413.t0 a_193_47.t2 a_465_369.t1 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 VGND.t8 a_724_21.t3 a_659_47.t0 VNB.t10 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 Q.t0 a_724_21.t4 VGND.t7 VNB.t9 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 VPWR.t1 GATE_N.t0 a_27_47.t0 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X8 a_659_47.t1 a_193_47.t3 a_561_413.t3 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X9 Q.t3 a_724_21.t5 VPWR.t6 VPB.t8 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 VPWR.t7 a_724_21.t6 a_682_413.t1 VPB.t9 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11 a_193_47.t0 a_27_47.t3 VGND.t2 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12 a_682_413.t0 a_27_47.t4 a_561_413.t1 VPB.t5 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13 VPWR.t8 a_724_21.t7 Q.t2 VPB.t10 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14 VGND.t6 a_724_21.t8 Q.t7 VNB.t8 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X15 a_193_47.t1 a_27_47.t5 VPWR.t4 VPB.t6 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X16 VPWR.t2 a_561_413.t4 a_724_21.t0 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17 VGND.t9 a_561_413.t5 a_724_21.t1 VNB.t11 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X18 VGND.t5 a_724_21.t9 Q.t6 VNB.t7 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X19 Q.t5 a_724_21.t10 VGND.t4 VNB.t6 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X20 VGND.t0 D.t1 a_299_47.t1 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21 VPWR.t9 a_724_21.t11 Q.t1 VPB.t11 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X22 a_465_369.t0 a_299_47.t3 VPWR.t3 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X23 VGND.t1 GATE_N.t1 a_27_47.t1 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
R0 D.n0 D.t0 327.642
R1 D.n0 D.t1 157.336
R2 D D.n0 78.594
R3 a_299_47.n0 a_299_47.t3 373.281
R4 a_299_47.t0 a_299_47.n1 292.715
R5 a_299_47.n1 a_299_47.t1 182.645
R6 a_299_47.n0 a_299_47.t2 132.281
R7 a_299_47.n1 a_299_47.n0 80.46
R8 VPWR.n10 VPWR.t7 373.741
R9 VPWR.n26 VPWR.n25 311.893
R10 VPWR.n2 VPWR.t8 260.943
R11 VPWR.n1 VPWR.n0 173.868
R12 VPWR.n6 VPWR.n5 169.982
R13 VPWR.n19 VPWR.n18 165.066
R14 VPWR.n18 VPWR.t3 41.554
R15 VPWR.n18 VPWR.t0 41.554
R16 VPWR.n25 VPWR.t4 41.554
R17 VPWR.n25 VPWR.t1 41.554
R18 VPWR.n0 VPWR.t9 33.49
R19 VPWR.n5 VPWR.t2 29.55
R20 VPWR.n0 VPWR.t5 26.595
R21 VPWR.n5 VPWR.t6 26.595
R22 VPWR.n4 VPWR.n3 4.65
R23 VPWR.n7 VPWR.n6 4.65
R24 VPWR.n9 VPWR.n8 4.65
R25 VPWR.n11 VPWR.n10 4.65
R26 VPWR.n13 VPWR.n12 4.65
R27 VPWR.n15 VPWR.n14 4.65
R28 VPWR.n17 VPWR.n16 4.65
R29 VPWR.n20 VPWR.n19 4.65
R30 VPWR.n22 VPWR.n21 4.65
R31 VPWR.n24 VPWR.n23 4.65
R32 VPWR.n27 VPWR.n26 3.932
R33 VPWR.n2 VPWR.n1 3.778
R34 VPWR.n4 VPWR.n2 0.24
R35 VPWR.n27 VPWR.n24 0.137
R36 VPWR VPWR.n27 0.123
R37 VPWR.n7 VPWR.n4 0.119
R38 VPWR.n9 VPWR.n7 0.119
R39 VPWR.n11 VPWR.n9 0.119
R40 VPWR.n13 VPWR.n11 0.119
R41 VPWR.n15 VPWR.n13 0.119
R42 VPWR.n17 VPWR.n15 0.119
R43 VPWR.n20 VPWR.n17 0.119
R44 VPWR.n22 VPWR.n20 0.119
R45 VPWR.n24 VPWR.n22 0.119
R46 VPB.t9 VPB.t3 583.021
R47 VPB.t6 VPB.t1 556.386
R48 VPB.t0 VPB.t5 358.099
R49 VPB.t4 VPB.t0 284.112
R50 VPB.t11 VPB.t7 269.314
R51 VPB.t7 VPB.t10 260.436
R52 VPB.t3 VPB.t8 257.476
R53 VPB.t8 VPB.t11 248.598
R54 VPB.t1 VPB.t4 248.598
R55 VPB.t2 VPB.t6 248.598
R56 VPB.t5 VPB.t9 213.084
R57 VPB VPB.t2 192.367
R58 a_724_21.t0 a_724_21.n7 466.769
R59 a_724_21.n6 a_724_21.t3 368.328
R60 a_724_21.n0 a_724_21.t7 212.079
R61 a_724_21.n1 a_724_21.t2 212.079
R62 a_724_21.n2 a_724_21.t11 212.079
R63 a_724_21.n3 a_724_21.t5 212.079
R64 a_724_21.n6 a_724_21.t6 149.821
R65 a_724_21.n4 a_724_21.t1 145.846
R66 a_724_21.n0 a_724_21.t9 139.779
R67 a_724_21.n1 a_724_21.t4 139.779
R68 a_724_21.n2 a_724_21.t8 139.779
R69 a_724_21.n3 a_724_21.t10 139.779
R70 a_724_21.n4 a_724_21.n3 100.686
R71 a_724_21.n7 a_724_21.n6 97.139
R72 a_724_21.n2 a_724_21.n1 66.457
R73 a_724_21.n1 a_724_21.n0 64.266
R74 a_724_21.n3 a_724_21.n2 61.345
R75 a_724_21.n5 a_724_21.n4 16.78
R76 a_724_21.n7 a_724_21.n5 0.969
R77 Q.n1 Q.n0 144.894
R78 Q.n5 Q.n4 144.822
R79 Q.n3 Q.n2 92.5
R80 Q.n7 Q.n6 92.5
R81 Q.n4 Q.t2 30.535
R82 Q.n6 Q.t6 28.615
R83 Q.n0 Q.t1 26.595
R84 Q.n0 Q.t3 26.595
R85 Q.n4 Q.t4 26.595
R86 Q.n9 Q.n3 26.233
R87 Q Q.n9 25.824
R88 Q.n2 Q.t7 24.923
R89 Q.n2 Q.t5 24.923
R90 Q.n6 Q.t0 24.923
R91 Q.n8 Q 21.807
R92 Q.n8 Q 14.351
R93 Q.n8 Q 10.903
R94 Q Q.n7 10.192
R95 Q.n9 Q 10.084
R96 Q Q.n5 9
R97 Q Q.n1 8.538
R98 Q.n3 Q 6.961
R99 Q.n5 Q 6.807
R100 Q.n1 Q 6.452
R101 Q.n7 Q 5.925
R102 Q Q.n8 3.49
R103 a_27_47.t0 a_27_47.n3 269.575
R104 a_27_47.n1 a_27_47.t5 263.171
R105 a_27_47.n0 a_27_47.t4 240.108
R106 a_27_47.n0 a_27_47.t2 239.726
R107 a_27_47.n1 a_27_47.t3 227.825
R108 a_27_47.n2 a_27_47.t1 202.368
R109 a_27_47.n2 a_27_47.n1 76
R110 a_27_47.n3 a_27_47.n2 18.97
R111 a_27_47.n3 a_27_47.n0 11.268
R112 a_465_47.n0 a_465_47.t0 88.333
R113 a_465_47.n0 a_465_47.t1 26.393
R114 a_465_47.n1 a_465_47.n0 14.4
R115 a_561_413.n3 a_561_413.n2 422.17
R116 a_561_413.n0 a_561_413.t4 212.079
R117 a_561_413.n2 a_561_413.n1 190.005
R118 a_561_413.n2 a_561_413.n0 179.229
R119 a_561_413.n0 a_561_413.t5 139.779
R120 a_561_413.t0 a_561_413.n3 121.952
R121 a_561_413.n3 a_561_413.t1 91.464
R122 a_561_413.n1 a_561_413.t3 46.666
R123 a_561_413.n1 a_561_413.t2 46.666
R124 VNB VNB.t1 6470.59
R125 VNB.t2 VNB.t0 6082.35
R126 VNB.t10 VNB.t11 5613.06
R127 VNB.t5 VNB.t3 3494.12
R128 VNB.t4 VNB.t10 3073.53
R129 VNB.t3 VNB.t4 2782.35
R130 VNB.t0 VNB.t5 2717.65
R131 VNB.t1 VNB.t2 2717.65
R132 VNB.t8 VNB.t9 2200
R133 VNB.t9 VNB.t7 2127.47
R134 VNB.t11 VNB.t6 2103.3
R135 VNB.t6 VNB.t8 2030.77
R136 VGND.n2 VGND.t5 148.607
R137 VGND.n10 VGND.t8 148.331
R138 VGND.n1 VGND.n0 120.66
R139 VGND.n6 VGND.n5 117.201
R140 VGND.n26 VGND.n25 107.239
R141 VGND.n19 VGND.n18 106.463
R142 VGND.n18 VGND.t3 38.571
R143 VGND.n18 VGND.t0 38.571
R144 VGND.n25 VGND.t2 38.571
R145 VGND.n25 VGND.t1 38.571
R146 VGND.n0 VGND.t6 31.384
R147 VGND.n5 VGND.t9 27.692
R148 VGND.n0 VGND.t7 24.923
R149 VGND.n5 VGND.t4 24.923
R150 VGND.n4 VGND.n3 4.65
R151 VGND.n7 VGND.n6 4.65
R152 VGND.n9 VGND.n8 4.65
R153 VGND.n11 VGND.n10 4.65
R154 VGND.n13 VGND.n12 4.65
R155 VGND.n15 VGND.n14 4.65
R156 VGND.n17 VGND.n16 4.65
R157 VGND.n20 VGND.n19 4.65
R158 VGND.n22 VGND.n21 4.65
R159 VGND.n24 VGND.n23 4.65
R160 VGND.n27 VGND.n26 3.932
R161 VGND.n2 VGND.n1 3.778
R162 VGND.n4 VGND.n2 0.24
R163 VGND.n27 VGND.n24 0.137
R164 VGND VGND.n27 0.123
R165 VGND.n7 VGND.n4 0.119
R166 VGND.n9 VGND.n7 0.119
R167 VGND.n11 VGND.n9 0.119
R168 VGND.n13 VGND.n11 0.119
R169 VGND.n15 VGND.n13 0.119
R170 VGND.n17 VGND.n15 0.119
R171 VGND.n20 VGND.n17 0.119
R172 VGND.n22 VGND.n20 0.119
R173 VGND.n24 VGND.n22 0.119
R174 a_193_47.n0 a_193_47.t3 464.325
R175 a_193_47.n0 a_193_47.t2 242.606
R176 a_193_47.n1 a_193_47.t0 230.004
R177 a_193_47.t1 a_193_47.n1 121.759
R178 a_193_47.n1 a_193_47.n0 99.063
R179 a_465_369.t0 a_465_369.t1 134.63
R180 a_659_47.t0 a_659_47.t1 93.059
R181 GATE_N.n0 GATE_N.t0 269.919
R182 GATE_N.n0 GATE_N.t1 234.573
R183 GATE_N.n1 GATE_N.n0 76
R184 GATE_N GATE_N.n1 10.971
R185 GATE_N.n1 GATE_N 6.791
R186 a_682_413.t0 a_682_413.t1 98.5
C0 VGND Q 0.38fF
C1 VPWR Q 0.82fF
C2 VPWR VGND 0.12fF
C3 VPWR VPB 0.15fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__dlxtp_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__dlxtp_1 D GATE Q VGND VPWR VNB VPB
X0 a_560_47.t0 a_193_47.t2 a_465_47.t1 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X1 VPWR.t1 D.t0 a_299_47.t0 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X2 VGND.t3 a_713_21.t2 a_659_47.t0 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X3 Q.t0 a_713_21.t3 VGND.t2 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 a_465_47.t0 a_299_47.t2 VGND.t4 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 VPWR.t5 GATE.t0 a_27_47.t1 VPB.t6 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X6 a_659_47.t1 a_27_47.t2 a_560_47.t2 VNB.t6 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X7 VGND.t0 a_560_47.t4 a_713_21.t1 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 VPWR.t2 a_713_21.t4 a_644_413.t0 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9 a_193_47.t0 a_27_47.t3 VGND.t6 VNB.t7 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10 VPWR.t0 a_560_47.t5 a_713_21.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 a_193_47.t1 a_27_47.t4 VPWR.t6 VPB.t7 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X12 Q.t1 a_713_21.t5 VPWR.t3 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13 VGND.t1 D.t1 a_299_47.t1 VNB.t8 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14 a_644_413.t1 a_193_47.t3 a_560_47.t1 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15 a_465_369.t1 a_299_47.t3 VPWR.t4 VPB.t5 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X16 a_560_47.t3 a_27_47.t5 a_465_369.t0 VPB.t8 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17 VGND.t5 GATE.t1 a_27_47.t0 VNB.t5 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
R0 a_193_47.n0 a_193_47.t2 254.216
R1 a_193_47.n1 a_193_47.t0 230.004
R2 a_193_47.n0 a_193_47.t3 146.481
R3 a_193_47.t1 a_193_47.n1 121.759
R4 a_193_47.n1 a_193_47.n0 6.199
R5 a_465_47.n0 a_465_47.t1 66.666
R6 a_465_47.n0 a_465_47.t0 26.393
R7 a_465_47.n1 a_465_47.n0 14.4
R8 a_560_47.n3 a_560_47.n2 429.37
R9 a_560_47.n0 a_560_47.t5 212.079
R10 a_560_47.n2 a_560_47.n1 187.369
R11 a_560_47.n2 a_560_47.n0 170.488
R12 a_560_47.n0 a_560_47.t4 139.779
R13 a_560_47.n1 a_560_47.t0 68.333
R14 a_560_47.t1 a_560_47.n3 63.321
R15 a_560_47.n3 a_560_47.t3 63.321
R16 a_560_47.n1 a_560_47.t2 46.666
R17 VNB.t7 VNB.t8 6082.35
R18 VNB.t2 VNB.t0 5690.29
R19 VNB VNB.t5 4270.59
R20 VNB.t4 VNB.t6 3512.9
R21 VNB.t1 VNB.t4 3011.81
R22 VNB.t6 VNB.t2 2980.65
R23 VNB.t8 VNB.t1 2717.65
R24 VNB.t5 VNB.t7 2717.65
R25 VNB.t0 VNB.t3 2103.3
R26 D.n0 D.t0 327.642
R27 D.n0 D.t1 157.336
R28 D D.n0 78.594
R29 a_299_47.n0 a_299_47.t3 373.281
R30 a_299_47.t0 a_299_47.n1 292.715
R31 a_299_47.n1 a_299_47.t1 182.645
R32 a_299_47.n0 a_299_47.t2 132.281
R33 a_299_47.n1 a_299_47.n0 80.46
R34 VPWR.n0 VPWR.t2 385.734
R35 VPWR.n17 VPWR.n16 311.893
R36 VPWR.n2 VPWR.n1 182.806
R37 VPWR.n10 VPWR.n9 165.066
R38 VPWR.n9 VPWR.t4 41.554
R39 VPWR.n9 VPWR.t1 41.554
R40 VPWR.n16 VPWR.t6 41.554
R41 VPWR.n16 VPWR.t5 41.554
R42 VPWR.n1 VPWR.t0 29.55
R43 VPWR.n1 VPWR.t3 26.595
R44 VPWR.n2 VPWR.n0 7.841
R45 VPWR.n4 VPWR.n3 4.65
R46 VPWR.n6 VPWR.n5 4.65
R47 VPWR.n8 VPWR.n7 4.65
R48 VPWR.n11 VPWR.n10 4.65
R49 VPWR.n13 VPWR.n12 4.65
R50 VPWR.n15 VPWR.n14 4.65
R51 VPWR.n18 VPWR.n17 3.932
R52 VPWR.n4 VPWR.n2 0.196
R53 VPWR.n18 VPWR.n15 0.137
R54 VPWR VPWR.n18 0.123
R55 VPWR.n6 VPWR.n4 0.119
R56 VPWR.n8 VPWR.n6 0.119
R57 VPWR.n11 VPWR.n8 0.119
R58 VPWR.n13 VPWR.n11 0.119
R59 VPWR.n15 VPWR.n13 0.119
R60 VPB.t2 VPB.t0 562.305
R61 VPB.t7 VPB.t1 556.386
R62 VPB.t4 VPB.t2 292.99
R63 VPB.t5 VPB.t8 281.152
R64 VPB.t0 VPB.t3 257.476
R65 VPB.t8 VPB.t4 248.598
R66 VPB.t1 VPB.t5 248.598
R67 VPB.t6 VPB.t7 248.598
R68 VPB VPB.t6 142.056
R69 a_713_21.t0 a_713_21.n4 466.769
R70 a_713_21.n3 a_713_21.t2 375.959
R71 a_713_21.n0 a_713_21.t5 241.534
R72 a_713_21.n0 a_713_21.t3 169.234
R73 a_713_21.n3 a_713_21.t4 147.812
R74 a_713_21.n1 a_713_21.t1 145.846
R75 a_713_21.n1 a_713_21.n0 98.496
R76 a_713_21.n4 a_713_21.n3 93.648
R77 a_713_21.n2 a_713_21.n1 16.78
R78 a_713_21.n4 a_713_21.n2 0.969
R79 a_659_47.t0 a_659_47.t1 90
R80 VGND.n1 VGND.t3 154.76
R81 VGND.n2 VGND.n0 130.535
R82 VGND.n17 VGND.n16 107.239
R83 VGND.n10 VGND.n9 106.463
R84 VGND.n9 VGND.t4 38.571
R85 VGND.n9 VGND.t1 38.571
R86 VGND.n16 VGND.t6 38.571
R87 VGND.n16 VGND.t5 38.571
R88 VGND.n0 VGND.t0 27.692
R89 VGND.n0 VGND.t2 24.923
R90 VGND.n4 VGND.n3 4.65
R91 VGND.n6 VGND.n5 4.65
R92 VGND.n8 VGND.n7 4.65
R93 VGND.n11 VGND.n10 4.65
R94 VGND.n13 VGND.n12 4.65
R95 VGND.n15 VGND.n14 4.65
R96 VGND.n2 VGND.n1 3.949
R97 VGND.n18 VGND.n17 3.932
R98 VGND.n4 VGND.n2 0.212
R99 VGND.n18 VGND.n15 0.137
R100 VGND VGND.n18 0.123
R101 VGND.n6 VGND.n4 0.119
R102 VGND.n8 VGND.n6 0.119
R103 VGND.n11 VGND.n8 0.119
R104 VGND.n13 VGND.n11 0.119
R105 VGND.n15 VGND.n13 0.119
R106 Q.n0 Q.t1 176.414
R107 Q.n1 Q.t0 122.038
R108 Q Q.n1 82.221
R109 Q Q.n0 8.538
R110 Q.n1 Q 6.961
R111 Q.n0 Q 6.452
R112 GATE.n0 GATE.t0 270.454
R113 GATE.n0 GATE.t1 235.108
R114 GATE.n1 GATE.n0 76
R115 GATE GATE.n1 11.2
R116 GATE.n1 GATE 6.933
R117 a_27_47.n0 a_27_47.t2 424.811
R118 a_27_47.t1 a_27_47.n3 269.575
R119 a_27_47.n1 a_27_47.t4 263.171
R120 a_27_47.n1 a_27_47.t3 227.825
R121 a_27_47.n0 a_27_47.t5 218.88
R122 a_27_47.n2 a_27_47.t0 202.368
R123 a_27_47.n2 a_27_47.n1 76
R124 a_27_47.n3 a_27_47.n2 18.97
R125 a_27_47.n3 a_27_47.n0 16.829
R126 a_644_413.t0 a_644_413.t1 161.821
R127 a_465_369.t1 a_465_369.t0 132.285
C0 VPWR Q 0.13fF
C1 VPB VPWR 0.12fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__dlygate4sd1_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__dlygate4sd1_1 A X VPWR VGND VNB VPB
X0 X.t0 a_299_93.t2 VGND.t0 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 VPWR.t2 a_193_47.t2 a_299_93.t0 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 VPWR.t1 A.t0 a_27_47.t1 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3 a_193_47.t0 a_27_47.t2 VGND.t3 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 a_193_47.t1 a_27_47.t3 VPWR.t3 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 VGND.t2 a_193_47.t3 a_299_93.t1 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 X.t1 a_299_93.t3 VPWR.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 VGND.t1 A.t1 a_27_47.t0 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
R0 a_299_93.t0 a_299_93.n1 423.981
R1 a_299_93.n0 a_299_93.t3 238.589
R2 a_299_93.n1 a_299_93.t1 178.739
R3 a_299_93.n0 a_299_93.t2 166.289
R4 a_299_93.n1 a_299_93.n0 76
R5 VGND.n2 VGND.n0 118.662
R6 VGND.n2 VGND.n1 113.607
R7 VGND.n1 VGND.t2 58.571
R8 VGND.n0 VGND.t3 38.571
R9 VGND.n0 VGND.t1 38.571
R10 VGND.n1 VGND.t0 24
R11 VGND VGND.n2 0.149
R12 X.n1 X.t1 170.811
R13 X.n0 X.t0 117.423
R14 X X.n0 78.626
R15 X.n1 X 10.286
R16 X X.n1 6.19
R17 X.n0 X 3.751
R18 VNB VNB.t1 6502.94
R19 VNB.t3 VNB.t2 5321.88
R20 VNB.t1 VNB.t3 2717.65
R21 VNB.t2 VNB.t0 2345.05
R22 a_193_47.n1 a_193_47.t1 429.07
R23 a_193_47.n0 a_193_47.t2 206.689
R24 a_193_47.t0 a_193_47.n1 176.461
R25 a_193_47.n0 a_193_47.t3 119.929
R26 a_193_47.n1 a_193_47.n0 101.28
R27 VPWR.n2 VPWR.n0 321.819
R28 VPWR.n2 VPWR.n1 318.662
R29 VPWR.n0 VPWR.t2 89.119
R30 VPWR.n1 VPWR.t3 63.321
R31 VPWR.n1 VPWR.t1 63.321
R32 VPWR.n0 VPWR.t0 37.313
R33 VPWR VPWR.n2 0.149
R34 VPB.t3 VPB.t2 562.305
R35 VPB.t2 VPB.t0 281.152
R36 VPB.t1 VPB.t3 248.598
R37 VPB VPB.t1 195.327
R38 A.n0 A.t0 326.76
R39 A.n0 A.t1 198.227
R40 A.n1 A.n0 76
R41 A.n1 A 7.761
R42 A A.n1 1.497
R43 a_27_47.n1 a_27_47.t1 437.423
R44 a_27_47.n0 a_27_47.t3 334.721
R45 a_27_47.n0 a_27_47.t2 206.188
R46 a_27_47.t0 a_27_47.n1 193.035
R47 a_27_47.n1 a_27_47.n0 76
C0 VPWR X 0.14fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__dlygate4sd2_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__dlygate4sd2_1 VGND VPWR X A VNB VPB
X0 VPWR.t0 A.t0 a_49_47.t1 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1 VPWR.t3 a_221_47.t2 a_327_47.t1 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=180000u
X2 X.t0 a_327_47.t2 VGND.t2 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 VGND.t1 A.t1 a_49_47.t0 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 X.t1 a_327_47.t3 VPWR.t1 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 a_221_47.t0 a_49_47.t2 VGND.t3 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=180000u
X6 a_221_47.t1 a_49_47.t3 VPWR.t2 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=180000u
X7 VGND.t0 a_221_47.t3 a_327_47.t0 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=180000u
R0 A.n0 A.t0 322.187
R1 A.n0 A.t1 193.654
R2 A.n1 A.n0 76
R3 A.n1 A 6.755
R4 A A.n1 1.303
R5 a_49_47.n1 a_49_47.t1 422.265
R6 a_49_47.n0 a_49_47.t3 283.843
R7 a_49_47.t0 a_49_47.n1 181.595
R8 a_49_47.n0 a_49_47.t2 176.732
R9 a_49_47.n1 a_49_47.n0 76
R10 VPWR.n2 VPWR.n0 313.931
R11 VPWR.n2 VPWR.n1 311.215
R12 VPWR.n1 VPWR.t3 75.047
R13 VPWR.n0 VPWR.t2 63.321
R14 VPWR.n0 VPWR.t0 63.321
R15 VPWR.n1 VPWR.t1 43.386
R16 VPWR VPWR.n2 0.159
R17 VPB.t2 VPB.t3 574.143
R18 VPB.t3 VPB.t1 290.031
R19 VPB.t0 VPB.t2 257.476
R20 VPB VPB.t0 257.476
R21 a_221_47.n1 a_221_47.t1 410.309
R22 a_221_47.n0 a_221_47.t2 272.061
R23 a_221_47.t0 a_221_47.n1 176.015
R24 a_221_47.n0 a_221_47.t3 164.95
R25 a_221_47.n1 a_221_47.n0 76
R26 a_327_47.n1 a_327_47.t1 432.419
R27 a_327_47.n0 a_327_47.t3 241.534
R28 a_327_47.t0 a_327_47.n1 189.221
R29 a_327_47.n0 a_327_47.t2 169.234
R30 a_327_47.n1 a_327_47.n0 76
R31 VGND.n2 VGND.n0 113.931
R32 VGND.n2 VGND.n1 111.215
R33 VGND.n1 VGND.t0 45.714
R34 VGND.n0 VGND.t3 38.571
R35 VGND.n0 VGND.t1 38.571
R36 VGND.n1 VGND.t2 34.505
R37 VGND VGND.n2 0.159
R38 X.n0 X.t1 171.895
R39 X.n2 X.t0 117.423
R40 X X.n3 7.791
R41 X.n1 X 6.569
R42 X X.n2 5.776
R43 X X.n0 4.776
R44 X.n0 X 2.87
R45 X.n2 X 1.925
R46 X.n3 X 1.669
R47 X X.n1 1.391
R48 X.n3 X 1.359
R49 X.n1 X 1.132
R50 VNB VNB.t1 7182.35
R51 VNB.t3 VNB.t0 6276.47
R52 VNB.t1 VNB.t3 2814.71
R53 VNB.t0 VNB.t2 2296.85
C0 X VGND 0.13fF
C1 VPWR X 0.14fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__dlygate4sd3_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__dlygate4sd3_1 A X VGND VPWR VNB VPB
X0 VPWR.t3 A.t0 a_49_47.t1 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1 VGND.t1 a_285_47.t2 a_391_47.t0 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=500000u
X2 X.t1 a_391_47.t2 VPWR.t2 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 VGND.t3 A.t1 a_49_47.t0 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 VPWR.t1 a_285_47.t3 a_391_47.t1 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=500000u
X5 a_285_47.t0 a_49_47.t2 VGND.t0 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=500000u
X6 a_285_47.t1 a_49_47.t3 VPWR.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=500000u
X7 X.t0 a_391_47.t3 VGND.t2 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
R0 A.n0 A.t0 331.776
R1 A.n0 A.t1 203.243
R2 A.n1 A.n0 76
R3 A A.n1 7.885
R4 A.n1 A 2.628
R5 a_49_47.n1 a_49_47.t1 440.935
R6 a_49_47.t0 a_49_47.n1 200.672
R7 a_49_47.n0 a_49_47.t3 107.486
R8 a_49_47.n1 a_49_47.n0 76
R9 a_49_47.n0 a_49_47.t2 68.926
R10 VPWR.n2 VPWR.n0 313.937
R11 VPWR.n2 VPWR.n1 311.362
R12 VPWR.n1 VPWR.t1 75.047
R13 VPWR.n0 VPWR.t0 63.321
R14 VPWR.n0 VPWR.t3 63.321
R15 VPWR.n1 VPWR.t2 43.386
R16 VPWR VPWR.n2 0.152
R17 VPB.t0 VPB.t1 763.551
R18 VPB.t1 VPB.t2 384.735
R19 VPB.t3 VPB.t0 352.18
R20 VPB VPB.t3 257.476
R21 a_285_47.n1 a_285_47.t1 380.179
R22 a_285_47.t0 a_285_47.n1 149.738
R23 a_285_47.n0 a_285_47.t3 107.486
R24 a_285_47.n1 a_285_47.n0 95.718
R25 a_285_47.n0 a_285_47.t2 68.926
R26 a_391_47.n1 a_391_47.t1 414.108
R27 a_391_47.n0 a_391_47.t2 241.534
R28 a_391_47.t0 a_391_47.n1 184.309
R29 a_391_47.n0 a_391_47.t3 169.234
R30 a_391_47.n1 a_391_47.n0 76.775
R31 VGND.n2 VGND.n1 113.937
R32 VGND.n2 VGND.n0 111.359
R33 VGND.n0 VGND.t1 45.714
R34 VGND.n1 VGND.t0 38.571
R35 VGND.n1 VGND.t3 38.571
R36 VGND.n0 VGND.t2 34.505
R37 VGND VGND.n2 0.152
R38 VNB.t0 VNB.t1 8347.06
R39 VNB VNB.t3 7182.35
R40 VNB.t3 VNB.t0 3850
R41 VNB.t1 VNB.t2 2739.62
R42 X X.t1 465.805
R43 X.n0 X.t0 117.423
R44 X X.n1 12.8
R45 X.n2 X 9.641
R46 X X.n0 8.477
R47 X.n0 X 2.825
R48 X.n1 X 2.742
R49 X.n2 X 2.285
R50 X.n1 X 1.994
R51 X X.n2 1.662
C0 X VGND 0.10fF
C1 VPWR X 0.11fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__dlymetal6s2s_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__dlymetal6s2s_1 VPWR VGND A X VNB VPB
X0 a_558_47.t1 a_381_47.t2 VPWR.t4 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 VGND.t0 X.t2 a_381_47.t0 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 a_841_47.t0 a_664_47.t2 VPWR.t5 VPB.t5 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 VPWR.t3 A.t0 a_62_47.t0 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 VGND.t3 A.t1 a_62_47.t1 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 a_558_47.t0 a_381_47.t3 VGND.t4 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 X.t0 a_62_47.t2 VPWR.t1 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 VPWR.t0 X.t3 a_381_47.t1 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 a_841_47.t1 a_664_47.t3 VGND.t5 VNB.t5 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 X.t1 a_62_47.t3 VGND.t2 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 VPWR.t2 a_558_47.t2 a_664_47.t0 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11 VGND.t1 a_558_47.t3 a_664_47.t1 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
R0 a_381_47.n1 a_381_47.t1 413.394
R1 a_381_47.n0 a_381_47.t2 241.534
R2 a_381_47.t0 a_381_47.n1 176.924
R3 a_381_47.n0 a_381_47.t3 169.234
R4 a_381_47.n1 a_381_47.n0 76
R5 VPWR.n3 VPWR.n2 296.548
R6 VPWR.n11 VPWR.n10 292.5
R7 VPWR.n1 VPWR.n0 292.5
R8 VPWR.n10 VPWR.t3 77.392
R9 VPWR.n0 VPWR.t0 77.392
R10 VPWR.n2 VPWR.t2 77.392
R11 VPWR.n10 VPWR.t1 41.041
R12 VPWR.n0 VPWR.t4 41.041
R13 VPWR.n2 VPWR.t5 41.041
R14 VPWR.n12 VPWR.n11 8.341
R15 VPWR.n3 VPWR.n1 5.099
R16 VPWR.n9 VPWR.n8 4.65
R17 VPWR.n5 VPWR.n4 4.65
R18 VPWR.n7 VPWR.n6 4.65
R19 VPWR.n5 VPWR.n3 0.146
R20 VPWR VPWR.n12 0.135
R21 VPWR.n12 VPWR.n9 0.132
R22 VPWR.n7 VPWR.n5 0.119
R23 VPWR.n9 VPWR.n7 0.119
R24 a_558_47.n0 a_558_47.t2 323.548
R25 a_558_47.t1 a_558_47.n1 218.553
R26 a_558_47.n0 a_558_47.t3 195.015
R27 a_558_47.n1 a_558_47.t0 153.586
R28 a_558_47.n1 a_558_47.n0 76
R29 VPB.t2 VPB.t0 662.928
R30 VPB.t4 VPB.t1 556.386
R31 VPB VPB.t3 310.747
R32 VPB.t1 VPB.t5 281.152
R33 VPB.t0 VPB.t4 281.152
R34 VPB.t3 VPB.t2 281.152
R35 X.n1 X.t3 323.548
R36 X.n1 X.t2 195.015
R37 X.n0 X.t0 172.919
R38 X.n4 X.t1 117.423
R39 X X.n1 77.408
R40 X.n2 X 16.711
R41 X.n2 X 16
R42 X X.n4 9.788
R43 X X.n0 7.712
R44 X.n3 X 6.345
R45 X X.n2 6.016
R46 X.n2 X 5.76
R47 X.n0 X 2.486
R48 X.n3 X 2.194
R49 X X.n3 1.807
R50 X.n4 X 0.451
R51 VGND.n3 VGND.n2 96.645
R52 VGND.n1 VGND.n0 92.5
R53 VGND.n11 VGND.n10 92.5
R54 VGND.n10 VGND.t3 45.714
R55 VGND.n0 VGND.t0 45.714
R56 VGND.n2 VGND.t1 45.714
R57 VGND.n10 VGND.t2 34.505
R58 VGND.n0 VGND.t4 34.505
R59 VGND.n2 VGND.t5 34.505
R60 VGND.n12 VGND.n11 8.413
R61 VGND.n3 VGND.n1 5.261
R62 VGND.n5 VGND.n4 4.65
R63 VGND.n7 VGND.n6 4.65
R64 VGND.n9 VGND.n8 4.65
R65 VGND.n5 VGND.n3 0.146
R66 VGND VGND.n12 0.135
R67 VGND.n12 VGND.n9 0.132
R68 VGND.n7 VGND.n5 0.119
R69 VGND.n9 VGND.n7 0.119
R70 VNB VNB.t3 7852.94
R71 VNB.t2 VNB.t0 5415.38
R72 VNB.t4 VNB.t1 4545.05
R73 VNB.t1 VNB.t5 2296.7
R74 VNB.t0 VNB.t4 2296.7
R75 VNB.t3 VNB.t2 2255.35
R76 a_664_47.t0 a_664_47.n1 414.617
R77 a_664_47.n0 a_664_47.t2 241.534
R78 a_664_47.n1 a_664_47.t1 176.924
R79 a_664_47.n0 a_664_47.t3 169.234
R80 a_664_47.n1 a_664_47.n0 76
R81 a_841_47.t0 a_841_47.t1 382.539
R82 A.n0 A.t0 323.548
R83 A.n0 A.t1 195.015
R84 A.n1 A.n0 76
R85 A.n1 A 7.521
R86 A A.n1 1.451
R87 a_62_47.t0 a_62_47.n1 412.177
R88 a_62_47.n0 a_62_47.t2 241.534
R89 a_62_47.n1 a_62_47.t1 172.362
R90 a_62_47.n0 a_62_47.t3 169.234
R91 a_62_47.n1 a_62_47.n0 76
C0 VPWR VGND 0.10fF
C1 X VGND 0.12fF
C2 X VPWR 0.12fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__dlymetal6s4s_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__dlymetal6s4s_1 VPWR VGND A X VNB VPB
X0 X.t0 a_345_47.t2 VGND.t4 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 VPWR.t0 a_239_47.t2 a_345_47.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 a_841_47.t1 a_664_47.t2 VPWR.t2 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 VGND.t3 a_239_47.t3 a_345_47.t1 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 VPWR.t3 A.t0 a_62_47.t1 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 VGND.t2 A.t1 a_62_47.t0 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 X.t1 a_345_47.t3 VPWR.t4 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 a_239_47.t0 a_62_47.t2 VPWR.t5 VPB.t5 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 a_841_47.t0 a_664_47.t3 VGND.t1 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 a_239_47.t1 a_62_47.t3 VGND.t5 VNB.t5 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 VPWR.t1 X.t2 a_664_47.t1 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11 VGND.t0 X.t3 a_664_47.t0 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
R0 a_345_47.t0 a_345_47.n1 414.954
R1 a_345_47.n0 a_345_47.t3 241.534
R2 a_345_47.n1 a_345_47.t1 177.226
R3 a_345_47.n0 a_345_47.t2 169.234
R4 a_345_47.n1 a_345_47.n0 76
R5 VGND.n1 VGND.n0 96.65
R6 VGND.n3 VGND.n2 92.5
R7 VGND.n11 VGND.n10 92.5
R8 VGND.n10 VGND.t2 45.714
R9 VGND.n2 VGND.t3 45.714
R10 VGND.n0 VGND.t0 45.714
R11 VGND.n10 VGND.t5 34.505
R12 VGND.n2 VGND.t4 34.505
R13 VGND.n0 VGND.t1 34.505
R14 VGND.n12 VGND.n11 8.413
R15 VGND.n4 VGND.n3 6.901
R16 VGND.n5 VGND.n4 4.65
R17 VGND.n7 VGND.n6 4.65
R18 VGND.n9 VGND.n8 4.65
R19 VGND.n5 VGND.n1 0.141
R20 VGND VGND.n12 0.135
R21 VGND.n12 VGND.n9 0.132
R22 VGND.n7 VGND.n5 0.119
R23 VGND.n9 VGND.n7 0.119
R24 X.n1 X.t2 323.548
R25 X.n1 X.t3 195.015
R26 X.n0 X.t1 172.916
R27 X.n5 X.t0 117.423
R28 X X.n1 77.792
R29 X.n2 X 17.777
R30 X.n2 X 14.933
R31 X X.n5 9.348
R32 X X.n0 7.367
R33 X.n3 X.n2 5.888
R34 X.n4 X.n3 5.881
R35 X.n2 X 5.376
R36 X.n0 X 2.375
R37 X.n4 X 2.075
R38 X X.n4 1.725
R39 X.n3 X 0.512
R40 X.n5 X 0.431
R41 VNB VNB.t2 7852.94
R42 VNB.t4 VNB.t0 5415.38
R43 VNB.t5 VNB.t3 4545.05
R44 VNB.t0 VNB.t1 2296.7
R45 VNB.t3 VNB.t4 2296.7
R46 VNB.t2 VNB.t5 2255.35
R47 a_239_47.n0 a_239_47.t2 323.548
R48 a_239_47.t0 a_239_47.n1 215.719
R49 a_239_47.n0 a_239_47.t3 195.015
R50 a_239_47.n1 a_239_47.t1 150.081
R51 a_239_47.n1 a_239_47.n0 76
R52 VPWR.n3 VPWR.n2 296.553
R53 VPWR.n11 VPWR.n10 292.5
R54 VPWR.n1 VPWR.n0 292.5
R55 VPWR.n10 VPWR.t3 77.392
R56 VPWR.n0 VPWR.t0 77.392
R57 VPWR.n2 VPWR.t1 77.392
R58 VPWR.n10 VPWR.t5 41.041
R59 VPWR.n0 VPWR.t4 41.041
R60 VPWR.n2 VPWR.t2 41.041
R61 VPWR.n3 VPWR.n1 11.231
R62 VPWR.n12 VPWR.n11 8.341
R63 VPWR.n9 VPWR.n8 4.65
R64 VPWR.n5 VPWR.n4 4.65
R65 VPWR.n7 VPWR.n6 4.65
R66 VPWR.n5 VPWR.n3 0.141
R67 VPWR VPWR.n12 0.135
R68 VPWR.n12 VPWR.n9 0.132
R69 VPWR.n7 VPWR.n5 0.119
R70 VPWR.n9 VPWR.n7 0.119
R71 VPB.t4 VPB.t1 662.928
R72 VPB.t5 VPB.t0 556.386
R73 VPB VPB.t3 310.747
R74 VPB.t1 VPB.t2 281.152
R75 VPB.t0 VPB.t4 281.152
R76 VPB.t3 VPB.t5 281.152
R77 a_664_47.n1 a_664_47.t1 414.617
R78 a_664_47.n0 a_664_47.t2 241.534
R79 a_664_47.t0 a_664_47.n1 176.924
R80 a_664_47.n0 a_664_47.t3 169.234
R81 a_664_47.n1 a_664_47.n0 76
R82 a_841_47.t1 a_841_47.t0 382.539
R83 A.n0 A.t0 323.548
R84 A.n0 A.t1 195.015
R85 A.n1 A.n0 76
R86 A.n1 A 7.521
R87 A A.n1 1.451
R88 a_62_47.n1 a_62_47.t1 412.177
R89 a_62_47.n0 a_62_47.t2 241.534
R90 a_62_47.t0 a_62_47.n1 172.362
R91 a_62_47.n0 a_62_47.t3 169.234
R92 a_62_47.n1 a_62_47.n0 76
C0 VPWR VGND 0.10fF
C1 X VGND 0.13fF
C2 X VPWR 0.13fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__dlymetal6s6s_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__dlymetal6s6s_1 VPWR VGND A X VNB VPB
X0 X.t0 a_629_47.t2 VGND.t1 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 a_523_47.t0 a_346_47.t2 VGND.t4 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 VGND.t5 a_240_47.t2 a_346_47.t0 VNB.t5 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3 a_240_47.t1 a_63_47.t2 VGND.t2 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 VPWR.t0 a_240_47.t3 a_346_47.t1 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 VGND.t3 A.t0 a_63_47.t0 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 VPWR.t5 A.t1 a_63_47.t1 VPB.t5 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7 VPWR.t2 a_523_47.t2 a_629_47.t0 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 VGND.t0 a_523_47.t3 a_629_47.t1 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9 a_523_47.t1 a_346_47.t3 VPWR.t4 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 a_240_47.t0 a_63_47.t3 VPWR.t1 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 X.t1 a_629_47.t3 VPWR.t3 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
R0 a_629_47.t0 a_629_47.n1 413.683
R1 a_629_47.n0 a_629_47.t3 241.534
R2 a_629_47.n1 a_629_47.t1 176.088
R3 a_629_47.n0 a_629_47.t2 169.234
R4 a_629_47.n1 a_629_47.n0 76
R5 VGND.n3 VGND.n2 98.056
R6 VGND.n1 VGND.n0 92.5
R7 VGND.n11 VGND.n10 92.5
R8 VGND.n10 VGND.t3 45.714
R9 VGND.n0 VGND.t5 45.714
R10 VGND.n2 VGND.t0 45.714
R11 VGND.n10 VGND.t2 34.505
R12 VGND.n0 VGND.t4 34.505
R13 VGND.n2 VGND.t1 34.505
R14 VGND.n3 VGND.n1 11.133
R15 VGND.n12 VGND.n11 8.789
R16 VGND.n5 VGND.n4 4.65
R17 VGND.n7 VGND.n6 4.65
R18 VGND.n9 VGND.n8 4.65
R19 VGND.n5 VGND.n3 0.154
R20 VGND VGND.n12 0.134
R21 VGND.n12 VGND.n9 0.132
R22 VGND.n7 VGND.n5 0.119
R23 VGND.n9 VGND.n7 0.119
R24 X.n0 X.t1 172.918
R25 X.n3 X.t0 117.423
R26 X.n2 X 9.955
R27 X.n3 X 9.563
R28 X.n1 X 8.533
R29 X X.n0 7.536
R30 X.n0 X 2.429
R31 X.n2 X 2.133
R32 X X.n1 1.777
R33 X X.n2 1.765
R34 X.n1 X 1.471
R35 X X.n3 0.441
R36 VNB VNB.t3 7852.94
R37 VNB.t4 VNB.t0 4545.05
R38 VNB.t2 VNB.t5 4545.05
R39 VNB.t0 VNB.t1 2296.7
R40 VNB.t5 VNB.t4 2296.7
R41 VNB.t3 VNB.t2 2255.35
R42 a_346_47.n1 a_346_47.t1 414.954
R43 a_346_47.n0 a_346_47.t3 241.534
R44 a_346_47.t0 a_346_47.n1 177.226
R45 a_346_47.n0 a_346_47.t2 169.234
R46 a_346_47.n1 a_346_47.n0 76
R47 a_523_47.n0 a_523_47.t2 323.548
R48 a_523_47.t1 a_523_47.n1 217.816
R49 a_523_47.n0 a_523_47.t3 195.015
R50 a_523_47.n1 a_523_47.t0 152.818
R51 a_523_47.n1 a_523_47.n0 76
R52 a_240_47.n0 a_240_47.t3 323.548
R53 a_240_47.t0 a_240_47.n1 215.719
R54 a_240_47.n0 a_240_47.t2 195.015
R55 a_240_47.n1 a_240_47.t1 150.081
R56 a_240_47.n1 a_240_47.n0 76
R57 a_63_47.n1 a_63_47.t1 412.07
R58 a_63_47.n0 a_63_47.t3 241.534
R59 a_63_47.t0 a_63_47.n1 172.263
R60 a_63_47.n0 a_63_47.t2 169.234
R61 a_63_47.n1 a_63_47.n0 76
R62 VPWR.n5 VPWR.n4 297.934
R63 VPWR.n1 VPWR.n0 292.5
R64 VPWR.n3 VPWR.n2 292.5
R65 VPWR.n0 VPWR.t5 77.392
R66 VPWR.n2 VPWR.t0 77.392
R67 VPWR.n4 VPWR.t2 77.392
R68 VPWR.n0 VPWR.t1 41.041
R69 VPWR.n2 VPWR.t4 41.041
R70 VPWR.n4 VPWR.t3 41.041
R71 VPWR.n5 VPWR.n3 10.842
R72 VPWR.n12 VPWR.n1 8.717
R73 VPWR.n11 VPWR.n10 4.65
R74 VPWR.n7 VPWR.n6 4.65
R75 VPWR.n9 VPWR.n8 4.65
R76 VPWR.n7 VPWR.n5 0.154
R77 VPWR VPWR.n12 0.134
R78 VPWR.n12 VPWR.n11 0.132
R79 VPWR.n9 VPWR.n7 0.119
R80 VPWR.n11 VPWR.n9 0.119
R81 VPB.t4 VPB.t2 556.386
R82 VPB.t1 VPB.t0 556.386
R83 VPB VPB.t5 310.747
R84 VPB.t2 VPB.t3 281.152
R85 VPB.t0 VPB.t4 281.152
R86 VPB.t5 VPB.t1 281.152
R87 A.n0 A.t1 323.548
R88 A.n0 A.t0 195.015
R89 A.n1 A.n0 76
R90 A.n1 A 7.444
R91 A A.n1 1.436
C0 VPWR X 0.11fF
C1 VGND X 0.11fF
C2 VGND VPWR 0.10fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__ebufn_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__ebufn_1 Z TE_B A VPWR VGND VNB VPB
X0 Z.t0 a_27_47.t2 a_383_297.t1 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_193_369.t1 TE_B.t0 VGND.t0 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 a_383_297.t0 TE_B.t1 VPWR.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 VPWR.t2 A.t0 a_27_47.t0 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X4 a_531_47.t0 a_193_369.t2 VGND.t1 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 Z.t1 a_27_47.t3 a_531_47.t1 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 a_193_369.t0 TE_B.t2 VPWR.t1 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X7 VGND.t2 A.t1 a_27_47.t1 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
R0 a_27_47.t0 a_27_47.n1 430.039
R1 a_27_47.n1 a_27_47.n0 253.918
R2 a_27_47.n0 a_27_47.t2 241.534
R3 a_27_47.n0 a_27_47.t3 169.234
R4 a_27_47.n1 a_27_47.t1 155.58
R5 a_383_297.t0 a_383_297.t1 187.15
R6 Z.n3 Z.t0 183.68
R7 Z Z.n0 94.27
R8 Z.n1 Z.n0 92.5
R9 Z.n0 Z.t1 50.769
R10 Z Z.n2 10.541
R11 Z.n1 Z 7.489
R12 Z Z.n3 3.892
R13 Z.n2 Z 2.258
R14 Z.n3 Z 2.177
R15 Z Z.n1 1.77
R16 Z.n2 Z 1.634
R17 VPB.t0 VPB.t2 651.09
R18 VPB.t1 VPB.t0 562.305
R19 VPB.t3 VPB.t1 248.598
R20 VPB VPB.t3 189.408
R21 TE_B.n1 TE_B.t1 323.815
R22 TE_B.n0 TE_B.t2 282.334
R23 TE_B.n0 TE_B.t0 102.826
R24 TE_B.n2 TE_B.n1 76
R25 TE_B.n1 TE_B.n0 14.606
R26 TE_B.n2 TE_B 11.054
R27 TE_B TE_B.n2 2.133
R28 VGND.n1 VGND.t1 139.887
R29 VGND.n1 VGND.n0 111.017
R30 VGND.n0 VGND.t0 88.797
R31 VGND.n0 VGND.t2 38.572
R32 VGND VGND.n1 0.143
R33 a_193_369.t0 a_193_369.n0 383.799
R34 a_193_369.n0 a_193_369.t2 275.379
R35 a_193_369.n0 a_193_369.t1 245.496
R36 VNB.t1 VNB.t0 9477.63
R37 VNB VNB.t3 6438.23
R38 VNB.t3 VNB.t1 2359.04
R39 VNB.t0 VNB.t2 1740.66
R40 VPWR.n1 VPWR.t0 512.796
R41 VPWR.n1 VPWR.n0 309.801
R42 VPWR.n0 VPWR.t1 41.554
R43 VPWR.n0 VPWR.t2 41.554
R44 VPWR VPWR.n1 0.217
R45 A.n0 A.t0 289.316
R46 A.n0 A.t1 196.13
R47 A.n1 A.n0 76
R48 A.n1 A 13.511
R49 A A.n1 2.607
R50 a_531_47.t0 a_531_47.t1 38.769
C0 Z VGND 0.12fF
C1 VPWR Z 0.32fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__ebufn_2.ext - technology: sky130A

.subckt sky130_fd_sc_hd__ebufn_2 Z A TE_B VGND VPWR VNB VPB
X0 a_320_309.t3 a_27_47.t2 Z.t3 VPB.t5 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 Z.t2 a_27_47.t3 a_320_309.t2 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 VPWR.t3 A.t0 a_27_47.t0 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X3 VGND.t2 a_214_47.t2 a_392_47.t1 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 a_214_47.t0 TE_B.t0 VPWR.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X5 a_320_309.t0 TE_B.t1 VPWR.t1 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=940000u l=150000u
X6 a_392_47.t0 a_214_47.t3 VGND.t1 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 VPWR.t2 TE_B.t2 a_320_309.t1 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=940000u l=150000u
X8 Z.t1 a_27_47.t4 a_392_47.t3 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 a_214_47.t1 TE_B.t3 VGND.t0 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10 a_392_47.t2 a_27_47.t5 Z.t0 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 VGND.t3 A.t1 a_27_47.t1 VNB.t5 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
R0 a_27_47.t0 a_27_47.n3 388.191
R1 a_27_47.n0 a_27_47.t2 221.719
R2 a_27_47.n1 a_27_47.t3 221.719
R3 a_27_47.n3 a_27_47.t1 170.759
R4 a_27_47.n0 a_27_47.t5 149.419
R5 a_27_47.n1 a_27_47.t4 149.419
R6 a_27_47.n2 a_27_47.n0 38.188
R7 a_27_47.n2 a_27_47.n1 35.511
R8 a_27_47.n3 a_27_47.n2 17.289
R9 Z.n1 Z.n0 147.009
R10 Z Z.n2 114.849
R11 Z.n0 Z.t3 26.595
R12 Z.n0 Z.t2 26.595
R13 Z.n2 Z.t0 24.923
R14 Z.n2 Z.t1 24.923
R15 Z.n3 Z 21.945
R16 Z Z.n3 15
R17 Z.n3 Z.n1 4.405
R18 Z.n1 Z 2.535
R19 a_320_309.n0 a_320_309.t1 579.456
R20 a_320_309.n2 a_320_309.n1 298.277
R21 a_320_309.n1 a_320_309.t3 235.163
R22 a_320_309.n4 a_320_309.n3 45.058
R23 a_320_309.n3 a_320_309.t0 40.867
R24 a_320_309.n2 a_320_309.t2 28.529
R25 a_320_309.n4 a_320_309.n2 16.982
R26 a_320_309.n5 a_320_309.n4 8.82
R27 a_320_309.n1 a_320_309.n0 8.211
R28 VPB.t0 VPB.t2 556.386
R29 VPB.t1 VPB.t4 529.75
R30 VPB.t3 VPB.t0 310.747
R31 VPB.t4 VPB.t5 248.598
R32 VPB.t2 VPB.t1 248.598
R33 VPB VPB.t3 189.408
R34 A.n0 A.t0 295.166
R35 A.n0 A.t1 201.98
R36 A.n1 A.n0 76
R37 A.n1 A 17.434
R38 A A.n1 12.579
R39 VPWR.n2 VPWR.n0 310.177
R40 VPWR.n2 VPWR.n1 162.537
R41 VPWR.n1 VPWR.t3 58.484
R42 VPWR.n1 VPWR.t0 56.945
R43 VPWR.n0 VPWR.t1 28.292
R44 VPWR.n0 VPWR.t2 28.292
R45 VPWR VPWR.n2 0.156
R46 a_214_47.t0 a_214_47.n1 380.385
R47 a_214_47.n0 a_214_47.t2 237.786
R48 a_214_47.n1 a_214_47.t1 170.836
R49 a_214_47.n1 a_214_47.n0 148.785
R50 a_214_47.n0 a_214_47.t3 139.487
R51 a_392_47.t2 a_392_47.n1 234.972
R52 a_392_47.n1 a_392_47.t1 178.304
R53 a_392_47.n1 a_392_47.n0 92.5
R54 a_392_47.n0 a_392_47.t3 36
R55 a_392_47.n0 a_392_47.t0 35.076
R56 VGND.n2 VGND.n0 110.339
R57 VGND.n2 VGND.n1 109.666
R58 VGND.n1 VGND.t0 68.571
R59 VGND.n1 VGND.t3 38.571
R60 VGND.n0 VGND.t1 24.923
R61 VGND.n0 VGND.t2 24.923
R62 VGND VGND.n2 0.142
R63 VNB.t0 VNB.t2 7651.29
R64 VNB VNB.t5 6438.23
R65 VNB.t5 VNB.t0 3397.06
R66 VNB.t1 VNB.t4 2586.81
R67 VNB.t4 VNB.t3 2030.77
R68 VNB.t2 VNB.t1 2030.77
R69 TE_B.n0 TE_B.t1 284.379
R70 TE_B.n1 TE_B.t0 233.367
R71 TE_B.n1 TE_B.n0 210.473
R72 TE_B.n2 TE_B.t3 204.448
R73 TE_B.n0 TE_B.t2 175.126
R74 TE_B TE_B.n2 91.321
R75 TE_B.n2 TE_B.n1 31.463
C0 A TE_B 0.16fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__ebufn_4.ext - technology: sky130A

.subckt sky130_fd_sc_hd__ebufn_4 A Z TE_B VGND VPWR VNB VPB
X0 a_214_47.t1 TE_B.t0 VPWR.t1 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 Z.t3 a_27_47.t2 a_320_309.t7 VPB.t5 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 VGND.t5 a_214_47.t2 a_393_47.t7 VNB.t9 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 a_320_309.t3 TE_B.t1 VPWR.t0 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=940000u l=150000u
X4 VGND.t4 a_214_47.t3 a_393_47.t6 VNB.t8 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 VPWR.t4 TE_B.t2 a_320_309.t2 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=940000u l=150000u
X6 a_320_309.t1 TE_B.t3 VPWR.t3 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=940000u l=150000u
X7 a_393_47.t5 a_214_47.t4 VGND.t3 VNB.t7 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 Z.t7 a_27_47.t3 a_393_47.t3 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 VPWR.t2 TE_B.t4 a_320_309.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=940000u l=150000u
X10 a_393_47.t4 a_214_47.t5 VGND.t2 VNB.t6 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 Z.t6 a_27_47.t4 a_393_47.t2 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 a_393_47.t1 a_27_47.t5 Z.t5 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 a_214_47.t0 TE_B.t5 VGND.t0 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14 Z.t2 a_27_47.t6 a_320_309.t6 VPB.t6 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 a_320_309.t5 a_27_47.t7 Z.t1 VPB.t7 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16 a_393_47.t0 a_27_47.t8 Z.t4 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X17 a_320_309.t4 a_27_47.t9 Z.t0 VPB.t9 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X18 VPWR.t5 A.t0 a_27_47.t0 VPB.t8 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X19 VGND.t1 A.t1 a_27_47.t1 VNB.t5 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
R0 TE_B.n4 TE_B.t5 365.811
R1 TE_B.n0 TE_B.t1 310.086
R2 TE_B.n3 TE_B.t0 194.279
R3 TE_B.n3 TE_B.n2 186.602
R4 TE_B.n0 TE_B.t2 175.126
R5 TE_B.n1 TE_B.t3 175.126
R6 TE_B.n2 TE_B.t4 175.126
R7 TE_B.n1 TE_B.n0 134.96
R8 TE_B.n2 TE_B.n1 134.96
R9 TE_B TE_B.n4 91.321
R10 TE_B.n4 TE_B.n3 22.197
R11 VPWR.n3 VPWR.n2 309.964
R12 VPWR.n1 VPWR.n0 306.463
R13 VPWR.n9 VPWR.n8 159.929
R14 VPWR.n8 VPWR.t1 39.4
R15 VPWR.n8 VPWR.t5 34.475
R16 VPWR.n2 VPWR.t0 28.292
R17 VPWR.n2 VPWR.t4 28.292
R18 VPWR.n0 VPWR.t3 28.292
R19 VPWR.n0 VPWR.t2 28.292
R20 VPWR.n5 VPWR.n4 4.65
R21 VPWR.n7 VPWR.n6 4.65
R22 VPWR.n10 VPWR.n9 3.932
R23 VPWR.n3 VPWR.n1 3.659
R24 VPWR.n5 VPWR.n3 0.256
R25 VPWR.n10 VPWR.n7 0.137
R26 VPWR VPWR.n10 0.121
R27 VPWR.n7 VPWR.n5 0.119
R28 a_214_47.n0 a_214_47.t2 263.493
R29 a_214_47.t1 a_214_47.n3 222.867
R30 a_214_47.n3 a_214_47.n2 192.561
R31 a_214_47.n3 a_214_47.t0 157.56
R32 a_214_47.n2 a_214_47.t5 139.487
R33 a_214_47.n1 a_214_47.n0 134.96
R34 a_214_47.n0 a_214_47.t4 128.533
R35 a_214_47.n1 a_214_47.t3 128.533
R36 a_214_47.n2 a_214_47.n1 109.253
R37 VPB.t4 VPB.t0 556.386
R38 VPB.t3 VPB.t5 535.669
R39 VPB.t8 VPB.t4 310.747
R40 VPB.t6 VPB.t7 248.598
R41 VPB.t9 VPB.t6 248.598
R42 VPB.t5 VPB.t9 248.598
R43 VPB.t2 VPB.t3 248.598
R44 VPB.t1 VPB.t2 248.598
R45 VPB.t0 VPB.t1 248.598
R46 VPB VPB.t8 189.408
R47 a_27_47.n4 a_27_47.t7 221.719
R48 a_27_47.n6 a_27_47.t6 221.719
R49 a_27_47.n2 a_27_47.t9 221.719
R50 a_27_47.n0 a_27_47.t2 221.719
R51 a_27_47.t0 a_27_47.n11 217.834
R52 a_27_47.n11 a_27_47.t1 156.848
R53 a_27_47.n4 a_27_47.t5 149.419
R54 a_27_47.n6 a_27_47.t4 149.419
R55 a_27_47.n2 a_27_47.t8 149.419
R56 a_27_47.n0 a_27_47.t3 149.419
R57 a_27_47.n8 a_27_47.n5 93.408
R58 a_27_47.n8 a_27_47.n7 76
R59 a_27_47.n3 a_27_47.n2 37.331
R60 a_27_47.n3 a_27_47.n0 35.276
R61 a_27_47.n9 a_27_47.n8 17.408
R62 a_27_47.n5 a_27_47.n4 16.066
R63 a_27_47.n2 a_27_47.n1 12.496
R64 a_27_47.n10 a_27_47.n9 10.546
R65 a_27_47.n11 a_27_47.n10 9.947
R66 a_27_47.n10 a_27_47.n3 8.822
R67 a_27_47.n7 a_27_47.n6 1.785
R68 a_320_309.n1 a_320_309.t0 570.308
R69 a_320_309.n1 a_320_309.n0 307.182
R70 a_320_309.n3 a_320_309.t5 191.708
R71 a_320_309.n3 a_320_309.n2 146.25
R72 a_320_309.t3 a_320_309.n4 82.781
R73 a_320_309.n4 a_320_309.n1 53.766
R74 a_320_309.n4 a_320_309.t7 49.897
R75 a_320_309.n0 a_320_309.t2 28.292
R76 a_320_309.n0 a_320_309.t1 28.292
R77 a_320_309.n2 a_320_309.t6 26.595
R78 a_320_309.n2 a_320_309.t4 26.595
R79 a_320_309.n4 a_320_309.n3 23.915
R80 Z.n6 Z.n3 292.5
R81 Z.n5 Z.n4 292.5
R82 Z.n2 Z.n1 137.3
R83 Z.n2 Z.n0 92.5
R84 Z Z.n2 28.8
R85 Z.n4 Z.t0 26.595
R86 Z.n4 Z.t3 26.595
R87 Z.n3 Z.t1 26.595
R88 Z.n3 Z.t2 26.595
R89 Z.n0 Z.t5 24.923
R90 Z.n0 Z.t6 24.923
R91 Z.n1 Z.t4 24.923
R92 Z.n1 Z.t7 24.923
R93 Z Z.n5 21.028
R94 Z.n5 Z 21.028
R95 Z.n6 Z 17.371
R96 Z.n7 Z 14.545
R97 Z Z.n7 5.236
R98 Z.n7 Z 5.066
R99 Z Z.n6 3.657
R100 a_393_47.n3 a_393_47.t1 234.803
R101 a_393_47.n1 a_393_47.t7 174.657
R102 a_393_47.n1 a_393_47.n0 99.652
R103 a_393_47.n3 a_393_47.n2 92.5
R104 a_393_47.n5 a_393_47.n4 92.5
R105 a_393_47.n4 a_393_47.n3 60.131
R106 a_393_47.n4 a_393_47.n1 56.926
R107 a_393_47.t3 a_393_47.n5 36
R108 a_393_47.n5 a_393_47.t4 36
R109 a_393_47.n0 a_393_47.t6 24.923
R110 a_393_47.n0 a_393_47.t5 24.923
R111 a_393_47.n2 a_393_47.t2 24.923
R112 a_393_47.n2 a_393_47.t0 24.923
R113 VGND.n3 VGND.n0 109.876
R114 VGND.n2 VGND.n1 106.463
R115 VGND.n11 VGND.n10 92.5
R116 VGND.n10 VGND.t0 44.307
R117 VGND.n10 VGND.t1 24.923
R118 VGND.n0 VGND.t2 24.923
R119 VGND.n0 VGND.t4 24.923
R120 VGND.n1 VGND.t3 24.923
R121 VGND.n1 VGND.t5 24.923
R122 VGND.n13 VGND.n12 4.65
R123 VGND.n5 VGND.n4 4.65
R124 VGND.n7 VGND.n6 4.65
R125 VGND.n9 VGND.n8 4.65
R126 VGND.n3 VGND.n2 3.842
R127 VGND.n5 VGND.n3 0.257
R128 VGND.n12 VGND.n11 0.188
R129 VGND.n7 VGND.n5 0.119
R130 VGND.n9 VGND.n7 0.119
R131 VGND.n13 VGND.n9 0.119
R132 VGND.n14 VGND.n13 0.119
R133 VGND VGND.n14 0.02
R134 VNB.t0 VNB.t9 6309.89
R135 VNB VNB.t5 6053.91
R136 VNB.t6 VNB.t4 2610.99
R137 VNB.t5 VNB.t0 2538.46
R138 VNB.t3 VNB.t2 2030.77
R139 VNB.t1 VNB.t3 2030.77
R140 VNB.t4 VNB.t1 2030.77
R141 VNB.t8 VNB.t6 2030.77
R142 VNB.t7 VNB.t8 2030.77
R143 VNB.t9 VNB.t7 2030.77
R144 A.n0 A.t0 237.326
R145 A.n0 A.t1 165.026
R146 A.n1 A.n0 76
R147 A.n1 A 17.434
R148 A A.n1 12.579
C0 A TE_B 0.16fF
C1 VPWR VPB 0.11fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__ebufn_8.ext - technology: sky130A

.subckt sky130_fd_sc_hd__ebufn_8 A Z TE_B VGND VPWR VNB VPB
X0 VPWR.t7 TE_B.t0 a_407_309.t6 VPB.t13 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=940000u l=150000u
X1 a_455_47.t15 a_301_47.t2 VGND.t8 VNB.t16 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 Z.t15 a_116_47.t4 a_407_309.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 Z.t7 a_116_47.t5 a_455_47.t0 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 a_116_47.t0 A.t0 VPWR.t9 VPB.t17 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 a_407_309.t1 a_116_47.t6 Z.t14 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 VPWR.t6 TE_B.t1 a_407_309.t5 VPB.t12 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=940000u l=150000u
X7 a_407_309.t12 TE_B.t2 VPWR.t5 VPB.t11 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=940000u l=150000u
X8 VGND.t7 a_301_47.t3 a_455_47.t14 VNB.t15 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 VGND.t6 a_301_47.t4 a_455_47.t13 VNB.t14 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 Z.t13 a_116_47.t7 a_407_309.t2 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 a_116_47.t1 A.t1 VGND.t9 VNB.t17 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 VGND.t5 a_301_47.t5 a_455_47.t12 VNB.t13 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 a_407_309.t11 TE_B.t3 VPWR.t4 VPB.t10 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=940000u l=150000u
X14 VGND.t4 a_301_47.t6 a_455_47.t11 VNB.t12 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X15 a_455_47.t1 a_116_47.t8 Z.t6 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X16 VPWR.t3 TE_B.t4 a_407_309.t10 VPB.t9 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=940000u l=150000u
X17 a_455_47.t2 a_116_47.t9 Z.t5 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X18 a_455_47.t3 a_116_47.t10 Z.t4 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X19 a_301_47.t0 TE_B.t5 VGND.t0 VNB.t6 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X20 a_455_47.t10 a_301_47.t7 VGND.t3 VNB.t11 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X21 a_301_47.t1 TE_B.t6 VPWR.t8 VPB.t8 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X22 a_455_47.t9 a_301_47.t8 VGND.t2 VNB.t10 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X23 a_455_47.t8 a_301_47.t9 VGND.t1 VNB.t9 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X24 a_407_309.t3 a_116_47.t11 Z.t12 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X25 Z.t3 a_116_47.t12 a_455_47.t4 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X26 Z.t2 a_116_47.t13 a_455_47.t5 VNB.t5 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X27 VPWR.t10 A.t2 a_116_47.t2 VPB.t18 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X28 Z.t11 a_116_47.t14 a_407_309.t4 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X29 Z.t1 a_116_47.t15 a_455_47.t6 VNB.t7 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X30 a_407_309.t9 TE_B.t7 VPWR.t2 VPB.t7 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=940000u l=150000u
X31 VGND.t10 A.t3 a_116_47.t3 VNB.t18 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X32 VPWR.t1 TE_B.t8 a_407_309.t8 VPB.t6 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=940000u l=150000u
X33 a_407_309.t13 a_116_47.t16 Z.t10 VPB.t14 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X34 Z.t9 a_116_47.t17 a_407_309.t14 VPB.t15 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X35 a_407_309.t7 TE_B.t9 VPWR.t0 VPB.t5 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=940000u l=150000u
X36 a_455_47.t7 a_116_47.t18 Z.t0 VNB.t8 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X37 a_407_309.t15 a_116_47.t19 Z.t8 VPB.t16 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
R0 TE_B.n0 TE_B.t2 310.086
R1 TE_B.n7 TE_B.n6 243.482
R2 TE_B.n7 TE_B.t6 212.079
R3 TE_B.n0 TE_B.t1 175.126
R4 TE_B.n1 TE_B.t3 175.126
R5 TE_B.n2 TE_B.t4 175.126
R6 TE_B.n3 TE_B.t7 175.126
R7 TE_B.n4 TE_B.t8 175.126
R8 TE_B.n5 TE_B.t9 175.126
R9 TE_B.n6 TE_B.t0 175.126
R10 TE_B.n7 TE_B.t5 139.779
R11 TE_B.n1 TE_B.n0 134.96
R12 TE_B.n2 TE_B.n1 134.96
R13 TE_B.n3 TE_B.n2 134.96
R14 TE_B.n4 TE_B.n3 134.96
R15 TE_B.n5 TE_B.n4 134.96
R16 TE_B.n6 TE_B.n5 134.96
R17 TE_B.n8 TE_B.n7 89.966
R18 TE_B.n8 TE_B 15.092
R19 TE_B TE_B.n8 10.889
R20 a_407_309.n7 a_407_309.t6 581.673
R21 a_407_309.n9 a_407_309.n4 310.194
R22 a_407_309.n8 a_407_309.n5 310.194
R23 a_407_309.n7 a_407_309.n6 310.194
R24 a_407_309.n12 a_407_309.n11 299.02
R25 a_407_309.n10 a_407_309.n3 292.5
R26 a_407_309.n1 a_407_309.t13 191.708
R27 a_407_309.n1 a_407_309.n0 146.25
R28 a_407_309.n13 a_407_309.n2 146.25
R29 a_407_309.n15 a_407_309.n14 146.25
R30 a_407_309.n9 a_407_309.n8 63.247
R31 a_407_309.n8 a_407_309.n7 63.247
R32 a_407_309.n10 a_407_309.n9 60.664
R33 a_407_309.n3 a_407_309.t12 46.106
R34 a_407_309.n4 a_407_309.t5 28.292
R35 a_407_309.n4 a_407_309.t11 28.292
R36 a_407_309.n5 a_407_309.t10 28.292
R37 a_407_309.n5 a_407_309.t9 28.292
R38 a_407_309.n6 a_407_309.t8 28.292
R39 a_407_309.n6 a_407_309.t7 28.292
R40 a_407_309.n11 a_407_309.t4 27.713
R41 a_407_309.n2 a_407_309.t2 26.595
R42 a_407_309.n2 a_407_309.t3 26.595
R43 a_407_309.n0 a_407_309.t14 26.595
R44 a_407_309.n0 a_407_309.t15 26.595
R45 a_407_309.t0 a_407_309.n15 26.595
R46 a_407_309.n15 a_407_309.t1 26.595
R47 a_407_309.n13 a_407_309.n12 20.547
R48 a_407_309.n14 a_407_309.n1 18.863
R49 a_407_309.n14 a_407_309.n13 18.863
R50 a_407_309.n12 a_407_309.n10 7.635
R51 VPWR.n3 VPWR.n0 310.446
R52 VPWR.n12 VPWR.n11 306.463
R53 VPWR.n7 VPWR.n6 306.463
R54 VPWR.n2 VPWR.n1 306.463
R55 VPWR.n23 VPWR.t9 191.562
R56 VPWR.n19 VPWR.n18 163.183
R57 VPWR.n18 VPWR.t8 43.34
R58 VPWR.n11 VPWR.t0 28.292
R59 VPWR.n11 VPWR.t7 28.292
R60 VPWR.n6 VPWR.t2 28.292
R61 VPWR.n6 VPWR.t1 28.292
R62 VPWR.n1 VPWR.t4 28.292
R63 VPWR.n1 VPWR.t3 28.292
R64 VPWR.n0 VPWR.t5 28.292
R65 VPWR.n0 VPWR.t6 28.292
R66 VPWR.n18 VPWR.t10 26.595
R67 VPWR.n5 VPWR.n4 4.65
R68 VPWR.n8 VPWR.n7 4.65
R69 VPWR.n10 VPWR.n9 4.65
R70 VPWR.n13 VPWR.n12 4.65
R71 VPWR.n15 VPWR.n14 4.65
R72 VPWR.n17 VPWR.n16 4.65
R73 VPWR.n20 VPWR.n19 4.65
R74 VPWR.n22 VPWR.n21 4.65
R75 VPWR.n24 VPWR.n23 4.65
R76 VPWR.n3 VPWR.n2 3.895
R77 VPWR.n5 VPWR.n3 0.317
R78 VPWR.n8 VPWR.n5 0.119
R79 VPWR.n10 VPWR.n8 0.119
R80 VPWR.n13 VPWR.n10 0.119
R81 VPWR.n15 VPWR.n13 0.119
R82 VPWR.n17 VPWR.n15 0.119
R83 VPWR.n20 VPWR.n17 0.119
R84 VPWR.n22 VPWR.n20 0.119
R85 VPWR.n24 VPWR.n22 0.119
R86 VPWR VPWR.n24 0.022
R87 VPB.t8 VPB.t13 556.386
R88 VPB.t11 VPB.t4 544.548
R89 VPB.t18 VPB.t8 298.909
R90 VPB.t15 VPB.t14 248.598
R91 VPB.t16 VPB.t15 248.598
R92 VPB.t0 VPB.t16 248.598
R93 VPB.t1 VPB.t0 248.598
R94 VPB.t2 VPB.t1 248.598
R95 VPB.t3 VPB.t2 248.598
R96 VPB.t4 VPB.t3 248.598
R97 VPB.t12 VPB.t11 248.598
R98 VPB.t10 VPB.t12 248.598
R99 VPB.t9 VPB.t10 248.598
R100 VPB.t7 VPB.t9 248.598
R101 VPB.t6 VPB.t7 248.598
R102 VPB.t5 VPB.t6 248.598
R103 VPB.t13 VPB.t5 248.598
R104 VPB.t17 VPB.t18 248.598
R105 VPB VPB.t17 213.084
R106 a_301_47.n7 a_301_47.n6 300.654
R107 a_301_47.n0 a_301_47.t3 263.493
R108 a_301_47.t1 a_301_47.n7 152.349
R109 a_301_47.n5 a_301_47.n4 134.96
R110 a_301_47.n4 a_301_47.n3 134.96
R111 a_301_47.n3 a_301_47.n2 134.96
R112 a_301_47.n2 a_301_47.n1 134.96
R113 a_301_47.n1 a_301_47.n0 134.96
R114 a_301_47.n7 a_301_47.t0 134.878
R115 a_301_47.n6 a_301_47.n5 132.942
R116 a_301_47.n0 a_301_47.t2 128.533
R117 a_301_47.n1 a_301_47.t5 128.533
R118 a_301_47.n2 a_301_47.t8 128.533
R119 a_301_47.n3 a_301_47.t6 128.533
R120 a_301_47.n4 a_301_47.t9 128.533
R121 a_301_47.n5 a_301_47.t4 128.533
R122 a_301_47.n6 a_301_47.t7 126.61
R123 VGND.n3 VGND.n0 109.942
R124 VGND.n2 VGND.n1 106.463
R125 VGND.n7 VGND.n6 106.463
R126 VGND.n11 VGND.n10 106.463
R127 VGND.n21 VGND.n20 106.255
R128 VGND.n25 VGND.t9 89.58
R129 VGND.n20 VGND.t0 40.615
R130 VGND.n0 VGND.t3 24.923
R131 VGND.n0 VGND.t6 24.923
R132 VGND.n1 VGND.t1 24.923
R133 VGND.n1 VGND.t4 24.923
R134 VGND.n6 VGND.t2 24.923
R135 VGND.n6 VGND.t5 24.923
R136 VGND.n10 VGND.t8 24.923
R137 VGND.n10 VGND.t7 24.923
R138 VGND.n20 VGND.t10 24.923
R139 VGND.n26 VGND.n25 4.65
R140 VGND.n5 VGND.n4 4.65
R141 VGND.n9 VGND.n8 4.65
R142 VGND.n13 VGND.n12 4.65
R143 VGND.n15 VGND.n14 4.65
R144 VGND.n17 VGND.n16 4.65
R145 VGND.n19 VGND.n18 4.65
R146 VGND.n22 VGND.n21 4.65
R147 VGND.n24 VGND.n23 4.65
R148 VGND.n3 VGND.n2 3.488
R149 VGND.n8 VGND.n7 3.388
R150 VGND.n12 VGND.n11 0.376
R151 VGND.n5 VGND.n3 0.263
R152 VGND.n9 VGND.n5 0.119
R153 VGND.n13 VGND.n9 0.119
R154 VGND.n15 VGND.n13 0.119
R155 VGND.n17 VGND.n15 0.119
R156 VGND.n19 VGND.n17 0.119
R157 VGND.n22 VGND.n19 0.119
R158 VGND.n24 VGND.n22 0.119
R159 VGND.n26 VGND.n24 0.119
R160 VGND VGND.n26 0.022
R161 a_455_47.n4 a_455_47.t7 234.803
R162 a_455_47.t14 a_455_47.n13 173.306
R163 a_455_47.n13 a_455_47.n0 99.652
R164 a_455_47.n12 a_455_47.n1 99.652
R165 a_455_47.n11 a_455_47.n2 99.652
R166 a_455_47.n4 a_455_47.n3 92.5
R167 a_455_47.n6 a_455_47.n5 92.5
R168 a_455_47.n8 a_455_47.n7 92.5
R169 a_455_47.n10 a_455_47.n9 92.5
R170 a_455_47.n6 a_455_47.n4 56.589
R171 a_455_47.n8 a_455_47.n6 56.589
R172 a_455_47.n10 a_455_47.n8 55.343
R173 a_455_47.n12 a_455_47.n11 53.76
R174 a_455_47.n13 a_455_47.n12 53.76
R175 a_455_47.n11 a_455_47.n10 53.013
R176 a_455_47.n9 a_455_47.t10 49.846
R177 a_455_47.n9 a_455_47.t0 48
R178 a_455_47.n7 a_455_47.t4 24.923
R179 a_455_47.n7 a_455_47.t1 24.923
R180 a_455_47.n5 a_455_47.t5 24.923
R181 a_455_47.n5 a_455_47.t2 24.923
R182 a_455_47.n3 a_455_47.t6 24.923
R183 a_455_47.n3 a_455_47.t3 24.923
R184 a_455_47.n0 a_455_47.t12 24.923
R185 a_455_47.n0 a_455_47.t15 24.923
R186 a_455_47.n1 a_455_47.t11 24.923
R187 a_455_47.n1 a_455_47.t9 24.923
R188 a_455_47.n2 a_455_47.t13 24.923
R189 a_455_47.n2 a_455_47.t8 24.923
R190 VNB VNB.t17 6247.32
R191 VNB.t6 VNB.t15 5705.49
R192 VNB.t11 VNB.t0 3287.91
R193 VNB.t18 VNB.t6 2441.76
R194 VNB.t7 VNB.t8 2030.77
R195 VNB.t3 VNB.t7 2030.77
R196 VNB.t5 VNB.t3 2030.77
R197 VNB.t2 VNB.t5 2030.77
R198 VNB.t4 VNB.t2 2030.77
R199 VNB.t1 VNB.t4 2030.77
R200 VNB.t0 VNB.t1 2030.77
R201 VNB.t14 VNB.t11 2030.77
R202 VNB.t9 VNB.t14 2030.77
R203 VNB.t12 VNB.t9 2030.77
R204 VNB.t10 VNB.t12 2030.77
R205 VNB.t13 VNB.t10 2030.77
R206 VNB.t16 VNB.t13 2030.77
R207 VNB.t15 VNB.t16 2030.77
R208 VNB.t17 VNB.t18 2030.77
R209 a_116_47.n27 a_116_47.n26 361.559
R210 a_116_47.n0 a_116_47.t16 221.719
R211 a_116_47.n1 a_116_47.t17 221.719
R212 a_116_47.n2 a_116_47.t19 221.719
R213 a_116_47.n6 a_116_47.t4 221.719
R214 a_116_47.n9 a_116_47.t6 221.719
R215 a_116_47.n15 a_116_47.t7 221.719
R216 a_116_47.n21 a_116_47.t11 221.719
R217 a_116_47.n19 a_116_47.t14 221.719
R218 a_116_47.n0 a_116_47.t18 149.419
R219 a_116_47.n1 a_116_47.t15 149.419
R220 a_116_47.n2 a_116_47.t10 149.419
R221 a_116_47.n6 a_116_47.t13 149.419
R222 a_116_47.n9 a_116_47.t9 149.419
R223 a_116_47.n15 a_116_47.t12 149.419
R224 a_116_47.n21 a_116_47.t8 149.419
R225 a_116_47.n19 a_116_47.t5 149.419
R226 a_116_47.n26 a_116_47.n25 143.034
R227 a_116_47.n5 a_116_47.n4 76
R228 a_116_47.n8 a_116_47.n7 76
R229 a_116_47.n11 a_116_47.n10 76
R230 a_116_47.n1 a_116_47.n0 74.977
R231 a_116_47.n21 a_116_47.n20 51.77
R232 a_116_47.n17 a_116_47.n16 49.092
R233 a_116_47.n5 a_116_47.n3 48.26
R234 a_116_47.n7 a_116_47.n6 33.918
R235 a_116_47.n3 a_116_47.n2 32.544
R236 a_116_47.n27 a_116_47.t2 26.595
R237 a_116_47.t0 a_116_47.n27 26.595
R238 a_116_47.n3 a_116_47.n1 26.425
R239 a_116_47.n25 a_116_47.t3 24.923
R240 a_116_47.n25 a_116_47.t1 24.923
R241 a_116_47.n20 a_116_47.n19 23.207
R242 a_116_47.n10 a_116_47.n9 19.637
R243 a_116_47.n8 a_116_47.n5 17.408
R244 a_116_47.n11 a_116_47.n8 17.408
R245 a_116_47.n12 a_116_47.n11 17.408
R246 a_116_47.n13 a_116_47.n12 14.08
R247 a_116_47.n18 a_116_47.n17 11.603
R248 a_116_47.n26 a_116_47.n24 11.563
R249 a_116_47.n23 a_116_47.n22 9.3
R250 a_116_47.n16 a_116_47.n15 5.355
R251 a_116_47.n22 a_116_47.n21 5.355
R252 a_116_47.n22 a_116_47.n18 3.57
R253 a_116_47.n14 a_116_47.n13 3.328
R254 a_116_47.n24 a_116_47.n23 1.194
R255 a_116_47.n23 a_116_47.n14 1.024
R256 Z.n7 Z.n0 292.5
R257 Z.n6 Z.n1 292.5
R258 Z.n5 Z.n2 292.5
R259 Z.n4 Z.n3 292.5
R260 Z.n12 Z.n11 137.3
R261 Z.n12 Z.n10 92.5
R262 Z.n13 Z.n9 92.5
R263 Z.n14 Z.n8 92.5
R264 Z.n14 Z.n13 44.8
R265 Z.n13 Z.n12 44.8
R266 Z Z.n4 27.428
R267 Z.n3 Z.t12 26.595
R268 Z.n3 Z.t11 26.595
R269 Z.n2 Z.t14 26.595
R270 Z.n2 Z.t13 26.595
R271 Z.n1 Z.t8 26.595
R272 Z.n1 Z.t15 26.595
R273 Z.n0 Z.t10 26.595
R274 Z.n0 Z.t9 26.595
R275 Z.n8 Z.t0 24.923
R276 Z.n8 Z.t1 24.923
R277 Z.n9 Z.t4 24.923
R278 Z.n9 Z.t2 24.923
R279 Z.n10 Z.t5 24.923
R280 Z.n10 Z.t3 24.923
R281 Z.n11 Z.t6 24.923
R282 Z.n11 Z.t7 24.923
R283 Z Z.n14 21.002
R284 Z Z.n7 17.371
R285 Z.n4 Z 14.628
R286 Z Z.n6 13.714
R287 Z.n5 Z 10.971
R288 Z Z.n5 10.057
R289 Z.n6 Z 7.314
R290 Z.n7 Z 3.657
R291 A.n1 A.t0 231.014
R292 A.n0 A.t2 221.719
R293 A.n1 A.t1 158.714
R294 A.n0 A.t3 149.419
R295 A.n2 A.n1 76
R296 A.n1 A.n0 61.588
R297 A.n2 A 10.573
R298 A A.n2 2.04
C0 VPWR VGND 0.10fF
C1 TE_B VPWR 0.11fF
C2 VPB TE_B 0.11fF
C3 VPB VPWR 0.18fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__edfxbp_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__edfxbp_1 VPWR VGND CLK Q_N DE D Q VNB VPB
X0 a_381_369.t0 D.t0 a_299_47.t2 VPB.t9 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1 Q.t0 a_1591_413.t4 VGND.t0 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 VPWR.t7 DE.t0 a_423_343.t1 VPB.t6 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X3 VPWR.t9 CLK.t0 a_27_47.t1 VPB.t14 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X4 a_1591_413.t0 a_193_47.t2 a_1514_47.t0 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X5 Q_N.t1 a_791_264.t2 VPWR.t4 VPB.t10 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 a_986_413.t3 a_193_47.t3 a_299_47.t0 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7 a_1101_47.t0 a_193_47.t4 a_986_413.t2 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X8 VGND.t3 DE.t1 a_423_343.t0 VNB.t7 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9 a_1500_413.t0 a_1150_159.t2 VPWR.t3 VPB.t8 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10 a_1514_47.t1 a_1150_159.t3 VGND.t9 VNB.t15 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11 Q.t1 a_1591_413.t5 VPWR.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 a_1675_413.t0 a_193_47.t5 a_1591_413.t1 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13 VPWR.t1 a_1591_413.t6 a_791_264.t1 VPB.t13 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X14 a_193_47.t0 a_27_47.t2 VGND.t2 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15 a_1591_413.t2 a_27_47.t3 a_1500_413.t1 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16 a_729_47.t0 a_423_343.t2 VGND.t11 VNB.t17 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17 a_729_369.t0 DE.t2 VPWR.t6 VPB.t7 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X18 a_1077_413.t1 a_27_47.t4 a_986_413.t1 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19 VPWR.t5 a_791_264.t3 a_1675_413.t1 VPB.t11 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20 a_299_47.t4 a_791_264.t4 a_729_47.t1 VNB.t9 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21 VGND.t4 a_791_264.t5 a_1717_47.t1 VNB.t10 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22 a_193_47.t1 a_27_47.t5 VPWR.t2 VPB.t5 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X23 a_1717_47.t0 a_27_47.t6 a_1591_413.t3 VNB.t5 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X24 VPWR.t11 a_1150_159.t4 a_1077_413.t0 VPB.t16 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X25 a_1150_159.t1 a_986_413.t4 VPWR.t10 VPB.t15 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X26 a_986_413.t0 a_27_47.t7 a_299_47.t1 VNB.t6 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X27 a_299_47.t5 a_791_264.t6 a_729_369.t1 VPB.t12 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X28 VGND.t1 a_1591_413.t7 a_791_264.t0 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X29 a_381_47.t0 D.t1 a_299_47.t3 VNB.t8 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X30 VGND.t10 a_1150_159.t5 a_1101_47.t1 VNB.t16 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X31 VPWR.t8 a_423_343.t3 a_381_369.t1 VPB.t17 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X32 VGND.t7 CLK.t1 a_27_47.t0 VNB.t13 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X33 VGND.t6 DE.t3 a_381_47.t1 VNB.t12 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X34 a_1150_159.t0 a_986_413.t5 VGND.t8 VNB.t14 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X35 Q_N.t0 a_791_264.t7 VGND.t5 VNB.t11 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
R0 D.n0 D.t1 216.76
R1 D.n0 D.t0 215.106
R2 D D.n0 34.479
R3 a_299_47.t2 a_299_47.n3 321.627
R4 a_299_47.n2 a_299_47.n0 234.198
R5 a_299_47.n0 a_299_47.t0 231.018
R6 a_299_47.n1 a_299_47.t1 206.236
R7 a_299_47.n3 a_299_47.t3 139.932
R8 a_299_47.n0 a_299_47.t5 41.167
R9 a_299_47.n1 a_299_47.t4 26.96
R10 a_299_47.n2 a_299_47.n1 8.417
R11 a_299_47.n3 a_299_47.n2 8.177
R12 a_381_369.t0 a_381_369.t1 64.64
R13 VPB.t10 VPB.t13 787.227
R14 VPB.t15 VPB.t8 556.386
R15 VPB.t17 VPB.t6 556.386
R16 VPB.t5 VPB.t9 556.386
R17 VPB.t12 VPB.t1 458.722
R18 VPB.t16 VPB.t15 390.654
R19 VPB.t2 VPB.t11 337.383
R20 VPB.t4 VPB.t16 304.828
R21 VPB.t7 VPB.t12 301.869
R22 VPB.t13 VPB.t0 287.071
R23 VPB.t11 VPB.t10 287.071
R24 VPB.t8 VPB.t3 269.314
R25 VPB.t1 VPB.t4 269.314
R26 VPB.t6 VPB.t7 260.436
R27 VPB.t3 VPB.t2 248.598
R28 VPB.t14 VPB.t5 248.598
R29 VPB.t9 VPB.t17 213.084
R30 VPB VPB.t14 142.056
R31 a_1591_413.n5 a_1591_413.n4 349.52
R32 a_1591_413.n0 a_1591_413.t5 212.079
R33 a_1591_413.n4 a_1591_413.n3 193.388
R34 a_1591_413.n1 a_1591_413.t7 176.733
R35 a_1591_413.n4 a_1591_413.n2 176.238
R36 a_1591_413.n2 a_1591_413.t6 163.879
R37 a_1591_413.n0 a_1591_413.t4 139.779
R38 a_1591_413.n3 a_1591_413.t3 76.666
R39 a_1591_413.n1 a_1591_413.n0 70.839
R40 a_1591_413.t1 a_1591_413.n5 63.321
R41 a_1591_413.n5 a_1591_413.t2 63.321
R42 a_1591_413.n3 a_1591_413.t0 50
R43 a_1591_413.n2 a_1591_413.n1 33.74
R44 VGND.n12 VGND.t9 152.016
R45 VGND.n35 VGND.t6 145.81
R46 VGND.n31 VGND.n30 109.76
R47 VGND.n44 VGND.n43 107.239
R48 VGND.n18 VGND.n17 106.11
R49 VGND.n3 VGND.n0 74.893
R50 VGND.n17 VGND.t8 74.865
R51 VGND.n2 VGND.n1 70.639
R52 VGND.n1 VGND.t4 57.782
R53 VGND.n0 VGND.t1 57.781
R54 VGND.n30 VGND.t11 41.428
R55 VGND.n30 VGND.t3 41.428
R56 VGND.n17 VGND.t10 40
R57 VGND.n43 VGND.t2 38.571
R58 VGND.n43 VGND.t7 38.571
R59 VGND.n0 VGND.t0 24.78
R60 VGND.n1 VGND.t5 24.778
R61 VGND.n3 VGND.n2 10.535
R62 VGND.n5 VGND.n4 4.65
R63 VGND.n7 VGND.n6 4.65
R64 VGND.n9 VGND.n8 4.65
R65 VGND.n11 VGND.n10 4.65
R66 VGND.n14 VGND.n13 4.65
R67 VGND.n16 VGND.n15 4.65
R68 VGND.n19 VGND.n18 4.65
R69 VGND.n21 VGND.n20 4.65
R70 VGND.n23 VGND.n22 4.65
R71 VGND.n25 VGND.n24 4.65
R72 VGND.n27 VGND.n26 4.65
R73 VGND.n29 VGND.n28 4.65
R74 VGND.n32 VGND.n31 4.65
R75 VGND.n34 VGND.n33 4.65
R76 VGND.n36 VGND.n35 4.65
R77 VGND.n38 VGND.n37 4.65
R78 VGND.n40 VGND.n39 4.65
R79 VGND.n42 VGND.n41 4.65
R80 VGND.n45 VGND.n44 3.932
R81 VGND.n13 VGND.n12 2.635
R82 VGND.n5 VGND.n3 0.138
R83 VGND.n45 VGND.n42 0.137
R84 VGND VGND.n45 0.123
R85 VGND.n7 VGND.n5 0.119
R86 VGND.n9 VGND.n7 0.119
R87 VGND.n11 VGND.n9 0.119
R88 VGND.n14 VGND.n11 0.119
R89 VGND.n16 VGND.n14 0.119
R90 VGND.n19 VGND.n16 0.119
R91 VGND.n21 VGND.n19 0.119
R92 VGND.n23 VGND.n21 0.119
R93 VGND.n25 VGND.n23 0.119
R94 VGND.n27 VGND.n25 0.119
R95 VGND.n29 VGND.n27 0.119
R96 VGND.n32 VGND.n29 0.119
R97 VGND.n34 VGND.n32 0.119
R98 VGND.n36 VGND.n34 0.119
R99 VGND.n38 VGND.n36 0.119
R100 VGND.n40 VGND.n38 0.119
R101 VGND.n42 VGND.n40 0.119
R102 Q Q.t1 153.46
R103 Q Q.t0 100.27
R104 VNB.t9 VNB.t6 6166.89
R105 VNB.t12 VNB.t7 6082.35
R106 VNB.t4 VNB.t8 6082.35
R107 VNB.t11 VNB.t2 5874.73
R108 VNB.t14 VNB.t15 5346.86
R109 VNB VNB.t13 4270.59
R110 VNB.t1 VNB.t16 3476.38
R111 VNB.t0 VNB.t5 3429.41
R112 VNB.t17 VNB.t9 3300
R113 VNB.t15 VNB.t0 3138.24
R114 VNB.t16 VNB.t14 3130.33
R115 VNB.t6 VNB.t1 3122.58
R116 VNB.t5 VNB.t10 3073.53
R117 VNB.t7 VNB.t17 2847.06
R118 VNB.t13 VNB.t4 2717.65
R119 VNB.t2 VNB.t3 2345.05
R120 VNB.t8 VNB.t12 2329.41
R121 VNB.t10 VNB.t11 2303.7
R122 DE.n0 DE.t2 319.725
R123 DE.n2 DE.n1 238.689
R124 DE.n0 DE.t0 178.339
R125 DE.n1 DE.n0 147.813
R126 DE.n2 DE.t3 130.384
R127 DE.n1 DE.t1 130.14
R128 DE DE.n2 82.892
R129 a_423_343.n1 a_423_343.t3 299.566
R130 a_423_343.n0 a_423_343.t2 258.036
R131 a_423_343.t1 a_423_343.n1 230.699
R132 a_423_343.n0 a_423_343.t0 151.679
R133 a_423_343.n1 a_423_343.n0 11.133
R134 VPWR.n12 VPWR.t3 375.462
R135 VPWR.n43 VPWR.n42 311.893
R136 VPWR.n34 VPWR.t8 228.681
R137 VPWR.n30 VPWR.n29 176.72
R138 VPWR.n17 VPWR.n16 171.436
R139 VPWR.n1 VPWR.n0 143.182
R140 VPWR.n3 VPWR.n2 132.968
R141 VPWR.n16 VPWR.t11 106.098
R142 VPWR.n2 VPWR.t5 95.255
R143 VPWR.n0 VPWR.t1 61.912
R144 VPWR.n29 VPWR.t6 44.632
R145 VPWR.n29 VPWR.t7 44.632
R146 VPWR.n16 VPWR.t10 43.34
R147 VPWR.n42 VPWR.t2 41.554
R148 VPWR.n42 VPWR.t9 41.554
R149 VPWR.n0 VPWR.t0 30.241
R150 VPWR.n2 VPWR.t4 26.498
R151 VPWR.n4 VPWR.n3 13.176
R152 VPWR.n5 VPWR.n4 4.65
R153 VPWR.n7 VPWR.n6 4.65
R154 VPWR.n9 VPWR.n8 4.65
R155 VPWR.n11 VPWR.n10 4.65
R156 VPWR.n13 VPWR.n12 4.65
R157 VPWR.n15 VPWR.n14 4.65
R158 VPWR.n18 VPWR.n17 4.65
R159 VPWR.n20 VPWR.n19 4.65
R160 VPWR.n22 VPWR.n21 4.65
R161 VPWR.n24 VPWR.n23 4.65
R162 VPWR.n26 VPWR.n25 4.65
R163 VPWR.n28 VPWR.n27 4.65
R164 VPWR.n31 VPWR.n30 4.65
R165 VPWR.n33 VPWR.n32 4.65
R166 VPWR.n35 VPWR.n34 4.65
R167 VPWR.n37 VPWR.n36 4.65
R168 VPWR.n39 VPWR.n38 4.65
R169 VPWR.n41 VPWR.n40 4.65
R170 VPWR.n44 VPWR.n43 3.932
R171 VPWR.n5 VPWR.n1 0.139
R172 VPWR.n44 VPWR.n41 0.137
R173 VPWR VPWR.n44 0.123
R174 VPWR.n7 VPWR.n5 0.119
R175 VPWR.n9 VPWR.n7 0.119
R176 VPWR.n11 VPWR.n9 0.119
R177 VPWR.n13 VPWR.n11 0.119
R178 VPWR.n15 VPWR.n13 0.119
R179 VPWR.n18 VPWR.n15 0.119
R180 VPWR.n20 VPWR.n18 0.119
R181 VPWR.n22 VPWR.n20 0.119
R182 VPWR.n24 VPWR.n22 0.119
R183 VPWR.n26 VPWR.n24 0.119
R184 VPWR.n28 VPWR.n26 0.119
R185 VPWR.n31 VPWR.n28 0.119
R186 VPWR.n33 VPWR.n31 0.119
R187 VPWR.n35 VPWR.n33 0.119
R188 VPWR.n37 VPWR.n35 0.119
R189 VPWR.n39 VPWR.n37 0.119
R190 VPWR.n41 VPWR.n39 0.119
R191 CLK.n0 CLK.t0 292.947
R192 CLK.n0 CLK.t1 209.401
R193 CLK CLK.n0 78.067
R194 a_27_47.n1 a_27_47.t6 443.438
R195 a_27_47.n0 a_27_47.t7 269.985
R196 a_27_47.n3 a_27_47.t5 263.405
R197 a_27_47.n1 a_27_47.t3 254.388
R198 a_27_47.t1 a_27_47.n5 244.156
R199 a_27_47.n3 a_27_47.t2 228.059
R200 a_27_47.n4 a_27_47.t0 195.871
R201 a_27_47.n0 a_27_47.t4 142.49
R202 a_27_47.n2 a_27_47.n1 113.844
R203 a_27_47.n4 a_27_47.n3 76
R204 a_27_47.n5 a_27_47.n4 35.339
R205 a_27_47.n5 a_27_47.n2 8.636
R206 a_27_47.n2 a_27_47.n0 2.9
R207 a_193_47.n1 a_193_47.t4 389.542
R208 a_193_47.n1 a_193_47.t3 273.571
R209 a_193_47.t1 a_193_47.n3 249.337
R210 a_193_47.n0 a_193_47.t5 232.651
R211 a_193_47.n0 a_193_47.t2 222.372
R212 a_193_47.n3 a_193_47.t0 207.871
R213 a_193_47.n2 a_193_47.n1 93.104
R214 a_193_47.n3 a_193_47.n2 7.926
R215 a_193_47.n2 a_193_47.n0 7.6
R216 a_1514_47.n0 a_1514_47.t0 70
R217 a_1514_47.n0 a_1514_47.t1 26.393
R218 a_1514_47.n1 a_1514_47.n0 14.4
R219 a_791_264.n0 a_791_264.t3 368.968
R220 a_791_264.n3 a_791_264.t4 310.621
R221 a_791_264.t1 a_791_264.n5 248.537
R222 a_791_264.n1 a_791_264.t2 245.819
R223 a_791_264.n5 a_791_264.n2 232.442
R224 a_791_264.n3 a_791_264.t6 194.941
R225 a_791_264.n0 a_791_264.t5 189.586
R226 a_791_264.n2 a_791_264.t7 152.633
R227 a_791_264.n4 a_791_264.t0 148.576
R228 a_791_264.n4 a_791_264.n3 134.221
R229 a_791_264.n1 a_791_264.n0 96.4
R230 a_791_264.n2 a_791_264.n1 29.962
R231 a_791_264.n5 a_791_264.n4 7.717
R232 Q_N Q_N.t1 148.433
R233 Q_N Q_N.t0 102.677
R234 a_986_413.n3 a_986_413.n2 388.236
R235 a_986_413.n0 a_986_413.t5 230.482
R236 a_986_413.n0 a_986_413.t4 196.013
R237 a_986_413.n2 a_986_413.n1 183.768
R238 a_986_413.n2 a_986_413.n0 95.938
R239 a_986_413.t1 a_986_413.n3 72.702
R240 a_986_413.n3 a_986_413.t3 70.357
R241 a_986_413.n1 a_986_413.t2 51.666
R242 a_986_413.n1 a_986_413.t0 45
R243 a_1101_47.t1 a_1101_47.t0 111.393
R244 a_1150_159.n1 a_1150_159.t4 406.399
R245 a_1150_159.n0 a_1150_159.t2 318.12
R246 a_1150_159.t1 a_1150_159.n3 262.563
R247 a_1150_159.n0 a_1150_159.t3 194.476
R248 a_1150_159.n1 a_1150_159.t5 130.052
R249 a_1150_159.n2 a_1150_159.n1 100.533
R250 a_1150_159.n2 a_1150_159.t0 93.987
R251 a_1150_159.n3 a_1150_159.n0 92.484
R252 a_1150_159.n3 a_1150_159.n2 9.323
R253 a_1500_413.t0 a_1500_413.t1 143.059
R254 a_1675_413.t0 a_1675_413.t1 197
R255 a_729_47.t0 a_729_47.t1 102.857
R256 a_729_369.t0 a_729_369.t1 110.812
R257 a_1077_413.t0 a_1077_413.t1 171.202
R258 a_1717_47.t1 a_1717_47.t0 93.059
R259 a_381_47.t0 a_381_47.t1 60
C0 VPWR VPB 0.26fF
C1 VGND Q 0.17fF
C2 VGND Q_N 0.17fF
C3 D DE 0.13fF
C4 VPWR VGND 0.14fF
C5 VPWR Q 0.21fF
C6 VPWR Q_N 0.16fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__edfxtp_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__edfxtp_1 VPWR VGND CLK DE D Q VNB VPB
X0 a_381_369.t0 D.t0 a_299_47.t2 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1 VGND.t3 a_1591_413.t4 a_791_264.t0 VNB.t8 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 VPWR.t9 DE.t0 a_423_343.t1 VPB.t7 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X3 VPWR.t7 CLK.t0 a_27_47.t1 VPB.t14 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X4 a_1591_413.t0 a_193_47.t2 a_1514_47.t0 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X5 a_986_413.t3 a_193_47.t3 a_299_47.t4 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 a_1101_47.t0 a_193_47.t4 a_986_413.t2 VNB.t5 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X7 Q.t1 a_1591_413.t5 VPWR.t3 VPB.t15 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 VGND.t5 DE.t1 a_423_343.t0 VNB.t9 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9 a_1500_413.t1 a_1150_159.t2 VPWR.t4 VPB.t9 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10 a_1514_47.t1 a_1150_159.t3 VGND.t7 VNB.t11 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11 a_1675_413.t0 a_193_47.t5 a_1591_413.t1 VPB.t5 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12 a_193_47.t0 a_27_47.t2 VGND.t9 VNB.t13 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13 a_1591_413.t2 a_27_47.t3 a_1500_413.t0 VPB.t11 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14 a_729_47.t1 a_423_343.t2 VGND.t2 VNB.t6 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15 a_729_369.t1 DE.t2 VPWR.t8 VPB.t8 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X16 a_1077_413.t0 a_27_47.t4 a_986_413.t0 VPB.t12 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17 VPWR.t1 a_791_264.t2 a_1675_413.t1 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18 Q.t0 a_1591_413.t6 VGND.t4 VNB.t7 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X19 a_299_47.t0 a_791_264.t3 a_729_47.t0 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20 VPWR.t2 a_1591_413.t7 a_791_264.t1 VPB.t16 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X21 VGND.t1 a_791_264.t4 a_1717_47.t1 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22 a_193_47.t1 a_27_47.t5 VPWR.t6 VPB.t13 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X23 a_1717_47.t0 a_27_47.t6 a_1591_413.t3 VNB.t14 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X24 VPWR.t5 a_1150_159.t4 a_1077_413.t1 VPB.t10 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X25 a_1150_159.t1 a_986_413.t4 VPWR.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X26 a_986_413.t1 a_27_47.t7 a_299_47.t5 VNB.t15 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X27 a_299_47.t1 a_791_264.t5 a_729_369.t0 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X28 a_381_47.t0 D.t1 a_299_47.t3 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X29 VGND.t8 a_1150_159.t5 a_1101_47.t1 VNB.t12 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X30 VPWR.t10 a_423_343.t3 a_381_369.t1 VPB.t6 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X31 VGND.t10 CLK.t1 a_27_47.t0 VNB.t16 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X32 VGND.t6 DE.t3 a_381_47.t1 VNB.t10 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X33 a_1150_159.t0 a_986_413.t5 VGND.t0 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
R0 D.n0 D.t1 216.76
R1 D.n0 D.t0 215.106
R2 D D.n0 34.479
R3 a_299_47.n1 a_299_47.t2 321.627
R4 a_299_47.n3 a_299_47.n2 244.917
R5 a_299_47.n3 a_299_47.t4 230.936
R6 a_299_47.n0 a_299_47.t5 206.236
R7 a_299_47.n1 a_299_47.t3 139.932
R8 a_299_47.t1 a_299_47.n3 35.02
R9 a_299_47.n0 a_299_47.t0 26.96
R10 a_299_47.n2 a_299_47.n0 8.417
R11 a_299_47.n2 a_299_47.n1 8.177
R12 a_381_369.t0 a_381_369.t1 64.64
R13 VPB.t1 VPB.t16 624.454
R14 VPB.t0 VPB.t9 556.386
R15 VPB.t6 VPB.t7 556.386
R16 VPB.t13 VPB.t3 556.386
R17 VPB.t2 VPB.t4 458.722
R18 VPB.t10 VPB.t0 390.654
R19 VPB.t5 VPB.t1 337.383
R20 VPB.t12 VPB.t10 304.828
R21 VPB.t8 VPB.t2 301.869
R22 VPB.t16 VPB.t15 287.071
R23 VPB.t9 VPB.t11 269.314
R24 VPB.t4 VPB.t12 269.314
R25 VPB.t7 VPB.t8 260.436
R26 VPB.t11 VPB.t5 248.598
R27 VPB.t14 VPB.t13 248.598
R28 VPB.t3 VPB.t6 213.084
R29 VPB VPB.t14 142.056
R30 a_1591_413.n4 a_1591_413.n3 398.525
R31 a_1591_413.n2 a_1591_413.t7 269.919
R32 a_1591_413.n1 a_1591_413.t5 212.079
R33 a_1591_413.n2 a_1591_413.t4 176.733
R34 a_1591_413.n3 a_1591_413.n2 176.181
R35 a_1591_413.n3 a_1591_413.n0 159.603
R36 a_1591_413.n1 a_1591_413.t6 139.779
R37 a_1591_413.n0 a_1591_413.t3 76.666
R38 a_1591_413.n2 a_1591_413.n1 70.839
R39 a_1591_413.t1 a_1591_413.n4 63.321
R40 a_1591_413.n4 a_1591_413.t2 63.321
R41 a_1591_413.n0 a_1591_413.t0 50
R42 a_791_264.n2 a_791_264.t4 382.743
R43 a_791_264.n0 a_791_264.t3 310.621
R44 a_791_264.t1 a_791_264.n3 216.537
R45 a_791_264.n0 a_791_264.t5 194.941
R46 a_791_264.n1 a_791_264.t0 149.821
R47 a_791_264.n2 a_791_264.t2 138.53
R48 a_791_264.n1 a_791_264.n0 133.605
R49 a_791_264.n3 a_791_264.n2 98.016
R50 a_791_264.n3 a_791_264.n1 48.37
R51 VGND.n11 VGND.t7 152.016
R52 VGND.n0 VGND.t1 149.356
R53 VGND.n34 VGND.t6 145.81
R54 VGND.n30 VGND.n29 109.76
R55 VGND.n43 VGND.n42 107.239
R56 VGND.n17 VGND.n16 106.11
R57 VGND.n2 VGND.n1 76.596
R58 VGND.n16 VGND.t0 74.865
R59 VGND.n1 VGND.t3 57.781
R60 VGND.n29 VGND.t2 41.428
R61 VGND.n29 VGND.t5 41.428
R62 VGND.n16 VGND.t8 40
R63 VGND.n42 VGND.t9 38.571
R64 VGND.n42 VGND.t10 38.571
R65 VGND.n1 VGND.t4 24.78
R66 VGND.n2 VGND.n0 8.863
R67 VGND.n4 VGND.n3 4.65
R68 VGND.n6 VGND.n5 4.65
R69 VGND.n8 VGND.n7 4.65
R70 VGND.n10 VGND.n9 4.65
R71 VGND.n13 VGND.n12 4.65
R72 VGND.n15 VGND.n14 4.65
R73 VGND.n18 VGND.n17 4.65
R74 VGND.n20 VGND.n19 4.65
R75 VGND.n22 VGND.n21 4.65
R76 VGND.n24 VGND.n23 4.65
R77 VGND.n26 VGND.n25 4.65
R78 VGND.n28 VGND.n27 4.65
R79 VGND.n31 VGND.n30 4.65
R80 VGND.n33 VGND.n32 4.65
R81 VGND.n35 VGND.n34 4.65
R82 VGND.n37 VGND.n36 4.65
R83 VGND.n39 VGND.n38 4.65
R84 VGND.n41 VGND.n40 4.65
R85 VGND.n44 VGND.n43 3.932
R86 VGND.n12 VGND.n11 2.635
R87 VGND.n4 VGND.n2 0.3
R88 VGND.n44 VGND.n41 0.137
R89 VGND VGND.n44 0.123
R90 VGND.n6 VGND.n4 0.119
R91 VGND.n8 VGND.n6 0.119
R92 VGND.n10 VGND.n8 0.119
R93 VGND.n13 VGND.n10 0.119
R94 VGND.n15 VGND.n13 0.119
R95 VGND.n18 VGND.n15 0.119
R96 VGND.n20 VGND.n18 0.119
R97 VGND.n22 VGND.n20 0.119
R98 VGND.n24 VGND.n22 0.119
R99 VGND.n26 VGND.n24 0.119
R100 VGND.n28 VGND.n26 0.119
R101 VGND.n31 VGND.n28 0.119
R102 VGND.n33 VGND.n31 0.119
R103 VGND.n35 VGND.n33 0.119
R104 VGND.n37 VGND.n35 0.119
R105 VGND.n39 VGND.n37 0.119
R106 VGND.n41 VGND.n39 0.119
R107 VNB.t3 VNB.t15 6166.89
R108 VNB.t2 VNB.t8 6082.35
R109 VNB.t10 VNB.t9 6082.35
R110 VNB.t13 VNB.t1 6082.35
R111 VNB.t0 VNB.t11 5346.86
R112 VNB VNB.t16 4270.59
R113 VNB.t5 VNB.t12 3476.38
R114 VNB.t4 VNB.t14 3429.41
R115 VNB.t6 VNB.t3 3300
R116 VNB.t11 VNB.t4 3138.24
R117 VNB.t12 VNB.t0 3130.33
R118 VNB.t15 VNB.t5 3122.58
R119 VNB.t14 VNB.t2 3073.53
R120 VNB.t9 VNB.t6 2847.06
R121 VNB.t16 VNB.t13 2717.65
R122 VNB.t1 VNB.t10 2329.41
R123 VNB.t8 VNB.t7 2303.7
R124 DE.n0 DE.t2 319.725
R125 DE.n2 DE.n1 238.689
R126 DE.n0 DE.t0 178.339
R127 DE.n1 DE.n0 147.813
R128 DE.n2 DE.t3 130.384
R129 DE.n1 DE.t1 130.14
R130 DE DE.n2 82.892
R131 a_423_343.n1 a_423_343.t3 299.566
R132 a_423_343.n0 a_423_343.t2 258.036
R133 a_423_343.t1 a_423_343.n1 230.699
R134 a_423_343.n0 a_423_343.t0 151.679
R135 a_423_343.n1 a_423_343.n0 11.133
R136 VPWR.n2 VPWR.t1 378.842
R137 VPWR.n11 VPWR.t4 375.462
R138 VPWR.n42 VPWR.n41 311.893
R139 VPWR.n33 VPWR.t10 228.681
R140 VPWR.n29 VPWR.n28 176.72
R141 VPWR.n16 VPWR.n15 171.436
R142 VPWR.n1 VPWR.n0 144.883
R143 VPWR.n15 VPWR.t5 106.098
R144 VPWR.n0 VPWR.t2 61.912
R145 VPWR.n28 VPWR.t8 44.632
R146 VPWR.n28 VPWR.t9 44.632
R147 VPWR.n15 VPWR.t0 43.34
R148 VPWR.n41 VPWR.t6 41.554
R149 VPWR.n41 VPWR.t7 41.554
R150 VPWR.n0 VPWR.t3 30.241
R151 VPWR.n4 VPWR.n3 4.65
R152 VPWR.n6 VPWR.n5 4.65
R153 VPWR.n8 VPWR.n7 4.65
R154 VPWR.n10 VPWR.n9 4.65
R155 VPWR.n12 VPWR.n11 4.65
R156 VPWR.n14 VPWR.n13 4.65
R157 VPWR.n17 VPWR.n16 4.65
R158 VPWR.n19 VPWR.n18 4.65
R159 VPWR.n21 VPWR.n20 4.65
R160 VPWR.n23 VPWR.n22 4.65
R161 VPWR.n25 VPWR.n24 4.65
R162 VPWR.n27 VPWR.n26 4.65
R163 VPWR.n30 VPWR.n29 4.65
R164 VPWR.n32 VPWR.n31 4.65
R165 VPWR.n34 VPWR.n33 4.65
R166 VPWR.n36 VPWR.n35 4.65
R167 VPWR.n38 VPWR.n37 4.65
R168 VPWR.n40 VPWR.n39 4.65
R169 VPWR.n43 VPWR.n42 3.932
R170 VPWR.n3 VPWR.n2 0.752
R171 VPWR.n4 VPWR.n1 0.3
R172 VPWR.n43 VPWR.n40 0.137
R173 VPWR VPWR.n43 0.123
R174 VPWR.n6 VPWR.n4 0.119
R175 VPWR.n8 VPWR.n6 0.119
R176 VPWR.n10 VPWR.n8 0.119
R177 VPWR.n12 VPWR.n10 0.119
R178 VPWR.n14 VPWR.n12 0.119
R179 VPWR.n17 VPWR.n14 0.119
R180 VPWR.n19 VPWR.n17 0.119
R181 VPWR.n21 VPWR.n19 0.119
R182 VPWR.n23 VPWR.n21 0.119
R183 VPWR.n25 VPWR.n23 0.119
R184 VPWR.n27 VPWR.n25 0.119
R185 VPWR.n30 VPWR.n27 0.119
R186 VPWR.n32 VPWR.n30 0.119
R187 VPWR.n34 VPWR.n32 0.119
R188 VPWR.n36 VPWR.n34 0.119
R189 VPWR.n38 VPWR.n36 0.119
R190 VPWR.n40 VPWR.n38 0.119
R191 CLK.n0 CLK.t0 292.947
R192 CLK.n0 CLK.t1 209.401
R193 CLK CLK.n0 78.067
R194 a_27_47.n1 a_27_47.t6 443.438
R195 a_27_47.n0 a_27_47.t7 269.985
R196 a_27_47.n3 a_27_47.t5 263.405
R197 a_27_47.n1 a_27_47.t3 254.388
R198 a_27_47.t1 a_27_47.n5 244.156
R199 a_27_47.n3 a_27_47.t2 228.059
R200 a_27_47.n4 a_27_47.t0 195.871
R201 a_27_47.n0 a_27_47.t4 142.49
R202 a_27_47.n2 a_27_47.n1 113.844
R203 a_27_47.n4 a_27_47.n3 76
R204 a_27_47.n5 a_27_47.n4 35.339
R205 a_27_47.n5 a_27_47.n2 8.636
R206 a_27_47.n2 a_27_47.n0 2.9
R207 a_193_47.n1 a_193_47.t4 389.542
R208 a_193_47.n1 a_193_47.t3 273.571
R209 a_193_47.t1 a_193_47.n3 249.337
R210 a_193_47.n0 a_193_47.t5 232.651
R211 a_193_47.n0 a_193_47.t2 222.372
R212 a_193_47.n3 a_193_47.t0 207.871
R213 a_193_47.n2 a_193_47.n1 93.104
R214 a_193_47.n3 a_193_47.n2 7.926
R215 a_193_47.n2 a_193_47.n0 7.6
R216 a_1514_47.n0 a_1514_47.t0 70
R217 a_1514_47.n0 a_1514_47.t1 26.393
R218 a_1514_47.n1 a_1514_47.n0 14.4
R219 a_986_413.n3 a_986_413.n2 388.236
R220 a_986_413.n0 a_986_413.t5 230.482
R221 a_986_413.n0 a_986_413.t4 196.013
R222 a_986_413.n2 a_986_413.n1 183.768
R223 a_986_413.n2 a_986_413.n0 95.938
R224 a_986_413.t0 a_986_413.n3 72.702
R225 a_986_413.n3 a_986_413.t3 70.357
R226 a_986_413.n1 a_986_413.t2 51.666
R227 a_986_413.n1 a_986_413.t1 45
R228 a_1101_47.t1 a_1101_47.t0 111.393
R229 Q Q.t1 153.46
R230 Q Q.t0 100.27
R231 a_1150_159.n1 a_1150_159.t4 406.399
R232 a_1150_159.n0 a_1150_159.t2 318.12
R233 a_1150_159.t1 a_1150_159.n3 262.563
R234 a_1150_159.n0 a_1150_159.t3 194.476
R235 a_1150_159.n1 a_1150_159.t5 130.052
R236 a_1150_159.n2 a_1150_159.n1 100.533
R237 a_1150_159.n2 a_1150_159.t0 93.987
R238 a_1150_159.n3 a_1150_159.n0 92.484
R239 a_1150_159.n3 a_1150_159.n2 9.323
R240 a_1500_413.t0 a_1500_413.t1 143.059
R241 a_1675_413.t0 a_1675_413.t1 197
R242 a_729_47.t0 a_729_47.t1 102.857
R243 a_729_369.t0 a_729_369.t1 110.812
R244 a_1077_413.t0 a_1077_413.t1 171.202
R245 a_1717_47.t1 a_1717_47.t0 93.059
R246 a_381_47.t0 a_381_47.t1 60
C0 VPWR Q 0.21fF
C1 VGND Q 0.15fF
C2 D DE 0.13fF
C3 VPWR VPB 0.24fF
C4 VPWR VGND 0.12fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__einvn_0.ext - technology: sky130A

.subckt sky130_fd_sc_hd__einvn_0 A TE_B Z VPWR VGND VNB VPB
X0 VGND.t0 TE_B.t0 a_30_47.t0 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1 Z.t0 A.t0 a_215_369.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X2 a_215_369.t1 TE_B.t1 VPWR.t0 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X3 a_215_47.t1 a_30_47.t2 VGND.t1 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 Z.t1 A.t1 a_215_47.t0 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 VPWR.t1 TE_B.t2 a_30_47.t1 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
R0 TE_B.n0 TE_B.t1 292.412
R1 TE_B.n1 TE_B.t0 206.188
R2 TE_B.n0 TE_B.t2 162.273
R3 TE_B.n1 TE_B.n0 124.248
R4 TE_B.n2 TE_B.n1 76
R5 TE_B.n2 TE_B 6.456
R6 TE_B TE_B.n2 1.246
R7 a_30_47.n0 a_30_47.t1 461.172
R8 a_30_47.n0 a_30_47.t2 278.808
R9 a_30_47.t0 a_30_47.n0 211.059
R10 VGND VGND.n0 96.798
R11 VGND.n0 VGND.t1 52.857
R12 VGND.n0 VGND.t0 51.428
R13 VNB VNB.t1 6567.65
R14 VNB.t1 VNB.t2 3332.35
R15 VNB.t2 VNB.t0 2329.41
R16 A.n0 A.t0 288.201
R17 A.n0 A.t1 195.015
R18 A.n1 A.n0 76
R19 A.n1 A 14.305
R20 A A.n1 2.76
R21 a_215_369.t0 a_215_369.t1 64.64
R22 Z Z.t0 335.748
R23 Z Z.t1 132.765
R24 VPB.t1 VPB.t2 304.828
R25 VPB.t2 VPB.t0 213.084
R26 VPB VPB.t1 201.246
R27 VPWR VPWR.n0 296.892
R28 VPWR.n0 VPWR.t1 86.773
R29 VPWR.n0 VPWR.t0 61.048
R30 a_215_47.t0 a_215_47.t1 60
C0 Z VGND 0.13fF
C1 VPWR Z 0.13fF
C2 A Z 0.30fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__einvn_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__einvn_1 Z A TE_B VGND VPWR VNB VPB
X0 VPWR.t1 TE_B.t0 a_27_47.t1 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1 a_204_297.t1 TE_B.t1 VPWR.t0 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 Z.t0 A.t0 a_204_297.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 Z.t1 A.t1 a_286_47.t1 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 a_286_47.t0 a_27_47.t2 VGND.t0 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 VGND.t1 TE_B.t2 a_27_47.t0 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
R0 TE_B.n0 TE_B.t1 313.299
R1 TE_B.n0 TE_B.t0 266.706
R2 TE_B.n1 TE_B.t2 229.753
R3 TE_B.n2 TE_B.n1 76
R4 TE_B.n1 TE_B.n0 56.233
R5 TE_B.n2 TE_B 8.583
R6 TE_B TE_B.n2 1.656
R7 a_27_47.t1 a_27_47.n0 398.946
R8 a_27_47.n0 a_27_47.t2 241.026
R9 a_27_47.n0 a_27_47.t0 173.936
R10 VPWR VPWR.n0 310.024
R11 VPWR.n0 VPWR.t1 49.25
R12 VPWR.n0 VPWR.t0 40.839
R13 VPB.t1 VPB.t0 523.831
R14 VPB.t2 VPB.t1 281.152
R15 VPB VPB.t2 192.367
R16 a_204_297.t0 a_204_297.t1 144.795
R17 A.n0 A.t0 230.361
R18 A.n0 A.t1 158.061
R19 A.n1 A.n0 76
R20 A.n1 A 14.889
R21 A A.n1 2.873
R22 Z Z.t0 173.974
R23 Z Z.t1 119.681
R24 Z.n0 Z 94.786
R25 Z.n0 Z 5.082
R26 Z Z.n0 3.576
R27 a_286_47.t0 a_286_47.t1 60
R28 VNB VNB.t1 6470.59
R29 VNB.t1 VNB.t0 4237.76
R30 VNB.t0 VNB.t2 2296.7
R31 VGND.n0 VGND.t1 67.138
R32 VGND.n0 VGND.t0 60.53
R33 VGND VGND.n0 37.326
C0 Z VGND 0.13fF
C1 VPWR Z 0.23fF
C2 A Z 0.25fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__einvn_2.ext - technology: sky130A

.subckt sky130_fd_sc_hd__einvn_2 TE_B A Z VPWR VGND VNB VPB
X0 Z.t3 A.t0 a_204_309.t1 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 VGND.t1 a_27_47.t2 a_214_120.t1 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 a_204_309.t0 A.t1 Z.t2 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 Z.t1 A.t2 a_214_120.t3 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 VPWR.t0 TE_B.t0 a_27_47.t0 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X5 VPWR.t2 TE_B.t1 a_204_309.t2 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=940000u l=150000u
X6 a_204_309.t3 TE_B.t2 VPWR.t1 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=940000u l=150000u
X7 a_214_120.t0 a_27_47.t3 VGND.t0 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 a_214_120.t2 A.t3 Z.t0 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 VGND.t2 TE_B.t3 a_27_47.t1 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
R0 A.n1 A.t0 234.037
R1 A.n0 A.t1 221.719
R2 A.n1 A.t3 161.737
R3 A.n0 A.t2 149.419
R4 A A.n1 78.011
R5 A.n1 A.n0 61.588
R6 a_204_309.n1 a_204_309.n0 511.94
R7 a_204_309.n0 a_204_309.t2 28.292
R8 a_204_309.n0 a_204_309.t3 28.292
R9 a_204_309.n1 a_204_309.t1 26.595
R10 a_204_309.t0 a_204_309.n1 26.595
R11 Z.n3 Z.t2 493.283
R12 Z.n1 Z.t3 208.131
R13 Z.n5 Z.n0 94.548
R14 Z.n0 Z.t0 24.923
R15 Z.n0 Z.t1 24.923
R16 Z Z.n4 17.408
R17 Z Z.n3 17.152
R18 Z.n4 Z.n2 15.104
R19 Z.n5 Z 13.312
R20 Z.n2 Z 7.862
R21 Z Z.n1 6.684
R22 Z.n3 Z 6.4
R23 Z.n1 Z 5.601
R24 Z.n2 Z 4.571
R25 Z Z.n5 4.096
R26 Z.n4 Z 2.304
R27 Z.n5 Z 2.304
R28 VPB.t3 VPB.t0 565.264
R29 VPB.t2 VPB.t4 281.152
R30 VPB.t0 VPB.t1 248.598
R31 VPB.t4 VPB.t3 248.598
R32 VPB VPB.t2 192.367
R33 a_27_47.t0 a_27_47.n1 387.354
R34 a_27_47.n0 a_27_47.t2 224.933
R35 a_27_47.n1 a_27_47.t1 170.828
R36 a_27_47.n1 a_27_47.n0 151.468
R37 a_27_47.n0 a_27_47.t3 147.071
R38 a_214_120.t2 a_214_120.n1 189.792
R39 a_214_120.n1 a_214_120.t1 181.546
R40 a_214_120.n1 a_214_120.n0 92.5
R41 a_214_120.n0 a_214_120.t0 32.307
R42 a_214_120.n0 a_214_120.t3 31.384
R43 VGND.n1 VGND.t2 150.43
R44 VGND.n1 VGND.n0 110.029
R45 VGND.n0 VGND.t0 24.923
R46 VGND.n0 VGND.t1 24.923
R47 VGND VGND.n1 0.218
R48 VNB VNB.t4 6470.59
R49 VNB.t4 VNB.t1 5289.53
R50 VNB.t0 VNB.t3 2393.41
R51 VNB.t3 VNB.t2 2030.77
R52 VNB.t1 VNB.t0 2030.77
R53 TE_B.n0 TE_B.t1 310.086
R54 TE_B.n1 TE_B.t0 247.426
R55 TE_B.n2 TE_B.t3 229.753
R56 TE_B.n0 TE_B.t2 175.126
R57 TE_B.n1 TE_B.n0 128.533
R58 TE_B TE_B.n2 101.756
R59 TE_B.n2 TE_B.n1 75.513
R60 VPWR.n1 VPWR.t2 491.965
R61 VPWR.n1 VPWR.n0 164.438
R62 VPWR.n0 VPWR.t0 49.25
R63 VPWR.n0 VPWR.t1 42.203
R64 VPWR VPWR.n1 0.236
C0 A Z 0.12fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__einvn_4.ext - technology: sky130A

.subckt sky130_fd_sc_hd__einvn_4 TE_B Z A VGND VPWR VNB VPB
X0 VGND.t3 a_27_47.t2 a_215_47.t7 VNB.t7 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 a_204_309.t7 A.t0 Z.t3 VPB.t8 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 VGND.t2 a_27_47.t3 a_215_47.t6 VNB.t6 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 VPWR.t4 TE_B.t0 a_204_309.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=940000u l=150000u
X4 Z.t7 A.t1 a_215_47.t0 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 a_204_309.t1 TE_B.t1 VPWR.t3 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=940000u l=150000u
X6 a_215_47.t5 a_27_47.t4 VGND.t1 VNB.t5 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 Z.t6 A.t2 a_215_47.t1 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 Z.t2 A.t3 a_204_309.t6 VPB.t7 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 VPWR.t2 TE_B.t2 a_204_309.t2 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=940000u l=150000u
X10 a_204_309.t3 TE_B.t3 VPWR.t1 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=940000u l=150000u
X11 a_215_47.t2 A.t4 Z.t5 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 a_215_47.t3 A.t5 Z.t4 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 a_215_47.t4 a_27_47.t5 VGND.t0 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14 a_204_309.t5 A.t6 Z.t1 VPB.t6 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 VPWR.t0 TE_B.t4 a_27_47.t0 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16 Z.t0 A.t7 a_204_309.t4 VPB.t5 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17 VGND.t4 TE_B.t5 a_27_47.t1 VNB.t8 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
R0 a_27_47.n0 a_27_47.t2 263.493
R1 a_27_47.t0 a_27_47.n3 249.016
R2 a_27_47.n3 a_27_47.n2 151.442
R3 a_27_47.n3 a_27_47.t1 148.974
R4 a_27_47.n1 a_27_47.n0 134.96
R5 a_27_47.n2 a_27_47.t4 134.475
R6 a_27_47.n0 a_27_47.t5 128.533
R7 a_27_47.n1 a_27_47.t3 128.533
R8 a_27_47.n2 a_27_47.n1 94.947
R9 a_215_47.n3 a_215_47.t3 231.209
R10 a_215_47.n1 a_215_47.t7 182.803
R11 a_215_47.n1 a_215_47.n0 99.652
R12 a_215_47.n3 a_215_47.n2 92.5
R13 a_215_47.n5 a_215_47.n4 92.5
R14 a_215_47.n4 a_215_47.n1 72.657
R15 a_215_47.n4 a_215_47.n3 65.061
R16 a_215_47.n5 a_215_47.t5 30.461
R17 a_215_47.t0 a_215_47.n5 29.538
R18 a_215_47.n0 a_215_47.t6 24.923
R19 a_215_47.n0 a_215_47.t4 24.923
R20 a_215_47.n2 a_215_47.t1 24.923
R21 a_215_47.n2 a_215_47.t2 24.923
R22 VGND.n6 VGND.t4 190.315
R23 VGND.n3 VGND.n0 109.922
R24 VGND.n2 VGND.n1 106.463
R25 VGND.n0 VGND.t1 24.923
R26 VGND.n0 VGND.t2 24.923
R27 VGND.n1 VGND.t0 24.923
R28 VGND.n1 VGND.t3 24.923
R29 VGND.n5 VGND.n4 4.65
R30 VGND.n7 VGND.n6 3.932
R31 VGND.n3 VGND.n2 3.796
R32 VGND.n5 VGND.n3 0.255
R33 VGND.n7 VGND.n5 0.137
R34 VGND VGND.n7 0.121
R35 VNB VNB.t8 6053.91
R36 VNB.t8 VNB.t7 4545.05
R37 VNB.t5 VNB.t0 2296.7
R38 VNB.t1 VNB.t3 2030.77
R39 VNB.t2 VNB.t1 2030.77
R40 VNB.t0 VNB.t2 2030.77
R41 VNB.t6 VNB.t5 2030.77
R42 VNB.t4 VNB.t6 2030.77
R43 VNB.t7 VNB.t4 2030.77
R44 A.n3 A.t6 212.079
R45 A.n2 A.t7 212.079
R46 A.n1 A.t0 212.079
R47 A.n0 A.t3 212.079
R48 A.n3 A.t5 139.779
R49 A.n2 A.t2 139.779
R50 A.n1 A.t4 139.779
R51 A.n0 A.t1 139.779
R52 A A.n3 138.197
R53 A.n3 A.n2 61.345
R54 A.n2 A.n1 61.345
R55 A.n1 A.n0 61.345
R56 Z.n2 Z.n0 154.517
R57 Z.n5 Z.n3 154.517
R58 Z.n5 Z.n4 92.5
R59 Z.n2 Z.n1 92.5
R60 Z.n0 Z.t1 26.595
R61 Z.n0 Z.t0 26.595
R62 Z.n3 Z.t3 26.595
R63 Z.n3 Z.t2 26.595
R64 Z.n1 Z.t4 24.923
R65 Z.n1 Z.t6 24.923
R66 Z.n4 Z.t5 24.923
R67 Z.n4 Z.t7 24.923
R68 Z Z.n2 5.432
R69 Z Z.n5 0.223
R70 a_204_309.t6 a_204_309.n2 421.307
R71 a_204_309.t6 a_204_309.n6 421.307
R72 a_204_309.n1 a_204_309.t5 276.389
R73 a_204_309.n5 a_204_309.n4 221.147
R74 a_204_309.n5 a_204_309.n3 163.677
R75 a_204_309.n1 a_204_309.n0 162.924
R76 a_204_309.n6 a_204_309.n5 75.687
R77 a_204_309.n2 a_204_309.n1 70.561
R78 a_204_309.n4 a_204_309.t2 28.292
R79 a_204_309.n4 a_204_309.t3 28.292
R80 a_204_309.n3 a_204_309.t0 28.292
R81 a_204_309.n3 a_204_309.t1 28.292
R82 a_204_309.n0 a_204_309.t4 26.595
R83 a_204_309.n0 a_204_309.t7 26.595
R84 VPB.t0 VPB.t7 556.386
R85 VPB.t4 VPB.t3 281.152
R86 VPB.t5 VPB.t6 248.598
R87 VPB.t8 VPB.t5 248.598
R88 VPB.t7 VPB.t8 248.598
R89 VPB.t1 VPB.t0 248.598
R90 VPB.t2 VPB.t1 248.598
R91 VPB.t3 VPB.t2 248.598
R92 VPB VPB.t4 189.408
R93 TE_B.n0 TE_B.t0 310.086
R94 TE_B.n3 TE_B.t4 220.389
R95 TE_B.n2 TE_B.t3 199.226
R96 TE_B.n0 TE_B.t1 175.126
R97 TE_B.n1 TE_B.t2 175.126
R98 TE_B.n4 TE_B.t5 158.061
R99 TE_B.n3 TE_B.n2 151.026
R100 TE_B.n1 TE_B.n0 134.96
R101 TE_B.n2 TE_B.n1 110.86
R102 TE_B TE_B.n4 79.684
R103 TE_B.n4 TE_B.n3 9.972
R104 VPWR.n2 VPWR.t4 193.09
R105 VPWR.n1 VPWR.n0 163.438
R106 VPWR.n6 VPWR.n5 163.438
R107 VPWR.n5 VPWR.t1 39.819
R108 VPWR.n0 VPWR.t3 28.292
R109 VPWR.n0 VPWR.t2 28.292
R110 VPWR.n5 VPWR.t0 26.451
R111 VPWR.n4 VPWR.n3 4.65
R112 VPWR.n7 VPWR.n6 3.932
R113 VPWR.n2 VPWR.n1 3.864
R114 VPWR.n4 VPWR.n2 0.257
R115 VPWR.n7 VPWR.n4 0.137
R116 VPWR VPWR.n7 0.121
C0 VGND VPWR 0.11fF
C1 Z A 0.15fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__einvn_8.ext - technology: sky130A

.subckt sky130_fd_sc_hd__einvn_8 A TE_B Z VGND VPWR VNB VPB
X0 a_204_309.t7 A.t0 Z.t0 VPB.t7 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 VGND.t7 a_27_47.t2 a_215_47.t15 VNB.t15 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 a_215_47.t7 A.t1 Z.t15 VNB.t7 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 Z.t8 A.t2 a_204_309.t6 VPB.t6 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 VGND.t6 a_27_47.t3 a_215_47.t14 VNB.t14 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 VGND.t5 a_27_47.t4 a_215_47.t13 VNB.t13 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 a_204_309.t8 TE_B.t0 VPWR.t8 VPB.t8 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=940000u l=150000u
X7 a_204_309.t5 A.t3 Z.t7 VPB.t5 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 VGND.t4 a_27_47.t5 a_215_47.t12 VNB.t12 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 VPWR.t7 TE_B.t1 a_204_309.t9 VPB.t9 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=940000u l=150000u
X10 Z.t6 A.t4 a_204_309.t4 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 a_204_309.t10 TE_B.t2 VPWR.t6 VPB.t10 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=940000u l=150000u
X12 a_215_47.t11 a_27_47.t6 VGND.t3 VNB.t11 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 Z.t14 A.t5 a_215_47.t6 VNB.t6 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14 a_215_47.t10 a_27_47.t7 VGND.t2 VNB.t10 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X15 a_215_47.t9 a_27_47.t8 VGND.t1 VNB.t9 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X16 VPWR.t5 TE_B.t3 a_204_309.t11 VPB.t11 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=940000u l=150000u
X17 a_215_47.t5 A.t6 Z.t13 VNB.t5 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X18 a_204_309.t12 TE_B.t4 VPWR.t4 VPB.t12 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=940000u l=150000u
X19 a_215_47.t4 A.t7 Z.t12 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X20 a_215_47.t3 A.t8 Z.t11 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X21 a_204_309.t3 A.t9 Z.t5 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X22 VPWR.t3 TE_B.t5 a_204_309.t13 VPB.t13 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=940000u l=150000u
X23 a_204_309.t14 TE_B.t6 VPWR.t2 VPB.t14 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=940000u l=150000u
X24 Z.t4 A.t10 a_204_309.t2 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X25 Z.t10 A.t11 a_215_47.t2 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X26 Z.t3 A.t12 a_204_309.t1 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X27 a_204_309.t0 A.t13 Z.t2 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X28 Z.t9 A.t14 a_215_47.t1 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X29 VPWR.t1 TE_B.t7 a_204_309.t15 VPB.t15 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=940000u l=150000u
X30 Z.t1 A.t15 a_215_47.t0 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X31 a_215_47.t8 a_27_47.t9 VGND.t0 VNB.t8 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X32 VPWR.t0 TE_B.t8 a_27_47.t0 VPB.t16 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X33 VGND.t8 TE_B.t9 a_27_47.t1 VNB.t16 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
R0 A.n1 A.t0 212.079
R1 A.n3 A.t2 212.079
R2 A.n0 A.t3 212.079
R3 A.n10 A.t4 212.079
R4 A.n13 A.t9 212.079
R5 A.n22 A.t10 212.079
R6 A.n15 A.t13 212.079
R7 A.n16 A.t12 212.079
R8 A.n1 A.t1 139.779
R9 A.n3 A.t15 139.779
R10 A.n0 A.t8 139.779
R11 A.n10 A.t14 139.779
R12 A.n13 A.t7 139.779
R13 A.n22 A.t11 139.779
R14 A.n15 A.t6 139.779
R15 A.n16 A.t5 139.779
R16 A.n2 A 81.517
R17 A.n6 A.n5 76
R18 A.n9 A.n8 76
R19 A.n12 A.n11 76
R20 A.n24 A.n23 76
R21 A.n21 A.n20 76
R22 A.n18 A.n17 76
R23 A.n5 A.n4 49.66
R24 A.n21 A.n14 49.66
R25 A.n17 A.n15 48.2
R26 A.n9 A.n0 45.278
R27 A.n3 A.n2 42.357
R28 A.n23 A.n22 39.436
R29 A.n11 A.n10 33.593
R30 A.n23 A.n13 21.909
R31 A.n2 A.n1 18.987
R32 A.n10 A.n9 16.066
R33 A.n8 A.n7 15.006
R34 A.n20 A.n19 15.006
R35 A.n12 A 13.903
R36 A.n17 A.n16 13.145
R37 A A.n18 13.02
R38 A.n24 A 11.696
R39 A A.n6 10.813
R40 A.n22 A.n21 10.224
R41 A.n6 A 9.489
R42 A A.n24 8.606
R43 A.n5 A.n3 7.303
R44 A.n18 A 7.282
R45 A A.n12 6.4
R46 A.n4 A.n0 4.381
R47 A.n7 A 4.193
R48 A.n20 A 3.31
R49 A.n19 A 1.986
R50 A.n15 A.n14 1.46
R51 A.n8 A 1.103
R52 Z.n2 Z.n0 194.081
R53 Z.n2 Z.n1 155.681
R54 Z.n15 Z.n14 147.863
R55 Z.n11 Z.n10 147.863
R56 Z.n7 Z.n6 144.948
R57 Z.n9 Z.n3 92.5
R58 Z.n8 Z.n4 92.5
R59 Z.n7 Z.n5 92.5
R60 Z.n9 Z.n8 52.448
R61 Z.n8 Z.n7 52.448
R62 Z.n12 Z 43.569
R63 Z.n13 Z.n2 38.4
R64 Z.n13 Z.n12 38.4
R65 Z Z.n9 28.472
R66 Z.n10 Z.t0 26.595
R67 Z.n10 Z.t8 26.595
R68 Z.n0 Z.t2 26.595
R69 Z.n0 Z.t3 26.595
R70 Z.n1 Z.t5 26.595
R71 Z.n1 Z.t4 26.595
R72 Z.n14 Z.t7 26.595
R73 Z.n14 Z.t6 26.595
R74 Z.n6 Z.t13 24.923
R75 Z.n6 Z.t14 24.923
R76 Z.n5 Z.t12 24.923
R77 Z.n5 Z.t10 24.923
R78 Z.n4 Z.t11 24.923
R79 Z.n4 Z.t9 24.923
R80 Z.n3 Z.t15 24.923
R81 Z.n3 Z.t1 24.923
R82 Z.n15 Z.n13 7.818
R83 Z.n12 Z.n11 7.818
R84 Z Z.n15 1.667
R85 Z.n11 Z 1.667
R86 a_204_309.t7 a_204_309.n13 236.531
R87 a_204_309.n7 a_204_309.n6 221.147
R88 a_204_309.n10 a_204_309.t1 206.39
R89 a_204_309.n9 a_204_309.n3 163.677
R90 a_204_309.n8 a_204_309.n4 163.677
R91 a_204_309.n7 a_204_309.n5 163.677
R92 a_204_309.n13 a_204_309.n0 152.295
R93 a_204_309.n12 a_204_309.n1 152.295
R94 a_204_309.n11 a_204_309.n2 152.295
R95 a_204_309.n10 a_204_309.n9 78.912
R96 a_204_309.n11 a_204_309.n10 76.895
R97 a_204_309.n9 a_204_309.n8 63.247
R98 a_204_309.n8 a_204_309.n7 63.247
R99 a_204_309.n13 a_204_309.n12 63.247
R100 a_204_309.n12 a_204_309.n11 63.247
R101 a_204_309.n6 a_204_309.t11 28.292
R102 a_204_309.n6 a_204_309.t12 28.292
R103 a_204_309.n3 a_204_309.t13 28.292
R104 a_204_309.n3 a_204_309.t14 28.292
R105 a_204_309.n4 a_204_309.t15 28.292
R106 a_204_309.n4 a_204_309.t8 28.292
R107 a_204_309.n5 a_204_309.t9 28.292
R108 a_204_309.n5 a_204_309.t10 28.292
R109 a_204_309.n2 a_204_309.t2 26.595
R110 a_204_309.n2 a_204_309.t0 26.595
R111 a_204_309.n1 a_204_309.t4 26.595
R112 a_204_309.n1 a_204_309.t3 26.595
R113 a_204_309.n0 a_204_309.t6 26.595
R114 a_204_309.n0 a_204_309.t5 26.595
R115 VPB.t13 VPB.t1 556.386
R116 VPB.t16 VPB.t12 281.152
R117 VPB.t6 VPB.t7 248.598
R118 VPB.t5 VPB.t6 248.598
R119 VPB.t4 VPB.t5 248.598
R120 VPB.t3 VPB.t4 248.598
R121 VPB.t2 VPB.t3 248.598
R122 VPB.t0 VPB.t2 248.598
R123 VPB.t1 VPB.t0 248.598
R124 VPB.t14 VPB.t13 248.598
R125 VPB.t15 VPB.t14 248.598
R126 VPB.t8 VPB.t15 248.598
R127 VPB.t9 VPB.t8 248.598
R128 VPB.t10 VPB.t9 248.598
R129 VPB.t11 VPB.t10 248.598
R130 VPB.t12 VPB.t11 248.598
R131 VPB VPB.t16 189.408
R132 a_27_47.n0 a_27_47.t2 263.493
R133 a_27_47.t0 a_27_47.n7 249.322
R134 a_27_47.n7 a_27_47.n6 216.606
R135 a_27_47.n7 a_27_47.t1 149.148
R136 a_27_47.n5 a_27_47.n4 134.96
R137 a_27_47.n4 a_27_47.n3 134.96
R138 a_27_47.n3 a_27_47.n2 134.96
R139 a_27_47.n2 a_27_47.n1 134.96
R140 a_27_47.n1 a_27_47.n0 134.96
R141 a_27_47.n6 a_27_47.t8 134.475
R142 a_27_47.n0 a_27_47.t9 128.533
R143 a_27_47.n1 a_27_47.t3 128.533
R144 a_27_47.n2 a_27_47.t6 128.533
R145 a_27_47.n3 a_27_47.t4 128.533
R146 a_27_47.n4 a_27_47.t7 128.533
R147 a_27_47.n5 a_27_47.t5 128.533
R148 a_27_47.n6 a_27_47.n5 94.947
R149 a_215_47.t7 a_215_47.n13 231.209
R150 a_215_47.n6 a_215_47.t15 182.803
R151 a_215_47.n6 a_215_47.n5 99.652
R152 a_215_47.n7 a_215_47.n4 99.652
R153 a_215_47.n8 a_215_47.n3 99.652
R154 a_215_47.n10 a_215_47.n9 92.5
R155 a_215_47.n13 a_215_47.n0 92.5
R156 a_215_47.n12 a_215_47.n1 92.5
R157 a_215_47.n11 a_215_47.n2 92.5
R158 a_215_47.n10 a_215_47.n8 68.316
R159 a_215_47.n8 a_215_47.n7 63.247
R160 a_215_47.n7 a_215_47.n6 63.247
R161 a_215_47.n11 a_215_47.n10 62.06
R162 a_215_47.n13 a_215_47.n12 55.138
R163 a_215_47.n12 a_215_47.n11 55.138
R164 a_215_47.n9 a_215_47.t9 30.461
R165 a_215_47.n9 a_215_47.t6 29.538
R166 a_215_47.n2 a_215_47.t2 24.923
R167 a_215_47.n2 a_215_47.t5 24.923
R168 a_215_47.n1 a_215_47.t1 24.923
R169 a_215_47.n1 a_215_47.t4 24.923
R170 a_215_47.n0 a_215_47.t0 24.923
R171 a_215_47.n0 a_215_47.t3 24.923
R172 a_215_47.n5 a_215_47.t14 24.923
R173 a_215_47.n5 a_215_47.t8 24.923
R174 a_215_47.n4 a_215_47.t13 24.923
R175 a_215_47.n4 a_215_47.t11 24.923
R176 a_215_47.n3 a_215_47.t12 24.923
R177 a_215_47.n3 a_215_47.t10 24.923
R178 VGND.n16 VGND.t8 190.315
R179 VGND.n3 VGND.n2 110.262
R180 VGND.n1 VGND.n0 106.463
R181 VGND.n7 VGND.n6 106.463
R182 VGND.n12 VGND.n11 106.463
R183 VGND.n2 VGND.t1 24.923
R184 VGND.n2 VGND.t4 24.923
R185 VGND.n0 VGND.t2 24.923
R186 VGND.n0 VGND.t5 24.923
R187 VGND.n6 VGND.t3 24.923
R188 VGND.n6 VGND.t6 24.923
R189 VGND.n11 VGND.t0 24.923
R190 VGND.n11 VGND.t7 24.923
R191 VGND.n5 VGND.n4 4.65
R192 VGND.n8 VGND.n7 4.65
R193 VGND.n10 VGND.n9 4.65
R194 VGND.n13 VGND.n12 4.65
R195 VGND.n15 VGND.n14 4.65
R196 VGND.n17 VGND.n16 3.932
R197 VGND.n3 VGND.n1 3.876
R198 VGND.n5 VGND.n3 0.376
R199 VGND.n17 VGND.n15 0.137
R200 VGND VGND.n17 0.121
R201 VGND.n8 VGND.n5 0.119
R202 VGND.n10 VGND.n8 0.119
R203 VGND.n13 VGND.n10 0.119
R204 VGND.n15 VGND.n13 0.119
R205 VNB VNB.t16 6053.91
R206 VNB.t16 VNB.t15 4545.05
R207 VNB.t9 VNB.t6 2296.7
R208 VNB.t0 VNB.t7 2030.77
R209 VNB.t3 VNB.t0 2030.77
R210 VNB.t1 VNB.t3 2030.77
R211 VNB.t4 VNB.t1 2030.77
R212 VNB.t2 VNB.t4 2030.77
R213 VNB.t5 VNB.t2 2030.77
R214 VNB.t6 VNB.t5 2030.77
R215 VNB.t12 VNB.t9 2030.77
R216 VNB.t10 VNB.t12 2030.77
R217 VNB.t13 VNB.t10 2030.77
R218 VNB.t11 VNB.t13 2030.77
R219 VNB.t14 VNB.t11 2030.77
R220 VNB.t8 VNB.t14 2030.77
R221 VNB.t15 VNB.t8 2030.77
R222 TE_B.n0 TE_B.t5 310.086
R223 TE_B.n7 TE_B.t8 220.389
R224 TE_B.n6 TE_B.t4 199.226
R225 TE_B.n0 TE_B.t6 175.126
R226 TE_B.n1 TE_B.t7 175.126
R227 TE_B.n2 TE_B.t0 175.126
R228 TE_B.n3 TE_B.t1 175.126
R229 TE_B.n4 TE_B.t2 175.126
R230 TE_B.n5 TE_B.t3 175.126
R231 TE_B.n8 TE_B.t9 158.061
R232 TE_B.n7 TE_B.n6 151.026
R233 TE_B.n1 TE_B.n0 134.96
R234 TE_B.n2 TE_B.n1 134.96
R235 TE_B.n3 TE_B.n2 134.96
R236 TE_B.n4 TE_B.n3 134.96
R237 TE_B.n5 TE_B.n4 134.96
R238 TE_B.n6 TE_B.n5 110.86
R239 TE_B TE_B.n8 79.684
R240 TE_B.n8 TE_B.n7 9.972
R241 VPWR.n2 VPWR.t3 194.996
R242 VPWR.n1 VPWR.n0 163.438
R243 VPWR.n6 VPWR.n5 163.438
R244 VPWR.n11 VPWR.n10 163.438
R245 VPWR.n16 VPWR.n15 163.438
R246 VPWR.n15 VPWR.t4 39.819
R247 VPWR.n0 VPWR.t2 28.292
R248 VPWR.n0 VPWR.t1 28.292
R249 VPWR.n5 VPWR.t8 28.292
R250 VPWR.n5 VPWR.t7 28.292
R251 VPWR.n10 VPWR.t6 28.292
R252 VPWR.n10 VPWR.t5 28.292
R253 VPWR.n15 VPWR.t0 26.451
R254 VPWR.n2 VPWR.n1 6.066
R255 VPWR.n4 VPWR.n3 4.65
R256 VPWR.n7 VPWR.n6 4.65
R257 VPWR.n9 VPWR.n8 4.65
R258 VPWR.n12 VPWR.n11 4.65
R259 VPWR.n14 VPWR.n13 4.65
R260 VPWR.n17 VPWR.n16 3.932
R261 VPWR.n4 VPWR.n2 0.457
R262 VPWR.n17 VPWR.n14 0.137
R263 VPWR VPWR.n17 0.121
R264 VPWR.n7 VPWR.n4 0.119
R265 VPWR.n9 VPWR.n7 0.119
R266 VPWR.n12 VPWR.n9 0.119
R267 VPWR.n14 VPWR.n12 0.119
C0 VPB A 0.11fF
C1 A Z 1.08fF
C2 VPB VPWR 0.16fF
C3 VPWR VGND 0.17fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__einvp_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__einvp_1 TE A Z VPWR VGND VNB VPB
X0 a_276_297.t1 a_27_47.t2 VPWR.t1 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 Z.t1 A.t0 a_204_47.t1 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 VPWR.t0 TE.t0 a_27_47.t0 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3 Z.t0 A.t1 a_276_297.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 a_204_47.t0 TE.t1 VGND.t1 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 VGND.t0 TE.t2 a_27_47.t1 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
R0 a_27_47.t0 a_27_47.n0 412.482
R1 a_27_47.n0 a_27_47.t2 317.534
R2 a_27_47.n0 a_27_47.t1 180.766
R3 VPWR VPWR.n0 174.791
R4 VPWR.n0 VPWR.t1 93.655
R5 VPWR.n0 VPWR.t0 35.178
R6 a_276_297.t0 a_276_297.t1 71.905
R7 VPB.t1 VPB.t2 494.236
R8 VPB.t2 VPB.t0 304.828
R9 VPB VPB.t1 189.408
R10 A.n0 A.t1 229.752
R11 A.n0 A.t0 157.452
R12 A.n1 A.n0 76
R13 A.n1 A 15.2
R14 A A.n1 2.933
R15 a_204_47.t0 a_204_47.t1 133.846
R16 Z Z.t0 524.215
R17 Z.n0 Z 112.129
R18 Z.n0 Z.t1 82.642
R19 Z Z.n0 3.206
R20 VNB VNB.t1 6438.23
R21 VNB.t0 VNB.t2 4230.77
R22 VNB.t1 VNB.t0 2255.35
R23 TE.n1 TE.t0 358.286
R24 TE.n0 TE.t1 257.066
R25 TE.n0 TE.t2 189.586
R26 TE.n2 TE.n1 95.944
R27 TE.n1 TE.n0 40.166
R28 TE.n2 TE 7.93
R29 TE TE.n2 1.53
R30 VGND VGND.n0 95.934
R31 VGND.n0 VGND.t1 41.648
R32 VGND.n0 VGND.t0 38.571
C0 Z VGND 0.14fF
C1 VPWR Z 0.13fF
C2 A Z 0.26fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__einvp_2.ext - technology: sky130A

.subckt sky130_fd_sc_hd__einvp_2 A Z TE VGND VPWR VNB VPB
X0 VPWR.t2 a_27_47.t2 a_215_309.t3 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=940000u l=150000u
X1 a_204_47.t2 A.t0 Z.t3 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 VPWR.t0 TE.t0 a_27_47.t0 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X3 Z.t2 A.t1 a_204_47.t1 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 a_215_309.t0 A.t2 Z.t1 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 Z.t0 A.t3 a_215_309.t1 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 a_204_47.t0 TE.t1 VGND.t2 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 VGND.t1 TE.t2 a_204_47.t3 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 a_215_309.t2 a_27_47.t3 VPWR.t1 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=940000u l=150000u
X9 VGND.t0 TE.t3 a_27_47.t1 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
R0 a_27_47.t0 a_27_47.n1 384.481
R1 a_27_47.n0 a_27_47.t2 253.852
R2 a_27_47.n0 a_27_47.t3 189.586
R3 a_27_47.n1 a_27_47.t1 171.6
R4 a_27_47.n1 a_27_47.n0 156.798
R5 a_215_309.n1 a_215_309.t3 284.896
R6 a_215_309.t0 a_215_309.n1 250.977
R7 a_215_309.n1 a_215_309.n0 140.206
R8 a_215_309.n0 a_215_309.t2 34.579
R9 a_215_309.n0 a_215_309.t1 31.691
R10 VPWR.n1 VPWR.t0 441.901
R11 VPWR.n1 VPWR.n0 166.996
R12 VPWR.n0 VPWR.t1 28.292
R13 VPWR.n0 VPWR.t2 28.292
R14 VPWR VPWR.n1 0.222
R15 VPB.t2 VPB.t4 556.386
R16 VPB.t3 VPB.t1 281.152
R17 VPB.t1 VPB.t0 248.598
R18 VPB.t4 VPB.t3 248.598
R19 VPB VPB.t2 189.408
R20 A.n1 A.t2 212.079
R21 A.n0 A.t3 212.079
R22 A.n1 A.t0 139.779
R23 A.n0 A.t1 139.779
R24 A.n2 A.n1 113.245
R25 A.n1 A.n0 61.345
R26 A.n2 A 12.8
R27 A A.n2 2.47
R28 Z.n2 Z.n1 146.156
R29 Z Z.n0 92.693
R30 Z.n1 Z.t1 26.595
R31 Z.n1 Z.t0 26.595
R32 Z.n0 Z.t3 24.923
R33 Z.n0 Z.t2 24.923
R34 Z.n2 Z 9.719
R35 Z Z.n2 3.392
R36 a_204_47.t2 a_204_47.n1 221.162
R37 a_204_47.n1 a_204_47.n0 169.594
R38 a_204_47.n1 a_204_47.t1 117.423
R39 a_204_47.n0 a_204_47.t3 24.923
R40 a_204_47.n0 a_204_47.t0 24.923
R41 VNB VNB.t4 6438.23
R42 VNB.t3 VNB.t1 4545.05
R43 VNB.t4 VNB.t0 2255.35
R44 VNB.t1 VNB.t2 2030.77
R45 VNB.t0 VNB.t3 2030.77
R46 TE.n2 TE.t0 322.939
R47 TE.n0 TE.t2 263.493
R48 TE.n1 TE.t3 189.586
R49 TE.n0 TE.t1 128.533
R50 TE.n1 TE.n0 128.533
R51 TE.n3 TE.n2 97.909
R52 TE.n2 TE.n1 40.166
R53 TE.n3 TE 14.889
R54 TE TE.n3 2.873
R55 VGND.n1 VGND.t1 192.59
R56 VGND.n1 VGND.n0 96.248
R57 VGND.n0 VGND.t0 47.142
R58 VGND.n0 VGND.t2 33.077
R59 VGND VGND.n1 0.233
C0 A Z 0.13fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__einvp_4.ext - technology: sky130A

.subckt sky130_fd_sc_hd__einvp_4 TE A Z VPWR VGND VNB VPB
X0 VPWR.t4 a_27_47.t2 a_215_309.t3 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=940000u l=150000u
X1 a_215_309.t4 A.t0 Z.t7 VPB.t5 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 VGND.t4 TE.t0 a_193_47.t3 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 Z.t3 A.t1 a_193_47.t7 VNB.t8 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 Z.t2 A.t2 a_193_47.t6 VNB.t7 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 a_193_47.t2 TE.t1 VGND.t3 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 Z.t6 A.t3 a_215_309.t5 VPB.t6 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 a_193_47.t1 TE.t2 VGND.t2 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 a_193_47.t5 A.t4 Z.t1 VNB.t6 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 a_193_47.t4 A.t5 Z.t0 VNB.t5 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 VGND.t1 TE.t3 a_193_47.t0 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 a_215_309.t2 a_27_47.t3 VPWR.t3 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=940000u l=150000u
X12 VPWR.t2 a_27_47.t4 a_215_309.t1 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=940000u l=150000u
X13 a_215_309.t0 a_27_47.t5 VPWR.t1 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=940000u l=150000u
X14 a_215_309.t6 A.t6 Z.t5 VPB.t7 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 VPWR.t0 TE.t4 a_27_47.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16 Z.t4 A.t7 a_215_309.t7 VPB.t8 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17 VGND.t0 TE.t5 a_27_47.t1 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
R0 a_27_47.t0 a_27_47.n3 479.311
R1 a_27_47.n0 a_27_47.t2 310.086
R2 a_27_47.n2 a_27_47.t3 188.514
R3 a_27_47.n3 a_27_47.n2 185.247
R4 a_27_47.n1 a_27_47.t4 175.126
R5 a_27_47.n0 a_27_47.t5 175.126
R6 a_27_47.n3 a_27_47.t1 165.986
R7 a_27_47.n1 a_27_47.n0 134.96
R8 a_27_47.n2 a_27_47.n1 72.3
R9 a_215_309.n2 a_215_309.t3 556.398
R10 a_215_309.n4 a_215_309.t6 234.399
R11 a_215_309.n2 a_215_309.n1 170.077
R12 a_215_309.n5 a_215_309.n4 152.296
R13 a_215_309.n3 a_215_309.n0 140.206
R14 a_215_309.n3 a_215_309.n2 95.29
R15 a_215_309.n4 a_215_309.n3 77.22
R16 a_215_309.n0 a_215_309.t2 34.579
R17 a_215_309.n0 a_215_309.t5 31.691
R18 a_215_309.n1 a_215_309.t1 28.292
R19 a_215_309.n1 a_215_309.t0 28.292
R20 a_215_309.n5 a_215_309.t7 26.595
R21 a_215_309.t4 a_215_309.n5 26.595
R22 VPWR.n6 VPWR.t0 574.991
R23 VPWR.n3 VPWR.n2 165.445
R24 VPWR.n1 VPWR.n0 163.438
R25 VPWR.n2 VPWR.t3 28.292
R26 VPWR.n2 VPWR.t2 28.292
R27 VPWR.n0 VPWR.t1 28.292
R28 VPWR.n0 VPWR.t4 28.292
R29 VPWR.n5 VPWR.n4 4.65
R30 VPWR.n7 VPWR.n6 3.932
R31 VPWR.n3 VPWR.n1 3.796
R32 VPWR.n5 VPWR.n3 0.254
R33 VPWR.n7 VPWR.n5 0.137
R34 VPWR VPWR.n7 0.121
R35 VPB.t0 VPB.t4 556.386
R36 VPB.t3 VPB.t6 281.152
R37 VPB.t8 VPB.t7 248.598
R38 VPB.t5 VPB.t8 248.598
R39 VPB.t6 VPB.t5 248.598
R40 VPB.t2 VPB.t3 248.598
R41 VPB.t1 VPB.t2 248.598
R42 VPB.t4 VPB.t1 248.598
R43 VPB VPB.t0 189.408
R44 A.n1 A.t6 235.146
R45 A.n4 A.t7 221.719
R46 A.n6 A.t0 212.079
R47 A.n5 A.t3 212.079
R48 A.n1 A.t5 162.846
R49 A.n4 A.t2 149.419
R50 A.n6 A.t4 139.779
R51 A.n5 A.t1 139.779
R52 A.n1 A.n0 76
R53 A.n3 A.n2 76
R54 A.n8 A.n7 76
R55 A.n6 A.n5 61.345
R56 A.n7 A.n6 58.261
R57 A.n8 A.n3 17.066
R58 A.n2 A.n1 15.174
R59 A.n7 A.n4 14.281
R60 A.n0 A 13.803
R61 A.n0 A 9.286
R62 A.n3 A 3.262
R63 A A.n8 2.76
R64 Z Z.n1 166.13
R65 Z.n2 Z.n0 152.163
R66 Z.n5 Z.n4 130.382
R67 Z.n5 Z.n3 92.5
R68 Z.n0 Z.t7 26.595
R69 Z.n0 Z.t6 26.595
R70 Z.n1 Z.t5 26.595
R71 Z.n1 Z.t4 26.595
R72 Z.n3 Z.t1 24.923
R73 Z.n3 Z.t3 24.923
R74 Z.n4 Z.t0 24.923
R75 Z.n4 Z.t2 24.923
R76 Z.n2 Z 21.082
R77 Z Z.n2 2.863
R78 Z Z.n5 0.168
R79 TE.n4 TE.t4 265.099
R80 TE.n0 TE.t3 263.493
R81 TE.n3 TE.t5 152.633
R82 TE.n2 TE.n1 141.386
R83 TE.n1 TE.n0 134.96
R84 TE.n2 TE.t2 128.533
R85 TE.n1 TE.t0 128.533
R86 TE.n0 TE.t1 128.533
R87 TE.n3 TE.n2 110.86
R88 TE.n5 TE.n4 97.909
R89 TE.n4 TE.n3 40.166
R90 TE.n5 TE 14.889
R91 TE TE.n5 2.873
R92 a_193_47.n4 a_193_47.t4 229.414
R93 a_193_47.n2 a_193_47.n1 164.782
R94 a_193_47.n3 a_193_47.t7 117.423
R95 a_193_47.n2 a_193_47.n0 101.535
R96 a_193_47.n5 a_193_47.n4 92.5
R97 a_193_47.n3 a_193_47.n2 67.559
R98 a_193_47.n4 a_193_47.n3 53.878
R99 a_193_47.n1 a_193_47.t1 28.615
R100 a_193_47.n1 a_193_47.t3 24.923
R101 a_193_47.n0 a_193_47.t0 24.923
R102 a_193_47.n0 a_193_47.t2 24.923
R103 a_193_47.t6 a_193_47.n5 24.923
R104 a_193_47.n5 a_193_47.t5 24.923
R105 VGND.n2 VGND.t1 195.046
R106 VGND.n1 VGND.n0 106.463
R107 VGND.n6 VGND.n5 106.463
R108 VGND.n0 VGND.t3 24.923
R109 VGND.n0 VGND.t4 24.923
R110 VGND.n5 VGND.t2 24.923
R111 VGND.n5 VGND.t0 24.923
R112 VGND.n4 VGND.n3 4.65
R113 VGND.n7 VGND.n6 3.932
R114 VGND.n2 VGND.n1 3.902
R115 VGND.n4 VGND.n2 0.265
R116 VGND.n7 VGND.n4 0.137
R117 VGND VGND.n7 0.121
R118 VNB VNB.t0 6053.91
R119 VNB.t1 VNB.t8 4714.29
R120 VNB.t2 VNB.t4 2127.47
R121 VNB.t7 VNB.t5 2030.77
R122 VNB.t6 VNB.t7 2030.77
R123 VNB.t8 VNB.t6 2030.77
R124 VNB.t3 VNB.t1 2030.77
R125 VNB.t4 VNB.t3 2030.77
R126 VNB.t0 VNB.t2 2030.77
C0 VPWR VGND 0.11fF
C1 A Z 0.40fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__einvp_8.ext - technology: sky130A

.subckt sky130_fd_sc_hd__einvp_8 A Z TE VPWR VGND VNB VPB
X0 VPWR.t8 a_27_47.t2 a_215_309.t13 VPB.t14 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=940000u l=150000u
X1 a_215_309.t0 A.t0 Z.t8 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 a_193_47.t15 A.t1 Z.t15 VNB.t16 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 a_215_309.t12 a_27_47.t3 VPWR.t7 VPB.t13 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=940000u l=150000u
X4 Z.t7 A.t2 a_215_309.t1 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 VGND.t7 TE.t0 a_193_47.t0 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 a_215_309.t2 A.t3 Z.t6 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 VPWR.t6 a_27_47.t4 a_215_309.t11 VPB.t12 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=940000u l=150000u
X8 a_215_309.t10 a_27_47.t5 VPWR.t5 VPB.t11 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=940000u l=150000u
X9 Z.t5 A.t4 a_215_309.t3 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 a_193_47.t1 TE.t1 VGND.t6 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 Z.t14 A.t5 a_193_47.t14 VNB.t15 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 a_193_47.t2 TE.t2 VGND.t5 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 a_193_47.t3 TE.t3 VGND.t4 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14 a_193_47.t4 TE.t4 VGND.t3 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X15 a_193_47.t13 A.t6 Z.t13 VNB.t14 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X16 a_193_47.t12 A.t7 Z.t12 VNB.t13 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X17 a_193_47.t11 A.t8 Z.t11 VNB.t12 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X18 a_215_309.t4 A.t9 Z.t4 VPB.t5 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X19 VGND.t2 TE.t5 a_193_47.t5 VNB.t5 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X20 VPWR.t4 a_27_47.t6 a_215_309.t9 VPB.t10 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=940000u l=150000u
X21 VGND.t1 TE.t6 a_193_47.t6 VNB.t6 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X22 VGND.t0 TE.t7 a_193_47.t7 VNB.t7 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X23 Z.t3 A.t10 a_215_309.t5 VPB.t6 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X24 Z.t10 A.t11 a_193_47.t10 VNB.t11 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X25 a_215_309.t8 a_27_47.t7 VPWR.t3 VPB.t9 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=940000u l=150000u
X26 Z.t2 A.t12 a_215_309.t14 VPB.t15 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X27 a_215_309.t15 A.t13 Z.t1 VPB.t16 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X28 Z.t9 A.t14 a_193_47.t9 VNB.t10 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X29 VPWR.t2 a_27_47.t8 a_215_309.t7 VPB.t8 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=940000u l=150000u
X30 Z.t0 A.t15 a_193_47.t8 VNB.t9 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X31 a_215_309.t6 a_27_47.t9 VPWR.t1 VPB.t7 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=940000u l=150000u
X32 VPWR.t0 TE.t8 a_27_47.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X33 VGND.t8 TE.t9 a_27_47.t1 VNB.t8 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
R0 a_27_47.t0 a_27_47.n7 479.311
R1 a_27_47.n0 a_27_47.t2 310.086
R2 a_27_47.n7 a_27_47.n6 250.411
R3 a_27_47.n6 a_27_47.t3 188.514
R4 a_27_47.n5 a_27_47.t4 175.126
R5 a_27_47.n4 a_27_47.t5 175.126
R6 a_27_47.n3 a_27_47.t6 175.126
R7 a_27_47.n2 a_27_47.t7 175.126
R8 a_27_47.n1 a_27_47.t8 175.126
R9 a_27_47.n0 a_27_47.t9 175.126
R10 a_27_47.n7 a_27_47.t1 165.986
R11 a_27_47.n5 a_27_47.n4 134.96
R12 a_27_47.n4 a_27_47.n3 134.96
R13 a_27_47.n3 a_27_47.n2 134.96
R14 a_27_47.n2 a_27_47.n1 134.96
R15 a_27_47.n1 a_27_47.n0 134.96
R16 a_27_47.n6 a_27_47.n5 72.3
R17 a_215_309.n6 a_215_309.t13 556.398
R18 a_215_309.t0 a_215_309.n13 236.533
R19 a_215_309.n8 a_215_309.n3 170.077
R20 a_215_309.n7 a_215_309.n4 170.077
R21 a_215_309.n6 a_215_309.n5 170.077
R22 a_215_309.n11 a_215_309.n2 152.295
R23 a_215_309.n12 a_215_309.n1 152.295
R24 a_215_309.n13 a_215_309.n0 152.295
R25 a_215_309.n10 a_215_309.n9 141.57
R26 a_215_309.n10 a_215_309.n8 84.413
R27 a_215_309.n11 a_215_309.n10 70.76
R28 a_215_309.n8 a_215_309.n7 63.247
R29 a_215_309.n7 a_215_309.n6 63.247
R30 a_215_309.n13 a_215_309.n12 63.247
R31 a_215_309.n12 a_215_309.n11 63.247
R32 a_215_309.n9 a_215_309.t12 34.579
R33 a_215_309.n9 a_215_309.t14 31.691
R34 a_215_309.n3 a_215_309.t11 28.292
R35 a_215_309.n3 a_215_309.t10 28.292
R36 a_215_309.n4 a_215_309.t9 28.292
R37 a_215_309.n4 a_215_309.t8 28.292
R38 a_215_309.n5 a_215_309.t7 28.292
R39 a_215_309.n5 a_215_309.t6 28.292
R40 a_215_309.n0 a_215_309.t1 26.595
R41 a_215_309.n0 a_215_309.t2 26.595
R42 a_215_309.n1 a_215_309.t3 26.595
R43 a_215_309.n1 a_215_309.t4 26.595
R44 a_215_309.n2 a_215_309.t5 26.595
R45 a_215_309.n2 a_215_309.t15 26.595
R46 VPWR.n16 VPWR.t0 574.991
R47 VPWR.n3 VPWR.n2 167.831
R48 VPWR.n1 VPWR.n0 163.438
R49 VPWR.n7 VPWR.n6 163.438
R50 VPWR.n12 VPWR.n11 163.438
R51 VPWR.n2 VPWR.t7 28.292
R52 VPWR.n2 VPWR.t6 28.292
R53 VPWR.n0 VPWR.t5 28.292
R54 VPWR.n0 VPWR.t4 28.292
R55 VPWR.n6 VPWR.t3 28.292
R56 VPWR.n6 VPWR.t2 28.292
R57 VPWR.n11 VPWR.t1 28.292
R58 VPWR.n11 VPWR.t8 28.292
R59 VPWR.n5 VPWR.n4 4.65
R60 VPWR.n8 VPWR.n7 4.65
R61 VPWR.n10 VPWR.n9 4.65
R62 VPWR.n13 VPWR.n12 4.65
R63 VPWR.n15 VPWR.n14 4.65
R64 VPWR.n17 VPWR.n16 3.932
R65 VPWR.n3 VPWR.n1 3.866
R66 VPWR.n5 VPWR.n3 0.386
R67 VPWR.n17 VPWR.n15 0.137
R68 VPWR VPWR.n17 0.121
R69 VPWR.n8 VPWR.n5 0.119
R70 VPWR.n10 VPWR.n8 0.119
R71 VPWR.n13 VPWR.n10 0.119
R72 VPWR.n15 VPWR.n13 0.119
R73 VPB.t0 VPB.t14 556.386
R74 VPB.t13 VPB.t15 281.152
R75 VPB.t2 VPB.t1 248.598
R76 VPB.t3 VPB.t2 248.598
R77 VPB.t4 VPB.t3 248.598
R78 VPB.t5 VPB.t4 248.598
R79 VPB.t6 VPB.t5 248.598
R80 VPB.t16 VPB.t6 248.598
R81 VPB.t15 VPB.t16 248.598
R82 VPB.t12 VPB.t13 248.598
R83 VPB.t11 VPB.t12 248.598
R84 VPB.t10 VPB.t11 248.598
R85 VPB.t9 VPB.t10 248.598
R86 VPB.t8 VPB.t9 248.598
R87 VPB.t7 VPB.t8 248.598
R88 VPB.t14 VPB.t7 248.598
R89 VPB VPB.t0 189.408
R90 A.n1 A.t0 234.39
R91 A.n9 A.t9 221.719
R92 A.n13 A.t10 221.719
R93 A.n4 A.t2 221.719
R94 A.n11 A.t13 212.079
R95 A.n10 A.t12 212.079
R96 A.n19 A.t3 212.079
R97 A.n7 A.t4 212.079
R98 A.n1 A.t1 162.09
R99 A.n9 A.t7 149.419
R100 A.n13 A.t11 149.419
R101 A.n4 A.t15 149.419
R102 A.n11 A.t6 139.779
R103 A.n10 A.t5 139.779
R104 A.n19 A.t8 139.779
R105 A.n7 A.t14 139.779
R106 A.n12 A 81.27
R107 A.n1 A.n0 76
R108 A.n3 A.n2 76
R109 A.n6 A.n5 76
R110 A.n21 A.n20 76
R111 A.n18 A.n17 76
R112 A.n15 A.n14 76
R113 A.n11 A.n10 61.345
R114 A.n12 A.n11 58.261
R115 A.n4 A.n3 49.985
R116 A.n19 A.n18 46.739
R117 A.n14 A.n13 46.414
R118 A.n8 A.n7 40.409
R119 A.n9 A.n8 32.133
R120 A.n14 A.n9 28.562
R121 A.n17 A.n16 17.066
R122 A.n21 A 16.815
R123 A.n18 A.n7 14.606
R124 A.n13 A.n12 14.281
R125 A.n6 A 12.298
R126 A.n15 A 11.796
R127 A.n3 A.n1 11.603
R128 A A.n15 11.294
R129 A A.n6 10.792
R130 A.n5 A.n4 10.711
R131 A A.n21 6.274
R132 A.n16 A 5.772
R133 A.n2 A 4.768
R134 A.n20 A.n19 2.921
R135 A.n0 A 1.254
R136 A.n17 A 0.25
R137 Z.n10 Z.n9 152.578
R138 Z.n8 Z.n0 152.163
R139 Z.n12 Z.n11 146.156
R140 Z.n15 Z.n14 146.156
R141 Z.n4 Z.n2 142.509
R142 Z.n6 Z.n5 92.5
R143 Z.n4 Z.n3 92.5
R144 Z.n7 Z.n1 92.5
R145 Z.n6 Z.n4 50.009
R146 Z.n7 Z.n6 37.882
R147 Z Z.n8 33.129
R148 Z.n13 Z 30.117
R149 Z.n14 Z.t8 26.595
R150 Z.n14 Z.t7 26.595
R151 Z.n0 Z.t1 26.595
R152 Z.n0 Z.t2 26.595
R153 Z.n9 Z.t4 26.595
R154 Z.n9 Z.t3 26.595
R155 Z.n11 Z.t6 26.595
R156 Z.n11 Z.t5 26.595
R157 Z.n1 Z.t13 24.923
R158 Z.n1 Z.t14 24.923
R159 Z.n2 Z.t15 24.923
R160 Z.n2 Z.t0 24.923
R161 Z.n3 Z.t11 24.923
R162 Z.n3 Z.t9 24.923
R163 Z.n5 Z.t12 24.923
R164 Z.n5 Z.t10 24.923
R165 Z.n16 Z 24.094
R166 Z Z.n7 23.073
R167 Z Z.n13 14.305
R168 Z Z.n10 8.282
R169 Z.n13 Z.n12 6.422
R170 Z.n16 Z.n15 6.422
R171 Z.n12 Z 3.392
R172 Z.n15 Z 3.392
R173 Z.n10 Z 3.296
R174 Z.n13 Z 3.296
R175 Z Z.n16 3.296
R176 Z.n8 Z 2.863
R177 Z.n10 Z 1.505
R178 Z.n8 Z 1.505
R179 a_193_47.n8 a_193_47.t15 229.414
R180 a_193_47.n4 a_193_47.n3 164.782
R181 a_193_47.t14 a_193_47.n13 117.423
R182 a_193_47.n4 a_193_47.n2 101.535
R183 a_193_47.n5 a_193_47.n1 101.535
R184 a_193_47.n6 a_193_47.n0 101.535
R185 a_193_47.n12 a_193_47.n11 92.5
R186 a_193_47.n10 a_193_47.n9 92.5
R187 a_193_47.n8 a_193_47.n7 92.5
R188 a_193_47.n13 a_193_47.n6 66.494
R189 a_193_47.n6 a_193_47.n5 63.247
R190 a_193_47.n5 a_193_47.n4 63.247
R191 a_193_47.n13 a_193_47.n12 53.612
R192 a_193_47.n10 a_193_47.n8 51.2
R193 a_193_47.n12 a_193_47.n10 51.2
R194 a_193_47.n3 a_193_47.t4 28.615
R195 a_193_47.n3 a_193_47.t0 24.923
R196 a_193_47.n2 a_193_47.t5 24.923
R197 a_193_47.n2 a_193_47.t1 24.923
R198 a_193_47.n1 a_193_47.t6 24.923
R199 a_193_47.n1 a_193_47.t2 24.923
R200 a_193_47.n0 a_193_47.t7 24.923
R201 a_193_47.n0 a_193_47.t3 24.923
R202 a_193_47.n7 a_193_47.t8 24.923
R203 a_193_47.n7 a_193_47.t11 24.923
R204 a_193_47.n9 a_193_47.t9 24.923
R205 a_193_47.n9 a_193_47.t12 24.923
R206 a_193_47.n11 a_193_47.t10 24.923
R207 a_193_47.n11 a_193_47.t13 24.923
R208 VNB VNB.t8 6053.91
R209 VNB.t7 VNB.t15 4714.29
R210 VNB.t4 VNB.t0 2127.47
R211 VNB.t9 VNB.t16 2030.77
R212 VNB.t12 VNB.t9 2030.77
R213 VNB.t10 VNB.t12 2030.77
R214 VNB.t13 VNB.t10 2030.77
R215 VNB.t11 VNB.t13 2030.77
R216 VNB.t14 VNB.t11 2030.77
R217 VNB.t15 VNB.t14 2030.77
R218 VNB.t3 VNB.t7 2030.77
R219 VNB.t6 VNB.t3 2030.77
R220 VNB.t2 VNB.t6 2030.77
R221 VNB.t5 VNB.t2 2030.77
R222 VNB.t1 VNB.t5 2030.77
R223 VNB.t0 VNB.t1 2030.77
R224 VNB.t8 VNB.t4 2030.77
R225 TE.n8 TE.t8 265.099
R226 TE.n0 TE.t7 263.493
R227 TE.n7 TE.t9 152.633
R228 TE.n6 TE.n5 141.386
R229 TE.n1 TE.n0 134.96
R230 TE.n2 TE.n1 134.96
R231 TE.n3 TE.n2 134.96
R232 TE.n4 TE.n3 134.96
R233 TE.n5 TE.n4 134.96
R234 TE.n6 TE.t4 128.533
R235 TE.n5 TE.t0 128.533
R236 TE.n4 TE.t1 128.533
R237 TE.n3 TE.t5 128.533
R238 TE.n2 TE.t2 128.533
R239 TE.n1 TE.t6 128.533
R240 TE.n0 TE.t3 128.533
R241 TE.n7 TE.n6 110.86
R242 TE.n9 TE.n8 97.909
R243 TE.n8 TE.n7 40.166
R244 TE.n9 TE 14.889
R245 TE TE.n9 2.873
R246 VGND.n2 VGND.t0 194.682
R247 VGND.n1 VGND.n0 106.463
R248 VGND.n6 VGND.n5 106.463
R249 VGND.n11 VGND.n10 106.463
R250 VGND.n16 VGND.n15 106.463
R251 VGND.n0 VGND.t4 24.923
R252 VGND.n0 VGND.t1 24.923
R253 VGND.n5 VGND.t5 24.923
R254 VGND.n5 VGND.t2 24.923
R255 VGND.n10 VGND.t6 24.923
R256 VGND.n10 VGND.t7 24.923
R257 VGND.n15 VGND.t3 24.923
R258 VGND.n15 VGND.t8 24.923
R259 VGND.n2 VGND.n1 8.623
R260 VGND.n4 VGND.n3 4.65
R261 VGND.n7 VGND.n6 4.65
R262 VGND.n9 VGND.n8 4.65
R263 VGND.n12 VGND.n11 4.65
R264 VGND.n14 VGND.n13 4.65
R265 VGND.n17 VGND.n16 3.932
R266 VGND.n4 VGND.n2 0.524
R267 VGND.n17 VGND.n14 0.137
R268 VGND VGND.n17 0.121
R269 VGND.n7 VGND.n4 0.119
R270 VGND.n9 VGND.n7 0.119
R271 VGND.n12 VGND.n9 0.119
R272 VGND.n14 VGND.n12 0.119
C0 VGND VPWR 0.17fF
C1 VPB A 0.11fF
C2 Z A 0.97fF
C3 VPB VPWR 0.16fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__fa_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__fa_1 COUT CIN VGND VPWR SUM A B VNB VPB
X0 a_76_199.t2 B.t0 a_208_47.t1 VNB.t11 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1 VGND.t8 A.t0 a_382_47.t2 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 a_738_413.t3 A.t1 VPWR.t8 VPB.t13 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3 a_1091_47.t1 CIN.t0 a_995_47.t1 VNB.t5 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 VPWR.t1 CIN.t1 a_738_413.t0 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 a_382_413.t0 B.t1 VPWR.t2 VPB.t7 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 a_1163_47.t0 B.t2 a_1091_47.t0 VNB.t10 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7 VPWR.t5 A.t2 a_382_413.t2 VPB.t12 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 a_995_47.t2 a_76_199.t4 a_738_47.t2 VNB.t13 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9 a_382_413.t1 CIN.t2 a_76_199.t0 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10 SUM.t0 a_995_47.t4 VGND.t0 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 a_208_47.t0 A.t3 VGND.t6 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12 VGND.t1 CIN.t3 a_738_47.t1 VNB.t6 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13 a_76_199.t3 B.t3 a_208_413.t0 VPB.t6 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14 a_208_413.t1 A.t4 VPWR.t7 VPB.t11 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15 a_738_413.t1 B.t4 VPWR.t3 VPB.t5 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16 VGND.t7 A.t5 a_1163_47.t1 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17 a_738_47.t0 B.t5 VGND.t2 VNB.t9 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18 a_738_47.t3 A.t6 VGND.t5 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19 a_1163_413.t0 B.t6 a_1091_413.t0 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20 VPWR.t6 A.t7 a_1163_413.t1 VPB.t10 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21 a_382_47.t0 CIN.t4 a_76_199.t1 VNB.t7 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22 a_382_47.t1 B.t7 VGND.t3 VNB.t8 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23 SUM.t1 a_995_47.t5 VPWR.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X24 a_995_47.t3 a_76_199.t5 a_738_413.t2 VPB.t9 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X25 VPWR.t4 a_76_199.t6 COUT.t1 VPB.t8 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X26 a_1091_413.t1 CIN.t5 a_995_47.t0 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X27 VGND.t4 a_76_199.t7 COUT.t0 VNB.t12 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
R0 B.n0 B.t0 384.528
R1 B.n1 B.t2 361.151
R2 B.n2 B.t7 351.86
R3 B.n3 B.t1 297.233
R4 B.n4 B.n2 209.939
R5 B.n1 B.t6 177.693
R6 B.n0 B.t3 156.381
R7 B.n2 B.t5 109.214
R8 B.n3 B.t4 102.658
R9 B.n6 B.n0 81.92
R10 B.n4 B.n3 50.82
R11 B.n5 B.n1 11.366
R12 B.n5 B.n4 9.853
R13 B.n6 B.n5 6.213
R14 B B.n6 2.72
R15 a_208_47.t0 a_208_47.t1 85.714
R16 a_76_199.n1 a_76_199.t5 373.281
R17 a_76_199.n5 a_76_199.n4 368.565
R18 a_76_199.n0 a_76_199.t6 241.534
R19 a_76_199.n0 a_76_199.t7 169.234
R20 a_76_199.n1 a_76_199.t4 167.628
R21 a_76_199.n3 a_76_199.n1 103.72
R22 a_76_199.n3 a_76_199.n2 93.314
R23 a_76_199.n4 a_76_199.n0 76
R24 a_76_199.n4 a_76_199.n3 72.157
R25 a_76_199.t0 a_76_199.n5 63.321
R26 a_76_199.n5 a_76_199.t3 63.321
R27 a_76_199.n2 a_76_199.t1 38.571
R28 a_76_199.n2 a_76_199.t2 38.571
R29 VNB.t8 VNB.t9 6082.35
R30 VNB VNB.t12 6053.91
R31 VNB.t10 VNB.t3 3105.88
R32 VNB.t13 VNB.t5 3105.88
R33 VNB.t2 VNB.t11 2911.76
R34 VNB.t4 VNB.t13 2879.41
R35 VNB.t6 VNB.t4 2717.65
R36 VNB.t9 VNB.t6 2717.65
R37 VNB.t0 VNB.t8 2717.65
R38 VNB.t7 VNB.t0 2717.65
R39 VNB.t11 VNB.t7 2717.65
R40 VNB.t3 VNB.t1 2331.37
R41 VNB.t12 VNB.t2 2331.37
R42 VNB.t5 VNB.t10 2329.41
R43 A.n0 A.t1 361.136
R44 A.n1 A.t7 342.296
R45 A.n7 A.t4 332.043
R46 A.n3 A.t2 323.475
R47 A.n3 A.t0 217.435
R48 A.n1 A.t5 197.18
R49 A.n5 A.t3 193.692
R50 A.n0 A.t6 177.722
R51 A.n4 A.n3 89.183
R52 A.n6 A.n5 12.496
R53 A.n2 A.n1 11.988
R54 A.n2 A.n0 9.806
R55 A.n8 A.n7 8.764
R56 A.n8 A.n4 3.719
R57 A.n7 A.n6 2.677
R58 A A.n9 2.133
R59 A.n4 A.n2 1.557
R60 A.n9 A.n8 0.581
R61 a_382_47.n0 a_382_47.t1 312.418
R62 a_382_47.n0 a_382_47.t2 38.571
R63 a_382_47.t0 a_382_47.n0 38.571
R64 VGND.n6 VGND.t2 146.78
R65 VGND.n3 VGND.n2 111.433
R66 VGND.n20 VGND.n19 107.239
R67 VGND.n1 VGND.n0 106.463
R68 VGND.n11 VGND.n10 106.463
R69 VGND.n19 VGND.t6 60
R70 VGND.n2 VGND.t0 46.857
R71 VGND.n2 VGND.t7 38.571
R72 VGND.n0 VGND.t5 38.571
R73 VGND.n0 VGND.t1 38.571
R74 VGND.n10 VGND.t3 38.571
R75 VGND.n10 VGND.t8 38.571
R76 VGND.n19 VGND.t4 25.428
R77 VGND.n5 VGND.n4 4.65
R78 VGND.n7 VGND.n6 4.65
R79 VGND.n9 VGND.n8 4.65
R80 VGND.n12 VGND.n11 4.65
R81 VGND.n14 VGND.n13 4.65
R82 VGND.n16 VGND.n15 4.65
R83 VGND.n18 VGND.n17 4.65
R84 VGND.n3 VGND.n1 4.102
R85 VGND.n21 VGND.n20 3.932
R86 VGND.n21 VGND.n18 0.137
R87 VGND.n5 VGND.n3 0.135
R88 VGND VGND.n21 0.121
R89 VGND.n7 VGND.n5 0.119
R90 VGND.n9 VGND.n7 0.119
R91 VGND.n12 VGND.n9 0.119
R92 VGND.n14 VGND.n12 0.119
R93 VGND.n16 VGND.n14 0.119
R94 VGND.n18 VGND.n16 0.119
R95 VPWR.n6 VPWR.t3 370.56
R96 VPWR.n20 VPWR.n19 312.98
R97 VPWR.n3 VPWR.n2 310.197
R98 VPWR.n1 VPWR.n0 306.463
R99 VPWR.n11 VPWR.n10 306.463
R100 VPWR.n2 VPWR.t6 98.5
R101 VPWR.n19 VPWR.t7 98.5
R102 VPWR.n0 VPWR.t8 63.321
R103 VPWR.n0 VPWR.t1 63.321
R104 VPWR.n10 VPWR.t2 63.321
R105 VPWR.n10 VPWR.t5 63.321
R106 VPWR.n2 VPWR.t0 27.955
R107 VPWR.n19 VPWR.t4 27.955
R108 VPWR.n5 VPWR.n4 4.65
R109 VPWR.n7 VPWR.n6 4.65
R110 VPWR.n9 VPWR.n8 4.65
R111 VPWR.n12 VPWR.n11 4.65
R112 VPWR.n14 VPWR.n13 4.65
R113 VPWR.n16 VPWR.n15 4.65
R114 VPWR.n18 VPWR.n17 4.65
R115 VPWR.n3 VPWR.n1 4.102
R116 VPWR.n21 VPWR.n20 3.932
R117 VPWR.n21 VPWR.n18 0.137
R118 VPWR.n5 VPWR.n3 0.135
R119 VPWR VPWR.n21 0.121
R120 VPWR.n7 VPWR.n5 0.119
R121 VPWR.n9 VPWR.n7 0.119
R122 VPWR.n12 VPWR.n9 0.119
R123 VPWR.n14 VPWR.n12 0.119
R124 VPWR.n16 VPWR.n14 0.119
R125 VPWR.n18 VPWR.n16 0.119
R126 a_738_413.n1 a_738_413.n0 673.847
R127 a_738_413.n0 a_738_413.t2 75.047
R128 a_738_413.n0 a_738_413.t3 63.321
R129 a_738_413.t0 a_738_413.n1 63.321
R130 a_738_413.n1 a_738_413.t1 63.321
R131 VPB.t7 VPB.t5 556.386
R132 VPB.t10 VPB.t0 292.99
R133 VPB.t8 VPB.t11 292.99
R134 VPB.t4 VPB.t10 284.112
R135 VPB.t9 VPB.t3 284.112
R136 VPB.t11 VPB.t6 266.355
R137 VPB.t13 VPB.t9 263.395
R138 VPB.t1 VPB.t13 248.598
R139 VPB.t5 VPB.t1 248.598
R140 VPB.t12 VPB.t7 248.598
R141 VPB.t2 VPB.t12 248.598
R142 VPB.t6 VPB.t2 248.598
R143 VPB.t3 VPB.t4 213.084
R144 VPB VPB.t8 189.408
R145 CIN.n0 CIN.t0 373.281
R146 CIN.n1 CIN.t3 346.02
R147 CIN.n2 CIN.t2 325.081
R148 CIN.n3 CIN.n2 281.437
R149 CIN.n2 CIN.t4 215.828
R150 CIN.n1 CIN.t1 193.335
R151 CIN.n0 CIN.t5 167.628
R152 CIN.n4 CIN.n3 88.425
R153 CIN.n3 CIN.n1 76
R154 CIN.n4 CIN.n0 76
R155 CIN CIN.n4 5.376
R156 a_995_47.n3 a_995_47.n2 420.271
R157 a_995_47.n0 a_995_47.t5 241.534
R158 a_995_47.n2 a_995_47.n1 211.138
R159 a_995_47.n0 a_995_47.t4 169.234
R160 a_995_47.n3 a_995_47.t3 91.464
R161 a_995_47.n2 a_995_47.n0 76
R162 a_995_47.t0 a_995_47.n3 63.321
R163 a_995_47.n1 a_995_47.t2 55.714
R164 a_995_47.n1 a_995_47.t1 38.571
R165 a_1091_47.t0 a_1091_47.t1 60
R166 a_382_413.t0 a_382_413.n0 731.857
R167 a_382_413.n0 a_382_413.t2 63.321
R168 a_382_413.n0 a_382_413.t1 63.321
R169 a_1163_47.t0 a_1163_47.t1 94.285
R170 a_738_47.n1 a_738_47.n0 273.847
R171 a_738_47.n0 a_738_47.t2 45.714
R172 a_738_47.n0 a_738_47.t3 38.571
R173 a_738_47.n1 a_738_47.t1 38.571
R174 a_738_47.t0 a_738_47.n1 38.571
R175 SUM.t1 SUM 465.7
R176 SUM.n1 SUM.t1 462.98
R177 SUM.n0 SUM.t0 117.423
R178 SUM.n3 SUM 11.442
R179 SUM.n2 SUM.n1 8.8
R180 SUM SUM.n0 6.56
R181 SUM.n0 SUM 4.32
R182 SUM SUM.n3 1.745
R183 SUM SUM.n2 1.551
R184 SUM.n3 SUM 1.44
R185 SUM.n2 SUM 1.28
R186 SUM.n1 SUM 0.8
R187 a_208_413.t0 a_208_413.t1 140.714
R188 a_1091_413.t0 a_1091_413.t1 98.5
R189 a_1163_413.t0 a_1163_413.t1 154.785
R190 COUT COUT.t1 495.407
R191 COUT.n1 COUT.t1 451.615
R192 COUT.n0 COUT.t0 117.423
R193 COUT.n1 COUT.n0 75.476
R194 COUT.n0 COUT 6.646
R195 COUT COUT.n1 0.492
C0 B A 1.37fF
C1 B CIN 0.59fF
C2 VPWR SUM 0.10fF
C3 CIN A 0.49fF
C4 VPWR VPB 0.14fF
C5 B VPWR 0.26fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__fa_2.ext - technology: sky130A

.subckt sky130_fd_sc_hd__fa_2 COUT SUM A B CIN VGND VPWR VNB VPB
X0 a_1171_369.t0 CIN.t0 a_1086_47.t1 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1 VGND.t0 CIN.t1 a_829_47.t0 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 VGND.t8 a_1086_47.t4 SUM.t1 VNB.t13 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 COUT.t3 a_80_21.t4 VPWR.t8 VPB.t15 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 a_829_369.t3 A.t0 VPWR.t3 VPB.t9 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X5 VPWR.t0 CIN.t2 a_829_369.t0 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X6 a_473_371.t1 B.t0 VPWR.t1 VPB.t5 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=630000u l=150000u
X7 a_294_47.t1 A.t1 VGND.t3 VNB.t8 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 VPWR.t4 A.t2 a_473_371.t2 VPB.t10 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=630000u l=150000u
X9 a_829_369.t1 B.t1 VPWR.t2 VPB.t6 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X10 a_829_47.t2 B.t2 VGND.t1 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11 a_829_47.t3 A.t3 VGND.t4 VNB.t9 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12 a_473_371.t0 CIN.t3 a_80_21.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=630000u l=150000u
X13 a_473_47.t0 CIN.t4 a_80_21.t1 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14 a_473_47.t1 B.t3 VGND.t2 VNB.t5 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15 VPWR.t10 a_1086_47.t5 SUM.t3 VPB.t14 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16 VGND.t9 a_80_21.t5 COUT.t1 VNB.t14 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X17 COUT.t0 a_80_21.t6 VGND.t10 VNB.t15 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X18 SUM.t2 a_1086_47.t6 VPWR.t9 VPB.t13 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X19 a_80_21.t2 B.t4 a_289_371.t0 VPB.t7 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=630000u l=150000u
X20 a_80_21.t3 B.t5 a_294_47.t0 VNB.t6 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21 VGND.t5 A.t4 a_473_47.t2 VNB.t10 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22 SUM.t0 a_1086_47.t7 VGND.t7 VNB.t12 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X23 VPWR.t7 a_80_21.t7 COUT.t2 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X24 a_289_371.t1 A.t5 VPWR.t5 VPB.t11 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=630000u l=150000u
X25 a_1194_47.t0 CIN.t5 a_1086_47.t0 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X26 a_1086_47.t2 a_80_21.t8 a_829_47.t1 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X27 VGND.t6 A.t6 a_1266_47.t1 VNB.t11 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X28 a_1266_371.t0 B.t6 a_1171_369.t1 VPB.t8 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=630000u l=150000u
X29 VPWR.t6 A.t7 a_1266_371.t1 VPB.t12 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=630000u l=150000u
X30 a_1266_47.t0 B.t7 a_1194_47.t1 VNB.t7 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X31 a_1086_47.t3 a_80_21.t9 a_829_369.t2 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
R0 CIN.n3 CIN.t5 321.868
R1 CIN.n0 CIN.t1 320.313
R2 CIN.n1 CIN.t3 291.341
R3 CIN.n2 CIN.n1 267.328
R4 CIN.n1 CIN.t4 215.828
R5 CIN.n3 CIN.t0 183.694
R6 CIN.n0 CIN.t2 183.694
R7 CIN.n4 CIN.n2 84.871
R8 CIN.n4 CIN.n3 80.096
R9 CIN.n2 CIN.n0 76
R10 CIN CIN.n4 9.472
R11 a_1086_47.n5 a_1086_47.n4 416.706
R12 a_1086_47.n4 a_1086_47.n0 222.095
R13 a_1086_47.n1 a_1086_47.t5 212.079
R14 a_1086_47.n2 a_1086_47.t6 212.079
R15 a_1086_47.n1 a_1086_47.t4 151.463
R16 a_1086_47.n2 a_1086_47.t7 145.621
R17 a_1086_47.n0 a_1086_47.t0 55.714
R18 a_1086_47.n0 a_1086_47.t2 55.714
R19 a_1086_47.n5 a_1086_47.t3 43.093
R20 a_1086_47.t1 a_1086_47.n5 41.554
R21 a_1086_47.n4 a_1086_47.n3 40.001
R22 a_1086_47.n3 a_1086_47.n1 30.235
R23 a_1086_47.n3 a_1086_47.n2 20.259
R24 a_1171_369.t0 a_1171_369.t1 96.234
R25 VPB.t5 VPB.t6 556.386
R26 VPB.t8 VPB.t12 319.626
R27 VPB.t12 VPB.t13 281.152
R28 VPB.t2 VPB.t8 281.152
R29 VPB.t7 VPB.t0 281.152
R30 VPB.t3 VPB.t11 281.152
R31 VPB.t9 VPB.t4 263.395
R32 VPB.t11 VPB.t7 263.395
R33 VPB.t4 VPB.t2 251.557
R34 VPB.t13 VPB.t14 248.598
R35 VPB.t1 VPB.t9 248.598
R36 VPB.t6 VPB.t1 248.598
R37 VPB.t10 VPB.t5 248.598
R38 VPB.t0 VPB.t10 248.598
R39 VPB.t15 VPB.t3 248.598
R40 VPB VPB.t15 195.327
R41 a_829_47.n1 a_829_47.n0 273.847
R42 a_829_47.n0 a_829_47.t1 45.714
R43 a_829_47.n0 a_829_47.t3 38.571
R44 a_829_47.t0 a_829_47.n1 38.571
R45 a_829_47.n1 a_829_47.t2 38.571
R46 VGND.n2 VGND.t8 197.778
R47 VGND.n34 VGND.t10 190.063
R48 VGND.n16 VGND.t1 146.78
R49 VGND.n30 VGND.n29 107.239
R50 VGND.n1 VGND.n0 106.463
R51 VGND.n12 VGND.n11 106.463
R52 VGND.n21 VGND.n20 106.463
R53 VGND.n29 VGND.t9 48.285
R54 VGND.n0 VGND.t7 46.857
R55 VGND.n0 VGND.t6 38.571
R56 VGND.n11 VGND.t4 38.571
R57 VGND.n11 VGND.t0 38.571
R58 VGND.n20 VGND.t2 38.571
R59 VGND.n20 VGND.t5 38.571
R60 VGND.n29 VGND.t3 38.571
R61 VGND.n35 VGND.n34 7.285
R62 VGND.n2 VGND.n1 5.533
R63 VGND.n4 VGND.n3 4.65
R64 VGND.n6 VGND.n5 4.65
R65 VGND.n8 VGND.n7 4.65
R66 VGND.n10 VGND.n9 4.65
R67 VGND.n13 VGND.n12 4.65
R68 VGND.n15 VGND.n14 4.65
R69 VGND.n17 VGND.n16 4.65
R70 VGND.n19 VGND.n18 4.65
R71 VGND.n22 VGND.n21 4.65
R72 VGND.n24 VGND.n23 4.65
R73 VGND.n26 VGND.n25 4.65
R74 VGND.n28 VGND.n27 4.65
R75 VGND.n31 VGND.n30 4.65
R76 VGND.n33 VGND.n32 4.65
R77 VGND.n4 VGND.n2 0.245
R78 VGND.n6 VGND.n4 0.119
R79 VGND.n8 VGND.n6 0.119
R80 VGND.n10 VGND.n8 0.119
R81 VGND.n13 VGND.n10 0.119
R82 VGND.n15 VGND.n13 0.119
R83 VGND.n17 VGND.n15 0.119
R84 VGND.n19 VGND.n17 0.119
R85 VGND.n22 VGND.n19 0.119
R86 VGND.n24 VGND.n22 0.119
R87 VGND.n26 VGND.n24 0.119
R88 VGND.n28 VGND.n26 0.119
R89 VGND.n31 VGND.n28 0.119
R90 VGND.n33 VGND.n31 0.119
R91 VGND.n35 VGND.n33 0.119
R92 VGND VGND.n35 0.022
R93 VNB VNB.t15 6102.26
R94 VNB.t5 VNB.t4 6082.35
R95 VNB.t3 VNB.t0 3494.12
R96 VNB.t7 VNB.t11 3105.88
R97 VNB.t8 VNB.t6 3073.53
R98 VNB.t9 VNB.t3 2879.41
R99 VNB.t2 VNB.t9 2717.65
R100 VNB.t4 VNB.t2 2717.65
R101 VNB.t10 VNB.t5 2717.65
R102 VNB.t1 VNB.t10 2717.65
R103 VNB.t6 VNB.t1 2717.65
R104 VNB.t12 VNB.t13 2610.99
R105 VNB.t14 VNB.t8 2345.21
R106 VNB.t11 VNB.t12 2331.37
R107 VNB.t0 VNB.t7 2329.41
R108 VNB.t15 VNB.t14 2030.77
R109 SUM SUM.n0 229.955
R110 SUM SUM.n1 88.985
R111 SUM.n1 SUM.t0 47.076
R112 SUM.n0 SUM.t3 26.595
R113 SUM.n0 SUM.t2 26.595
R114 SUM.n1 SUM.t1 24.923
R115 a_80_21.n0 a_80_21.t9 337.934
R116 a_80_21.n7 a_80_21.n6 248.376
R117 a_80_21.n3 a_80_21.t7 212.079
R118 a_80_21.n4 a_80_21.t4 212.079
R119 a_80_21.n0 a_80_21.t8 167.628
R120 a_80_21.n3 a_80_21.t5 139.779
R121 a_80_21.n4 a_80_21.t6 139.779
R122 a_80_21.n2 a_80_21.n0 104.229
R123 a_80_21.n6 a_80_21.n5 97.458
R124 a_80_21.n2 a_80_21.n1 93.285
R125 a_80_21.n6 a_80_21.n2 71.31
R126 a_80_21.n7 a_80_21.t2 59.412
R127 a_80_21.t0 a_80_21.n7 42.214
R128 a_80_21.n1 a_80_21.t1 38.571
R129 a_80_21.n1 a_80_21.t3 38.571
R130 a_80_21.n5 a_80_21.n4 33.593
R131 a_80_21.n5 a_80_21.n3 27.751
R132 VPWR.n30 VPWR.n29 306.463
R133 VPWR.n21 VPWR.n20 306.463
R134 VPWR.n12 VPWR.n11 306.463
R135 VPWR.n1 VPWR.n0 306.463
R136 VPWR.n16 VPWR.t2 228.681
R137 VPWR.n2 VPWR.t10 214.209
R138 VPWR.n34 VPWR.t8 204.201
R139 VPWR.n0 VPWR.t6 57.849
R140 VPWR.n29 VPWR.t5 46.904
R141 VPWR.n29 VPWR.t7 43.926
R142 VPWR.n20 VPWR.t1 42.214
R143 VPWR.n20 VPWR.t4 42.214
R144 VPWR.n11 VPWR.t3 41.554
R145 VPWR.n11 VPWR.t0 41.554
R146 VPWR.n0 VPWR.t9 32.982
R147 VPWR.n35 VPWR.n34 7.285
R148 VPWR.n4 VPWR.n3 4.65
R149 VPWR.n6 VPWR.n5 4.65
R150 VPWR.n8 VPWR.n7 4.65
R151 VPWR.n10 VPWR.n9 4.65
R152 VPWR.n13 VPWR.n12 4.65
R153 VPWR.n15 VPWR.n14 4.65
R154 VPWR.n17 VPWR.n16 4.65
R155 VPWR.n19 VPWR.n18 4.65
R156 VPWR.n22 VPWR.n21 4.65
R157 VPWR.n24 VPWR.n23 4.65
R158 VPWR.n26 VPWR.n25 4.65
R159 VPWR.n28 VPWR.n27 4.65
R160 VPWR.n31 VPWR.n30 4.65
R161 VPWR.n33 VPWR.n32 4.65
R162 VPWR.n2 VPWR.n1 3.833
R163 VPWR.n4 VPWR.n2 0.349
R164 VPWR.n6 VPWR.n4 0.119
R165 VPWR.n8 VPWR.n6 0.119
R166 VPWR.n10 VPWR.n8 0.119
R167 VPWR.n13 VPWR.n10 0.119
R168 VPWR.n15 VPWR.n13 0.119
R169 VPWR.n17 VPWR.n15 0.119
R170 VPWR.n19 VPWR.n17 0.119
R171 VPWR.n22 VPWR.n19 0.119
R172 VPWR.n24 VPWR.n22 0.119
R173 VPWR.n26 VPWR.n24 0.119
R174 VPWR.n28 VPWR.n26 0.119
R175 VPWR.n31 VPWR.n28 0.119
R176 VPWR.n33 VPWR.n31 0.119
R177 VPWR.n35 VPWR.n33 0.119
R178 VPWR VPWR.n35 0.022
R179 COUT COUT.n0 198.878
R180 COUT.n2 COUT.n1 146.398
R181 COUT.n1 COUT.t2 26.595
R182 COUT.n1 COUT.t3 26.595
R183 COUT.n0 COUT.t1 24.923
R184 COUT.n0 COUT.t0 24.923
R185 COUT COUT.n3 10.057
R186 COUT.n3 COUT 8.62
R187 COUT.n3 COUT.n2 5.466
R188 COUT.n2 COUT 5.034
R189 A.n0 A.t0 325.789
R190 A.n5 A.t5 300.981
R191 A.n1 A.t7 300.981
R192 A.n3 A.t2 289.735
R193 A.n3 A.t4 217.435
R194 A.n1 A.t6 206.188
R195 A.n5 A.t1 205.7
R196 A.n0 A.t3 177.722
R197 A.n2 A.n1 107.608
R198 A.n4 A.n3 89.183
R199 A A.n5 84.914
R200 A.n2 A.n0 9.806
R201 A A.n4 9.664
R202 A.n4 A.n2 1.557
R203 a_829_369.n1 a_829_369.n0 673.847
R204 a_829_369.n0 a_829_369.t2 49.25
R205 a_829_369.n0 a_829_369.t3 41.554
R206 a_829_369.t0 a_829_369.n1 41.554
R207 a_829_369.n1 a_829_369.t1 41.554
R208 B.n0 B.t3 393.633
R209 B.n1 B.t0 334.186
R210 B.n5 B.t5 325.081
R211 B.n3 B.t7 325.081
R212 B.n5 B.t4 182.088
R213 B.n3 B.t6 182.088
R214 B.n2 B.n0 173.233
R215 B.n1 B.t1 136.566
R216 B.n4 B.n3 99.558
R217 B.n0 B.t2 91.58
R218 B B.n5 85.142
R219 B.n2 B.n1 22.407
R220 B B.n4 10.653
R221 B.n4 B.n2 10.135
R222 a_473_371.n0 a_473_371.t1 700.368
R223 a_473_371.n0 a_473_371.t2 42.214
R224 a_473_371.t0 a_473_371.n0 42.214
R225 a_294_47.t0 a_294_47.t1 92.857
R226 a_473_47.n0 a_473_47.t1 312.418
R227 a_473_47.n0 a_473_47.t2 38.571
R228 a_473_47.t0 a_473_47.n0 38.571
R229 a_289_371.t0 a_289_371.t1 92.246
R230 a_1194_47.t0 a_1194_47.t1 60
R231 a_1266_47.t0 a_1266_47.t1 94.285
R232 a_1266_371.t0 a_1266_371.t1 121.952
C0 VPWR COUT 0.19fF
C1 VPWR VPB 0.17fF
C2 VGND SUM 0.19fF
C3 CIN A 0.47fF
C4 A B 1.43fF
C5 COUT VGND 0.17fF
C6 VPWR SUM 0.20fF
C7 VPWR B 0.33fF
C8 CIN B 0.53fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__fa_4.ext - technology: sky130A

.subckt sky130_fd_sc_hd__fa_4 COUT SUM A B CIN VGND VPWR VNB VPB
X0 a_1014_369.t1 B.t0 VPWR.t8 VPB.t11 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1 VPWR.t13 CIN.t0 a_1014_369.t2 VPB.t15 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X2 VPWR.t0 A.t0 a_658_369.t2 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X3 VGND.t12 A.t1 a_658_47.t2 VNB.t17 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 a_79_21.t1 B.t1 a_456_371.t0 VPB.t10 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=630000u l=150000u
X5 a_658_369.t1 CIN.t1 a_79_21.t2 VPB.t16 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X6 VPWR.t4 a_1271_47.t4 SUM.t7 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 a_461_47.t1 A.t2 VGND.t10 VNB.t16 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 VPWR.t10 a_79_21.t4 COUT.t7 VPB.t12 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 SUM.t6 a_1271_47.t5 VPWR.t5 VPB.t5 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 a_1271_47.t0 a_79_21.t5 a_1014_47.t0 VNB.t11 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11 a_658_47.t1 CIN.t2 a_79_21.t3 VNB.t10 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12 a_658_47.t0 B.t2 VGND.t5 VNB.t7 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13 COUT.t6 a_79_21.t6 VPWR.t11 VPB.t13 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14 a_456_371.t1 A.t3 VPWR.t1 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=630000u l=150000u
X15 a_1451_47.t0 B.t3 a_1379_47.t0 VNB.t6 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16 VPWR.t12 a_79_21.t7 COUT.t5 VPB.t14 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17 VGND.t7 a_79_21.t8 COUT.t3 VNB.t12 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X18 VGND.t8 a_79_21.t9 COUT.t2 VNB.t13 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X19 VPWR.t6 a_1271_47.t6 SUM.t5 VPB.t6 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X20 VGND.t0 a_1271_47.t7 SUM.t3 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X21 VGND.t1 a_1271_47.t8 SUM.t2 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X22 a_1451_371.t0 B.t4 a_1356_369.t0 VPB.t9 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=630000u l=150000u
X23 a_79_21.t0 B.t5 a_461_47.t0 VNB.t5 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24 a_1014_47.t3 A.t4 VGND.t9 VNB.t15 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X25 a_1271_47.t1 a_79_21.t10 a_1014_369.t3 VPB.t18 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X26 COUT.t1 a_79_21.t11 VGND.t13 VNB.t18 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X27 a_658_369.t0 B.t6 VPWR.t9 VPB.t8 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X28 VPWR.t2 A.t5 a_1451_371.t1 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=630000u l=150000u
X29 a_1014_47.t1 B.t7 VGND.t4 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X30 a_1379_47.t1 CIN.t3 a_1271_47.t3 VNB.t9 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X31 VGND.t11 A.t6 a_1451_47.t1 VNB.t14 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X32 SUM.t1 a_1271_47.t9 VGND.t2 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X33 a_1356_369.t1 CIN.t4 a_1271_47.t2 VPB.t17 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X34 SUM.t0 a_1271_47.t10 VGND.t3 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X35 SUM.t4 a_1271_47.t11 VPWR.t7 VPB.t7 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X36 VGND.t6 CIN.t5 a_1014_47.t2 VNB.t8 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X37 a_1014_369.t0 A.t7 VPWR.t3 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X38 COUT.t4 a_79_21.t12 VPWR.t14 VPB.t19 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X39 COUT.t0 a_79_21.t13 VGND.t14 VNB.t19 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
R0 B.n0 B.t2 393.633
R1 B.n1 B.t6 332.579
R2 B.n5 B.t5 325.081
R3 B.n3 B.t3 325.081
R4 B.n5 B.t1 182.088
R5 B.n3 B.t4 182.088
R6 B.n2 B.n0 173.233
R7 B.n1 B.t0 136.566
R8 B.n4 B.n3 99.558
R9 B.n0 B.t7 91.58
R10 B B.n5 89.844
R11 B.n2 B.n1 22.407
R12 B B.n4 10.653
R13 B.n4 B.n2 10.135
R14 VPWR.n35 VPWR.n34 306.463
R15 VPWR.n26 VPWR.n25 306.463
R16 VPWR.n17 VPWR.n16 306.463
R17 VPWR.n6 VPWR.n5 306.463
R18 VPWR.n21 VPWR.t8 228.681
R19 VPWR.n2 VPWR.t6 214.161
R20 VPWR.n45 VPWR.t14 204.201
R21 VPWR.n40 VPWR.n39 177.606
R22 VPWR.n1 VPWR.n0 177.606
R23 VPWR.n5 VPWR.t2 57.849
R24 VPWR.n34 VPWR.t1 46.904
R25 VPWR.n34 VPWR.t10 43.926
R26 VPWR.n0 VPWR.t7 42.355
R27 VPWR.n25 VPWR.t9 41.554
R28 VPWR.n25 VPWR.t0 41.554
R29 VPWR.n16 VPWR.t3 41.554
R30 VPWR.n16 VPWR.t13 41.554
R31 VPWR.n5 VPWR.t5 32.982
R32 VPWR.n39 VPWR.t11 26.595
R33 VPWR.n39 VPWR.t12 26.595
R34 VPWR.n0 VPWR.t4 26.595
R35 VPWR.n2 VPWR.n1 14.882
R36 VPWR.n46 VPWR.n45 6.908
R37 VPWR.n4 VPWR.n3 4.65
R38 VPWR.n7 VPWR.n6 4.65
R39 VPWR.n9 VPWR.n8 4.65
R40 VPWR.n11 VPWR.n10 4.65
R41 VPWR.n13 VPWR.n12 4.65
R42 VPWR.n15 VPWR.n14 4.65
R43 VPWR.n18 VPWR.n17 4.65
R44 VPWR.n20 VPWR.n19 4.65
R45 VPWR.n22 VPWR.n21 4.65
R46 VPWR.n24 VPWR.n23 4.65
R47 VPWR.n27 VPWR.n26 4.65
R48 VPWR.n29 VPWR.n28 4.65
R49 VPWR.n31 VPWR.n30 4.65
R50 VPWR.n33 VPWR.n32 4.65
R51 VPWR.n36 VPWR.n35 4.65
R52 VPWR.n38 VPWR.n37 4.65
R53 VPWR.n42 VPWR.n41 4.65
R54 VPWR.n44 VPWR.n43 4.65
R55 VPWR.n41 VPWR.n40 3.764
R56 VPWR.n4 VPWR.n2 0.309
R57 VPWR.n7 VPWR.n4 0.119
R58 VPWR.n9 VPWR.n7 0.119
R59 VPWR.n11 VPWR.n9 0.119
R60 VPWR.n13 VPWR.n11 0.119
R61 VPWR.n15 VPWR.n13 0.119
R62 VPWR.n18 VPWR.n15 0.119
R63 VPWR.n20 VPWR.n18 0.119
R64 VPWR.n22 VPWR.n20 0.119
R65 VPWR.n24 VPWR.n22 0.119
R66 VPWR.n27 VPWR.n24 0.119
R67 VPWR.n29 VPWR.n27 0.119
R68 VPWR.n31 VPWR.n29 0.119
R69 VPWR.n33 VPWR.n31 0.119
R70 VPWR.n36 VPWR.n33 0.119
R71 VPWR.n38 VPWR.n36 0.119
R72 VPWR.n42 VPWR.n38 0.119
R73 VPWR.n44 VPWR.n42 0.119
R74 VPWR.n46 VPWR.n44 0.119
R75 VPWR VPWR.n46 0.02
R76 a_1014_369.n1 a_1014_369.n0 673.847
R77 a_1014_369.n1 a_1014_369.t3 49.25
R78 a_1014_369.n0 a_1014_369.t2 41.554
R79 a_1014_369.n0 a_1014_369.t1 41.554
R80 a_1014_369.t0 a_1014_369.n1 41.554
R81 VPB.t8 VPB.t11 556.386
R82 VPB.t10 VPB.t16 334.423
R83 VPB.t9 VPB.t2 319.626
R84 VPB.t4 VPB.t7 295.95
R85 VPB.t2 VPB.t5 281.152
R86 VPB.t17 VPB.t9 281.152
R87 VPB.t12 VPB.t1 281.152
R88 VPB.t3 VPB.t18 263.395
R89 VPB.t1 VPB.t10 263.395
R90 VPB.t18 VPB.t17 251.557
R91 VPB.t7 VPB.t6 248.598
R92 VPB.t5 VPB.t4 248.598
R93 VPB.t15 VPB.t3 248.598
R94 VPB.t11 VPB.t15 248.598
R95 VPB.t0 VPB.t8 248.598
R96 VPB.t16 VPB.t0 248.598
R97 VPB.t13 VPB.t12 248.598
R98 VPB.t14 VPB.t13 248.598
R99 VPB.t19 VPB.t14 248.598
R100 VPB VPB.t19 189.408
R101 CIN.n3 CIN.t3 321.868
R102 CIN.n0 CIN.t5 320.313
R103 CIN.n1 CIN.t1 289.734
R104 CIN.n2 CIN.n1 267.328
R105 CIN.n1 CIN.t2 215.828
R106 CIN.n3 CIN.t4 183.694
R107 CIN.n0 CIN.t0 183.694
R108 CIN.n4 CIN.n2 84.871
R109 CIN.n4 CIN.n3 80.096
R110 CIN.n2 CIN.n0 76
R111 CIN CIN.n4 9.472
R112 A.n0 A.t7 325.789
R113 A.n5 A.t3 300.981
R114 A.n1 A.t5 300.981
R115 A.n3 A.t0 288.127
R116 A.n3 A.t1 217.435
R117 A.n1 A.t6 206.188
R118 A.n5 A.t2 205.7
R119 A.n0 A.t4 177.722
R120 A.n2 A.n1 107.608
R121 A.n4 A.n3 89.183
R122 A A.n5 89.028
R123 A.n2 A.n0 9.806
R124 A A.n4 9.664
R125 A.n4 A.n2 1.557
R126 a_658_369.t0 a_658_369.n0 699.708
R127 a_658_369.n0 a_658_369.t2 41.554
R128 a_658_369.n0 a_658_369.t1 41.554
R129 a_658_47.t0 a_658_47.n0 312.418
R130 a_658_47.n0 a_658_47.t2 38.571
R131 a_658_47.n0 a_658_47.t1 38.571
R132 VGND.n2 VGND.t1 192.383
R133 VGND.n46 VGND.t14 190.063
R134 VGND.n22 VGND.t4 146.78
R135 VGND.n1 VGND.n0 116.217
R136 VGND.n41 VGND.n40 116.217
R137 VGND.n36 VGND.n35 107.239
R138 VGND.n6 VGND.n5 106.463
R139 VGND.n18 VGND.n17 106.463
R140 VGND.n27 VGND.n26 106.463
R141 VGND.n5 VGND.t3 56.263
R142 VGND.n35 VGND.t8 48.285
R143 VGND.n5 VGND.t11 38.571
R144 VGND.n17 VGND.t9 38.571
R145 VGND.n17 VGND.t6 38.571
R146 VGND.n26 VGND.t5 38.571
R147 VGND.n26 VGND.t12 38.571
R148 VGND.n35 VGND.t10 38.571
R149 VGND.n0 VGND.t2 24.923
R150 VGND.n0 VGND.t0 24.923
R151 VGND.n40 VGND.t13 24.923
R152 VGND.n40 VGND.t7 24.923
R153 VGND.n2 VGND.n1 8.859
R154 VGND.n47 VGND.n46 6.908
R155 VGND.n4 VGND.n3 4.65
R156 VGND.n8 VGND.n7 4.65
R157 VGND.n10 VGND.n9 4.65
R158 VGND.n12 VGND.n11 4.65
R159 VGND.n14 VGND.n13 4.65
R160 VGND.n16 VGND.n15 4.65
R161 VGND.n19 VGND.n18 4.65
R162 VGND.n21 VGND.n20 4.65
R163 VGND.n23 VGND.n22 4.65
R164 VGND.n25 VGND.n24 4.65
R165 VGND.n28 VGND.n27 4.65
R166 VGND.n30 VGND.n29 4.65
R167 VGND.n32 VGND.n31 4.65
R168 VGND.n34 VGND.n33 4.65
R169 VGND.n37 VGND.n36 4.65
R170 VGND.n39 VGND.n38 4.65
R171 VGND.n43 VGND.n42 4.65
R172 VGND.n45 VGND.n44 4.65
R173 VGND.n42 VGND.n41 3.764
R174 VGND.n7 VGND.n6 1.129
R175 VGND.n4 VGND.n2 0.309
R176 VGND.n8 VGND.n4 0.119
R177 VGND.n10 VGND.n8 0.119
R178 VGND.n12 VGND.n10 0.119
R179 VGND.n14 VGND.n12 0.119
R180 VGND.n16 VGND.n14 0.119
R181 VGND.n19 VGND.n16 0.119
R182 VGND.n21 VGND.n19 0.119
R183 VGND.n23 VGND.n21 0.119
R184 VGND.n25 VGND.n23 0.119
R185 VGND.n28 VGND.n25 0.119
R186 VGND.n30 VGND.n28 0.119
R187 VGND.n32 VGND.n30 0.119
R188 VGND.n34 VGND.n32 0.119
R189 VGND.n37 VGND.n34 0.119
R190 VGND.n39 VGND.n37 0.119
R191 VGND.n43 VGND.n39 0.119
R192 VGND.n45 VGND.n43 0.119
R193 VGND.n47 VGND.n45 0.119
R194 VGND VGND.n47 0.02
R195 VNB.t7 VNB.t4 6082.35
R196 VNB VNB.t19 6053.91
R197 VNB.t11 VNB.t9 3494.12
R198 VNB.t5 VNB.t10 3300
R199 VNB.t6 VNB.t14 3105.88
R200 VNB.t16 VNB.t5 3073.53
R201 VNB.t15 VNB.t11 2879.41
R202 VNB.t8 VNB.t15 2717.65
R203 VNB.t4 VNB.t8 2717.65
R204 VNB.t17 VNB.t7 2717.65
R205 VNB.t10 VNB.t17 2717.65
R206 VNB.t14 VNB.t3 2524.78
R207 VNB.t3 VNB.t0 2417.58
R208 VNB.t13 VNB.t16 2345.21
R209 VNB.t9 VNB.t6 2329.41
R210 VNB.t2 VNB.t1 2030.77
R211 VNB.t0 VNB.t2 2030.77
R212 VNB.t18 VNB.t13 2030.77
R213 VNB.t12 VNB.t18 2030.77
R214 VNB.t19 VNB.t12 2030.77
R215 a_456_371.t0 a_456_371.t1 92.246
R216 a_79_21.n0 a_79_21.t10 337.934
R217 a_79_21.n13 a_79_21.n12 247.748
R218 a_79_21.n8 a_79_21.t4 212.079
R219 a_79_21.n9 a_79_21.t6 212.079
R220 a_79_21.n3 a_79_21.t7 212.079
R221 a_79_21.n5 a_79_21.t12 212.079
R222 a_79_21.n0 a_79_21.t5 167.628
R223 a_79_21.n8 a_79_21.t9 139.779
R224 a_79_21.n9 a_79_21.t11 139.779
R225 a_79_21.n3 a_79_21.t8 139.779
R226 a_79_21.n5 a_79_21.t13 139.779
R227 a_79_21.n2 a_79_21.n0 104.229
R228 a_79_21.n7 a_79_21.n6 101.6
R229 a_79_21.n2 a_79_21.n1 93.285
R230 a_79_21.n7 a_79_21.n4 76
R231 a_79_21.n11 a_79_21.n10 76
R232 a_79_21.n12 a_79_21.n2 73.331
R233 a_79_21.n13 a_79_21.t1 67.23
R234 a_79_21.n1 a_79_21.t0 64.285
R235 a_79_21.n6 a_79_21.n5 43.818
R236 a_79_21.n10 a_79_21.n8 40.896
R237 a_79_21.n1 a_79_21.t3 38.571
R238 a_79_21.n14 a_79_21.t2 38.24
R239 a_79_21.n4 a_79_21.n3 32.133
R240 a_79_21.n12 a_79_21.n11 28.235
R241 a_79_21.n11 a_79_21.n7 25.6
R242 a_79_21.n10 a_79_21.n9 20.448
R243 a_79_21.n14 a_79_21.n13 15.634
R244 a_79_21.n15 a_79_21.n14 3.338
R245 a_1271_47.n14 a_1271_47.n13 416.706
R246 a_1271_47.n13 a_1271_47.n0 222.095
R247 a_1271_47.n1 a_1271_47.t6 212.079
R248 a_1271_47.n3 a_1271_47.t11 212.079
R249 a_1271_47.n7 a_1271_47.t4 212.079
R250 a_1271_47.n10 a_1271_47.t5 212.079
R251 a_1271_47.n1 a_1271_47.t8 139.779
R252 a_1271_47.n3 a_1271_47.t9 139.779
R253 a_1271_47.n10 a_1271_47.t10 139.779
R254 a_1271_47.n6 a_1271_47.t7 139.779
R255 a_1271_47.n5 a_1271_47.n2 101.6
R256 a_1271_47.n5 a_1271_47.n4 76
R257 a_1271_47.n9 a_1271_47.n8 76
R258 a_1271_47.n12 a_1271_47.n11 76
R259 a_1271_47.n0 a_1271_47.t3 55.714
R260 a_1271_47.n0 a_1271_47.t0 55.714
R261 a_1271_47.t1 a_1271_47.n14 43.093
R262 a_1271_47.n14 a_1271_47.t2 41.554
R263 a_1271_47.n2 a_1271_47.n1 37.245
R264 a_1271_47.n9 a_1271_47.n5 25.6
R265 a_1271_47.n12 a_1271_47.n9 25.6
R266 a_1271_47.n4 a_1271_47.n3 25.56
R267 a_1271_47.n7 a_1271_47.n6 11.684
R268 a_1271_47.n11 a_1271_47.n10 9.493
R269 a_1271_47.n13 a_1271_47.n12 9.035
R270 a_1271_47.n8 a_1271_47.n7 2.19
R271 SUM.n2 SUM.n0 227.437
R272 SUM.n2 SUM.n1 109.186
R273 SUM.n5 SUM.n3 92.725
R274 SUM.n5 SUM.n4 52.431
R275 SUM.n3 SUM.t0 39.692
R276 SUM SUM.n2 30.903
R277 SUM SUM.n5 26.7
R278 SUM.n0 SUM.t7 26.595
R279 SUM.n0 SUM.t6 26.595
R280 SUM.n1 SUM.t5 26.595
R281 SUM.n1 SUM.t4 26.595
R282 SUM.n3 SUM.t3 24.923
R283 SUM.n4 SUM.t2 24.923
R284 SUM.n4 SUM.t1 24.923
R285 a_461_47.t0 a_461_47.t1 92.857
R286 COUT.n5 COUT.n4 223.615
R287 COUT.n3 COUT.n1 159.419
R288 COUT COUT.n0 156.262
R289 COUT.n3 COUT.n2 52.431
R290 COUT.n5 COUT.n3 36.914
R291 COUT.n0 COUT.t5 26.595
R292 COUT.n0 COUT.t4 26.595
R293 COUT.n4 COUT.t7 26.595
R294 COUT.n4 COUT.t6 26.595
R295 COUT.n1 COUT.t2 24.923
R296 COUT.n1 COUT.t1 24.923
R297 COUT.n2 COUT.t3 24.923
R298 COUT.n2 COUT.t0 24.923
R299 COUT COUT.n6 6.4
R300 COUT.n6 COUT.n5 4.654
R301 a_1014_47.n1 a_1014_47.n0 273.847
R302 a_1014_47.t0 a_1014_47.n1 45.714
R303 a_1014_47.n0 a_1014_47.t2 38.571
R304 a_1014_47.n0 a_1014_47.t1 38.571
R305 a_1014_47.n1 a_1014_47.t3 38.571
R306 a_1379_47.t0 a_1379_47.t1 60
R307 a_1451_47.t0 a_1451_47.t1 94.285
R308 a_1356_369.t1 a_1356_369.t0 96.234
R309 a_1451_371.t0 a_1451_371.t1 121.952
C0 VPB VPWR 0.20fF
C1 A CIN 0.47fF
C2 VGND SUM 0.40fF
C3 COUT VPWR 0.51fF
C4 B CIN 0.51fF
C5 COUT VGND 0.39fF
C6 VGND VPWR 0.13fF
C7 B VPWR 0.33fF
C8 A B 1.45fF
C9 SUM VPWR 0.47fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__fah_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__fah_1 COUT B A SUM CI VPWR VGND VNB VPB
X0 a_508_297.t0 B.t0 VGND.t0 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 a_1332_297.t0 a_719_47.t4 a_1262_49.t3 VNB.t5 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X2 a_27_47.t4 a_508_297.t4 a_719_47.t2 VNB.t10 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X3 VGND.t4 CI.t0 a_1262_49.t0 VNB.t8 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X4 a_67_199.t0 A.t0 VPWR.t6 VPB.t14 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 a_508_297.t1 B.t1 VPWR.t0 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 VPWR.t7 A.t1 a_310_49.t4 VPB.t13 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 a_310_49.t1 B.t2 a_1008_47.t1 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X8 a_508_297.t3 a_1008_47.t4 a_1332_297.t2 VNB.t11 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X9 a_1332_297.t1 a_719_47.t5 a_508_297.t2 VPB.t6 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X10 a_719_47.t1 B.t3 a_310_49.t0 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X11 a_1640_380.t2 a_719_47.t6 a_1617_49.t0 VNB.t6 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X12 a_1008_47.t3 a_508_297.t5 a_310_49.t3 VNB.t9 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X13 VGND.t3 a_1332_297.t4 COUT.t1 VNB.t7 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14 a_719_47.t0 B.t4 a_27_47.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X15 a_1262_49.t2 a_719_47.t7 a_1617_49.t1 VPB.t5 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X16 SUM.t0 a_1617_49.t4 VPWR.t1 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17 a_1640_380.t0 a_1262_49.t6 VPWR.t2 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X18 a_1617_49.t2 a_1008_47.t5 a_1640_380.t3 VPB.t11 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X19 VPWR.t4 a_1332_297.t5 COUT.t0 VPB.t7 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X20 VPWR.t3 a_67_199.t2 a_27_47.t2 VPB.t15 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X21 a_310_49.t2 a_508_297.t6 a_719_47.t3 VPB.t10 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X22 a_67_199.t1 A.t2 VGND.t6 VNB.t14 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X23 VGND.t7 A.t3 a_310_49.t5 VNB.t15 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X24 a_27_47.t1 B.t5 a_1008_47.t0 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X25 a_1617_49.t3 a_1008_47.t6 a_1262_49.t4 VNB.t12 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X26 a_1640_380.t1 a_1262_49.t7 VGND.t5 VNB.t13 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X27 SUM.t1 a_1617_49.t5 VGND.t1 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X28 VPWR.t5 CI.t1 a_1262_49.t1 VPB.t8 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X29 a_1008_47.t2 a_508_297.t7 a_27_47.t5 VPB.t9 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X30 VGND.t2 a_67_199.t3 a_27_47.t3 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X31 a_1262_49.t5 a_1008_47.t7 a_1332_297.t3 VPB.t12 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
R0 B.n3 B.t2 241.626
R1 B.n2 B.t1 212.079
R2 B.n0 B.t4 186.373
R3 B.n3 B.t5 154.81
R4 B.n0 B.t3 141.386
R5 B.n1 B.t0 139.779
R6 B.n1 B.n0 139.487
R7 B.n4 B.n2 112.038
R8 B.n2 B.n1 14.606
R9 B B.n3 13.196
R10 B B.n4 5.44
R11 B.n4 B 4.65
R12 VGND.n3 VGND.n2 116.217
R13 VGND.n39 VGND.n38 114.711
R14 VGND.n47 VGND.n46 114.711
R15 VGND.n1 VGND.n0 68.138
R16 VGND.n38 VGND.t0 67.041
R17 VGND.n46 VGND.t6 35.625
R18 VGND.n2 VGND.t5 25.312
R19 VGND.n2 VGND.t4 25.312
R20 VGND.n38 VGND.t7 25.312
R21 VGND.n0 VGND.t1 24.923
R22 VGND.n0 VGND.t3 24.923
R23 VGND.n46 VGND.t2 22.167
R24 VGND.n4 VGND.n3 7.529
R25 VGND.n5 VGND.n4 4.65
R26 VGND.n7 VGND.n6 4.65
R27 VGND.n9 VGND.n8 4.65
R28 VGND.n11 VGND.n10 4.65
R29 VGND.n13 VGND.n12 4.65
R30 VGND.n15 VGND.n14 4.65
R31 VGND.n17 VGND.n16 4.65
R32 VGND.n19 VGND.n18 4.65
R33 VGND.n21 VGND.n20 4.65
R34 VGND.n23 VGND.n22 4.65
R35 VGND.n25 VGND.n24 4.65
R36 VGND.n27 VGND.n26 4.65
R37 VGND.n29 VGND.n28 4.65
R38 VGND.n31 VGND.n30 4.65
R39 VGND.n33 VGND.n32 4.65
R40 VGND.n35 VGND.n34 4.65
R41 VGND.n37 VGND.n36 4.65
R42 VGND.n41 VGND.n40 4.65
R43 VGND.n43 VGND.n42 4.65
R44 VGND.n45 VGND.n44 4.65
R45 VGND.n49 VGND.n48 4.65
R46 VGND.n40 VGND.n39 1.882
R47 VGND.n48 VGND.n47 0.752
R48 VGND.n5 VGND.n1 0.143
R49 VGND.n7 VGND.n5 0.119
R50 VGND.n9 VGND.n7 0.119
R51 VGND.n11 VGND.n9 0.119
R52 VGND.n13 VGND.n11 0.119
R53 VGND.n15 VGND.n13 0.119
R54 VGND.n17 VGND.n15 0.119
R55 VGND.n19 VGND.n17 0.119
R56 VGND.n21 VGND.n19 0.119
R57 VGND.n23 VGND.n21 0.119
R58 VGND.n25 VGND.n23 0.119
R59 VGND.n27 VGND.n25 0.119
R60 VGND.n29 VGND.n27 0.119
R61 VGND.n31 VGND.n29 0.119
R62 VGND.n33 VGND.n31 0.119
R63 VGND.n35 VGND.n33 0.119
R64 VGND.n37 VGND.n35 0.119
R65 VGND.n41 VGND.n37 0.119
R66 VGND.n43 VGND.n41 0.119
R67 VGND.n45 VGND.n43 0.119
R68 VGND.n49 VGND.n45 0.119
R69 VGND.n50 VGND.n49 0.119
R70 VGND VGND.n50 0.022
R71 a_508_297.n2 a_508_297.t3 310.11
R72 a_508_297.t1 a_508_297.n9 255.427
R73 a_508_297.n2 a_508_297.t2 213.063
R74 a_508_297.n3 a_508_297.t7 191.485
R75 a_508_297.n4 a_508_297.t6 186.373
R76 a_508_297.n0 a_508_297.t0 175.982
R77 a_508_297.n4 a_508_297.t4 141.386
R78 a_508_297.n3 a_508_297.t5 141.386
R79 a_508_297.n5 a_508_297.n3 106.624
R80 a_508_297.n6 a_508_297.n5 90.834
R81 a_508_297.n9 a_508_297.n8 50.85
R82 a_508_297.n5 a_508_297.n4 42.357
R83 a_508_297.n8 a_508_297.n7 9.3
R84 a_508_297.n6 a_508_297.n2 7.117
R85 a_508_297.n7 a_508_297.n6 5.405
R86 a_508_297.n7 a_508_297.n1 3.318
R87 a_508_297.n1 a_508_297.n0 0.711
R88 VNB.t6 VNB.t8 6502.22
R89 VNB VNB.t4 6078.09
R90 VNB.t13 VNB.t7 6012.26
R91 VNB.t10 VNB.t9 4986.67
R92 VNB.t2 VNB.t1 4642.83
R93 VNB.t11 VNB.t12 4595.56
R94 VNB.t0 VNB.t5 4595.56
R95 VNB.t14 VNB.t15 4545.05
R96 VNB.t9 VNB.t0 3594.41
R97 VNB.t15 VNB.t2 3287.91
R98 VNB.t4 VNB.t14 2296.7
R99 VNB.t12 VNB.t6 2151.11
R100 VNB.t5 VNB.t11 2077.78
R101 VNB.t1 VNB.t10 2077.78
R102 VNB.t8 VNB.t13 2053.33
R103 VNB.t7 VNB.t3 2030.77
R104 a_719_47.n5 a_719_47.n4 348.718
R105 a_719_47.n0 a_719_47.t6 289.199
R106 a_719_47.n0 a_719_47.t7 284.38
R107 a_719_47.n1 a_719_47.t5 186.373
R108 a_719_47.n1 a_719_47.t4 146.935
R109 a_719_47.n2 a_719_47.n1 138.683
R110 a_719_47.n4 a_719_47.n3 116.97
R111 a_719_47.n2 a_719_47.n0 73.072
R112 a_719_47.n5 a_719_47.t3 32.833
R113 a_719_47.t0 a_719_47.n5 31.66
R114 a_719_47.n3 a_719_47.t1 26.25
R115 a_719_47.n3 a_719_47.t2 25.312
R116 a_719_47.n4 a_719_47.n2 7.029
R117 a_1262_49.n5 a_1262_49.t5 464.875
R118 a_1262_49.n2 a_1262_49.n1 294.621
R119 a_1262_49.n7 a_1262_49.n6 292.5
R120 a_1262_49.n0 a_1262_49.t6 238.154
R121 a_1262_49.n3 a_1262_49.t0 234.604
R122 a_1262_49.n3 a_1262_49.t3 207.716
R123 a_1262_49.n0 a_1262_49.t7 164.247
R124 a_1262_49.n6 a_1262_49.n5 146.904
R125 a_1262_49.n1 a_1262_49.n0 139.492
R126 a_1262_49.n4 a_1262_49.t4 117.812
R127 a_1262_49.n7 a_1262_49.t2 84.428
R128 a_1262_49.n5 a_1262_49.n4 69.04
R129 a_1262_49.n2 a_1262_49.t1 25.45
R130 a_1262_49.n9 a_1262_49.n8 24.625
R131 a_1262_49.n10 a_1262_49.n9 21.621
R132 a_1262_49.n4 a_1262_49.n3 16.062
R133 a_1262_49.n9 a_1262_49.n2 13.196
R134 a_1262_49.n8 a_1262_49.n7 4.69
R135 a_1332_297.n3 a_1332_297.n2 322.505
R136 a_1332_297.n0 a_1332_297.t5 232.247
R137 a_1332_297.n0 a_1332_297.t4 161.878
R138 a_1332_297.n2 a_1332_297.n1 111.462
R139 a_1332_297.n3 a_1332_297.t3 31.66
R140 a_1332_297.t1 a_1332_297.n3 31.66
R141 a_1332_297.n1 a_1332_297.t2 26.25
R142 a_1332_297.n1 a_1332_297.t0 25.312
R143 a_1332_297.n2 a_1332_297.n0 18.534
R144 a_27_47.n12 a_27_47.t0 560.35
R145 a_27_47.n11 a_27_47.t5 247.164
R146 a_27_47.n13 a_27_47.n12 231.46
R147 a_27_47.n0 a_27_47.t1 198.987
R148 a_27_47.n10 a_27_47.t4 174.158
R149 a_27_47.n13 a_27_47.t3 156.146
R150 a_27_47.n12 a_27_47.n11 142.164
R151 a_27_47.t2 a_27_47.n13 122.686
R152 a_27_47.n8 a_27_47.n7 98.986
R153 a_27_47.n2 a_27_47.n0 80.082
R154 a_27_47.n11 a_27_47.n10 75.654
R155 a_27_47.n6 a_27_47.n5 54.4
R156 a_27_47.n4 a_27_47.n3 38.4
R157 a_27_47.n2 a_27_47.n1 25.6
R158 a_27_47.n9 a_27_47.n8 19.536
R159 a_27_47.n10 a_27_47.n9 18.248
R160 a_27_47.n9 a_27_47.n6 9.6
R161 a_27_47.n6 a_27_47.n4 5.12
R162 a_27_47.n4 a_27_47.n2 1.828
R163 CI.n0 CI.t1 233.868
R164 CI.n0 CI.t0 159.961
R165 CI CI.n0 99.952
R166 A.n0 A.t1 214.269
R167 A.n1 A.t0 212.809
R168 A.n1 A.t2 141.386
R169 A.n0 A.t3 138.172
R170 A.n2 A.n0 103.703
R171 A A.n2 83.04
R172 A.n2 A.n1 33.593
R173 VPWR.n37 VPWR.n36 308.015
R174 VPWR.n1 VPWR.n0 306.255
R175 VPWR.n44 VPWR.n43 305.65
R176 VPWR.n3 VPWR.n2 175.92
R177 VPWR.n36 VPWR.t7 50.235
R178 VPWR.n43 VPWR.t3 32.505
R179 VPWR.n36 VPWR.t0 31.52
R180 VPWR.n2 VPWR.t1 26.595
R181 VPWR.n2 VPWR.t4 26.595
R182 VPWR.n0 VPWR.t2 26.595
R183 VPWR.n0 VPWR.t5 26.595
R184 VPWR.n43 VPWR.t6 26.595
R185 VPWR.n5 VPWR.n4 4.65
R186 VPWR.n7 VPWR.n6 4.65
R187 VPWR.n9 VPWR.n8 4.65
R188 VPWR.n11 VPWR.n10 4.65
R189 VPWR.n13 VPWR.n12 4.65
R190 VPWR.n15 VPWR.n14 4.65
R191 VPWR.n17 VPWR.n16 4.65
R192 VPWR.n19 VPWR.n18 4.65
R193 VPWR.n21 VPWR.n20 4.65
R194 VPWR.n23 VPWR.n22 4.65
R195 VPWR.n25 VPWR.n24 4.65
R196 VPWR.n27 VPWR.n26 4.65
R197 VPWR.n29 VPWR.n28 4.65
R198 VPWR.n31 VPWR.n30 4.65
R199 VPWR.n33 VPWR.n32 4.65
R200 VPWR.n35 VPWR.n34 4.65
R201 VPWR.n38 VPWR.n37 4.65
R202 VPWR.n40 VPWR.n39 4.65
R203 VPWR.n42 VPWR.n41 4.65
R204 VPWR.n45 VPWR.n44 4.01
R205 VPWR.n3 VPWR.n1 3.642
R206 VPWR.n5 VPWR.n3 0.149
R207 VPWR.n45 VPWR.n42 0.135
R208 VPWR VPWR.n45 0.125
R209 VPWR.n7 VPWR.n5 0.119
R210 VPWR.n9 VPWR.n7 0.119
R211 VPWR.n11 VPWR.n9 0.119
R212 VPWR.n13 VPWR.n11 0.119
R213 VPWR.n15 VPWR.n13 0.119
R214 VPWR.n17 VPWR.n15 0.119
R215 VPWR.n19 VPWR.n17 0.119
R216 VPWR.n21 VPWR.n19 0.119
R217 VPWR.n23 VPWR.n21 0.119
R218 VPWR.n25 VPWR.n23 0.119
R219 VPWR.n27 VPWR.n25 0.119
R220 VPWR.n29 VPWR.n27 0.119
R221 VPWR.n31 VPWR.n29 0.119
R222 VPWR.n33 VPWR.n31 0.119
R223 VPWR.n35 VPWR.n33 0.119
R224 VPWR.n38 VPWR.n35 0.119
R225 VPWR.n40 VPWR.n38 0.119
R226 VPWR.n42 VPWR.n40 0.119
R227 a_67_199.t0 a_67_199.n1 601.052
R228 a_67_199.n0 a_67_199.t2 236.932
R229 a_67_199.n0 a_67_199.t3 164.632
R230 a_67_199.n1 a_67_199.t1 126.301
R231 a_67_199.n1 a_67_199.n0 76
R232 VPB.t12 VPB.t11 905.607
R233 VPB.t4 VPB.t7 722.118
R234 VPB.t1 VPB.t6 651.09
R235 VPB.t10 VPB.t9 624.454
R236 VPB.t2 VPB.t0 624.454
R237 VPB.t14 VPB.t13 568.224
R238 VPB.t5 VPB.t8 497.196
R239 VPB.t13 VPB.t2 334.423
R240 VPB.t9 VPB.t1 287.071
R241 VPB.t15 VPB.t14 266.355
R242 VPB.t0 VPB.t10 251.557
R243 VPB.t7 VPB.t3 248.598
R244 VPB.t8 VPB.t4 248.598
R245 VPB.t11 VPB.t5 248.598
R246 VPB.t6 VPB.t12 248.598
R247 VPB VPB.t15 204.205
R248 a_310_49.t4 a_310_49.n3 619.325
R249 a_310_49.n0 a_310_49.t2 327.36
R250 a_310_49.n1 a_310_49.t3 205.887
R251 a_310_49.n2 a_310_49.n0 180.893
R252 a_310_49.n0 a_310_49.t1 142.716
R253 a_310_49.n1 a_310_49.t0 120.147
R254 a_310_49.n3 a_310_49.n2 116.615
R255 a_310_49.n3 a_310_49.t5 91.103
R256 a_310_49.n2 a_310_49.n1 11.885
R257 a_1008_47.n4 a_1008_47.n2 340.852
R258 a_1008_47.n0 a_1008_47.t5 319.032
R259 a_1008_47.n5 a_1008_47.n4 292.5
R260 a_1008_47.n4 a_1008_47.n3 196.48
R261 a_1008_47.n1 a_1008_47.t7 195.866
R262 a_1008_47.n1 a_1008_47.t4 138.172
R263 a_1008_47.n0 a_1008_47.t6 138.172
R264 a_1008_47.n2 a_1008_47.n0 69.378
R265 a_1008_47.n2 a_1008_47.n1 67.918
R266 a_1008_47.n3 a_1008_47.t3 66.127
R267 a_1008_47.t1 a_1008_47.n5 50.157
R268 a_1008_47.n5 a_1008_47.t2 32.248
R269 a_1008_47.n3 a_1008_47.t0 26.063
R270 a_1617_49.n3 a_1617_49.n2 300.029
R271 a_1617_49.n0 a_1617_49.t4 241.534
R272 a_1617_49.n0 a_1617_49.t5 169.234
R273 a_1617_49.n2 a_1617_49.n1 146.583
R274 a_1617_49.n2 a_1617_49.n0 103.349
R275 a_1617_49.t1 a_1617_49.n3 31.66
R276 a_1617_49.n3 a_1617_49.t2 31.66
R277 a_1617_49.n1 a_1617_49.t3 29.062
R278 a_1617_49.n1 a_1617_49.t0 25.312
R279 a_1640_380.n0 a_1640_380.t3 395.287
R280 a_1640_380.t0 a_1640_380.n1 327.69
R281 a_1640_380.n0 a_1640_380.t2 284.87
R282 a_1640_380.n1 a_1640_380.t1 169.033
R283 a_1640_380.n1 a_1640_380.n0 10.482
R284 COUT.n1 COUT.n0 292.5
R285 COUT.n0 COUT.t1 179.316
R286 COUT.n2 COUT.n1 146.493
R287 COUT.n1 COUT.t0 26.595
R288 COUT.n2 COUT 6.496
R289 COUT.n0 COUT 3.692
R290  COUT.n2 1.85
R291 SUM.n2 SUM.t0 173.92
R292  SUM.n0 93.761
R293 SUM.n1 SUM.n0 92.5
R294 SUM.n0 SUM.t1 39.692
R295 SUM  19.342
R296 SUM.n3 SUM 15.928
R297 SUM.n1  10.997
R298  SUM.n2 9.355
R299  SUM.n3 3.413
R300 SUM.n2  3.019
R301 SUM.n3  2.163
R302  SUM.n1 1.261
C0 VPWR VPB 0.25fF
C1 VGND SUM 0.16fF
C2 VPWR COUT 0.16fF
C3 VPWR SUM 0.17fF
C4 VGND COUT 0.16fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__fahcin_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__fahcin_1 COUT B A SUM CIN VPWR VGND VNB VPB
X0 a_721_47.t2 a_489_21.t2 a_27_47.t2 VPB.t5 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X1 VGND.t1 a_1636_315.t4 a_1565_49.t0 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X2 SUM.t1 a_1647_49.t4 VPWR.t1 VPB.t10 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 VGND.t2 CIN.t0 a_1251_49.t1 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X4 VPWR.t4 a_67_199.t6 a_27_47.t3 VPB.t7 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 a_67_199.t4 B.t0 a_721_47.t3 VPB.t13 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X6 VPWR.t2 CIN.t1 a_1251_49.t2 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 a_67_199.t1 a_489_21.t3 a_434_49.t0 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X8 COUT.t1 a_434_49.t4 a_1251_49.t0 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X9 a_1647_49.t3 a_721_47.t4 a_1565_49.t3 VNB.t13 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X10 a_434_49.t2 B.t1 a_67_199.t5 VNB.t14 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X11 a_434_49.t3 B.t2 a_27_47.t5 VPB.t14 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X12 VPWR.t0 a_1636_315.t5 a_1565_49.t1 VPB.t6 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13 VGND.t7 B.t3 a_489_21.t0 VNB.t15 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14 SUM.t0 a_1647_49.t5 VGND.t6 VNB.t11 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X15 a_67_199.t3 A.t0 VPWR.t6 VPB.t9 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16 a_1142_49.t3 a_721_47.t5 COUT.t2 VNB.t12 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X17 VGND.t4 a_67_199.t7 a_27_47.t4 VNB.t9 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X18 a_27_47.t1 a_489_21.t4 a_434_49.t1 VNB.t8 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X19 a_67_199.t0 A.t1 VGND.t0 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X20 VPWR.t7 B.t4 a_489_21.t1 VPB.t15 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X21 a_27_47.t0 B.t5 a_721_47.t0 VNB.t5 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X22 a_1251_49.t3 a_721_47.t6 COUT.t3 VPB.t12 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X23 a_1142_49.t0 a_489_21.t5 VGND.t3 VNB.t7 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X24 a_1142_49.t1 a_489_21.t6 VPWR.t3 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X25 a_1565_49.t2 a_434_49.t5 a_1647_49.t0 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X26 a_721_47.t1 a_489_21.t7 a_67_199.t2 VNB.t6 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X27 a_1636_315.t0 a_434_49.t6 a_1647_49.t1 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X28 a_1647_49.t2 a_721_47.t7 a_1636_315.t3 VPB.t11 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X29 a_1636_315.t1 CIN.t2 VPWR.t5 VPB.t8 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X30 COUT.t0 a_434_49.t7 a_1142_49.t2 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X31 a_1636_315.t2 CIN.t3 VGND.t5 VNB.t10 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
R0 a_489_21.t1 a_489_21.n5 301.63
R1 a_489_21.n3 a_489_21.t6 238.589
R2 a_489_21.n0 a_489_21.t2 194.406
R3 a_489_21.n1 a_489_21.t3 186.373
R4 a_489_21.n3 a_489_21.t5 164.682
R5 a_489_21.n4 a_489_21.t0 161.414
R6 a_489_21.n0 a_489_21.t7 141.386
R7 a_489_21.n1 a_489_21.t4 138.172
R8 a_489_21.n5 a_489_21.n2 120.777
R9 a_489_21.n2 a_489_21.n0 105.893
R10 a_489_21.n4 a_489_21.n3 90.545
R11 a_489_21.n2 a_489_21.n1 41.627
R12 a_489_21.n5 a_489_21.n4 12.675
R13 a_27_47.n2 a_27_47.t5 452.585
R14 a_27_47.n1 a_27_47.t2 241.787
R15 a_27_47.n0 a_27_47.t0 219.798
R16 a_27_47.n3 a_27_47.t4 169.635
R17 a_27_47.n0 a_27_47.t1 166.13
R18 a_27_47.n2 a_27_47.n1 132.581
R19 a_27_47.t3 a_27_47.n3 123.83
R20 a_27_47.n3 a_27_47.n2 119.578
R21 a_27_47.n1 a_27_47.n0 74.577
R22 a_721_47.n4 a_721_47.n2 504.943
R23 a_721_47.n5 a_721_47.n4 292.5
R24 a_721_47.n0 a_721_47.t7 282.084
R25 a_721_47.n1 a_721_47.t6 195.136
R26 a_721_47.n4 a_721_47.n3 187.636
R27 a_721_47.n0 a_721_47.t4 144.744
R28 a_721_47.n1 a_721_47.t5 138.172
R29 a_721_47.n2 a_721_47.n1 130.724
R30 a_721_47.n3 a_721_47.t1 62.592
R31 a_721_47.n5 a_721_47.t3 50.157
R32 a_721_47.t2 a_721_47.n5 32.248
R33 a_721_47.n2 a_721_47.n0 24.1
R34 a_721_47.n3 a_721_47.t0 20.109
R35 VPB.t12 VPB.t11 899.688
R36 VPB.t1 VPB.t6 668.847
R37 VPB.t9 VPB.t14 662.928
R38 VPB.t4 VPB.t5 630.373
R39 VPB.t13 VPB.t15 624.454
R40 VPB.t8 VPB.t0 571.183
R41 VPB.t3 VPB.t2 556.386
R42 VPB.t15 VPB.t3 301.869
R43 VPB.t7 VPB.t9 295.95
R44 VPB.t5 VPB.t13 287.071
R45 VPB.t14 VPB.t4 251.557
R46 VPB.t0 VPB.t10 248.598
R47 VPB.t6 VPB.t8 248.598
R48 VPB.t11 VPB.t1 248.598
R49 VPB.t2 VPB.t12 248.598
R50 VPB VPB.t7 195.327
R51 a_1636_315.n2 a_1636_315.t3 432.959
R52 a_1636_315.n0 a_1636_315.t5 241.534
R53 a_1636_315.n2 a_1636_315.t0 198.302
R54 a_1636_315.n0 a_1636_315.t4 167.627
R55 a_1636_315.t1 a_1636_315.n3 125.311
R56 a_1636_315.n1 a_1636_315.t2 123.471
R57 a_1636_315.n1 a_1636_315.n0 76
R58 a_1636_315.n3 a_1636_315.n2 72.604
R59 a_1636_315.n3 a_1636_315.n1 21.778
R60 a_1565_49.n1 a_1565_49.n0 369.458
R61 a_1565_49.n0 a_1565_49.t3 260.93
R62 a_1565_49.n2 a_1565_49.t2 174.72
R63 a_1565_49.n0 a_1565_49.t0 80.931
R64 a_1565_49.n1 a_1565_49.t1 20.908
R65 a_1565_49.n3 a_1565_49.n2 18.861
R66 a_1565_49.n2 a_1565_49.n1 12.978
R67 VGND.n2 VGND.n1 116.217
R68 VGND.n46 VGND.n45 114.711
R69 VGND.n3 VGND.n0 111.331
R70 VGND.n25 VGND.n24 64.067
R71 VGND.n24 VGND.t3 40.312
R72 VGND.n0 VGND.t6 32.479
R73 VGND.n45 VGND.t4 30.937
R74 VGND.n1 VGND.t1 29.062
R75 VGND.n1 VGND.t5 28.729
R76 VGND.n45 VGND.t0 26.854
R77 VGND.n0 VGND.t2 25.312
R78 VGND.n24 VGND.t7 24.042
R79 VGND.n3 VGND.n2 10.531
R80 VGND.n47 VGND.n46 6.029
R81 VGND.n5 VGND.n4 4.65
R82 VGND.n7 VGND.n6 4.65
R83 VGND.n9 VGND.n8 4.65
R84 VGND.n11 VGND.n10 4.65
R85 VGND.n13 VGND.n12 4.65
R86 VGND.n15 VGND.n14 4.65
R87 VGND.n17 VGND.n16 4.65
R88 VGND.n19 VGND.n18 4.65
R89 VGND.n21 VGND.n20 4.65
R90 VGND.n23 VGND.n22 4.65
R91 VGND.n26 VGND.n25 4.65
R92 VGND.n28 VGND.n27 4.65
R93 VGND.n30 VGND.n29 4.65
R94 VGND.n32 VGND.n31 4.65
R95 VGND.n34 VGND.n33 4.65
R96 VGND.n36 VGND.n35 4.65
R97 VGND.n38 VGND.n37 4.65
R98 VGND.n40 VGND.n39 4.65
R99 VGND.n42 VGND.n41 4.65
R100 VGND.n44 VGND.n43 4.65
R101 VGND.n5 VGND.n3 0.142
R102 VGND.n47 VGND.n44 0.132
R103 VGND VGND.n47 0.129
R104 VGND.n7 VGND.n5 0.119
R105 VGND.n9 VGND.n7 0.119
R106 VGND.n11 VGND.n9 0.119
R107 VGND.n13 VGND.n11 0.119
R108 VGND.n15 VGND.n13 0.119
R109 VGND.n17 VGND.n15 0.119
R110 VGND.n19 VGND.n17 0.119
R111 VGND.n21 VGND.n19 0.119
R112 VGND.n23 VGND.n21 0.119
R113 VGND.n26 VGND.n23 0.119
R114 VGND.n28 VGND.n26 0.119
R115 VGND.n30 VGND.n28 0.119
R116 VGND.n32 VGND.n30 0.119
R117 VGND.n34 VGND.n32 0.119
R118 VGND.n36 VGND.n34 0.119
R119 VGND.n38 VGND.n36 0.119
R120 VGND.n40 VGND.n38 0.119
R121 VGND.n42 VGND.n40 0.119
R122 VGND.n44 VGND.n42 0.119
R123 VNB.t4 VNB.t1 7015.56
R124 VNB VNB.t9 6115.42
R125 VNB.t0 VNB.t14 5556.41
R126 VNB.t12 VNB.t13 5402.22
R127 VNB.t8 VNB.t6 4911.99
R128 VNB.t7 VNB.t3 4864.44
R129 VNB.t10 VNB.t2 4545.05
R130 VNB.t5 VNB.t15 4496.7
R131 VNB.t6 VNB.t5 3215.38
R132 VNB.t15 VNB.t7 2333.7
R133 VNB.t2 VNB.t11 2296.7
R134 VNB.t1 VNB.t10 2248.62
R135 VNB.t9 VNB.t0 2248.62
R136 VNB.t13 VNB.t4 2151.11
R137 VNB.t3 VNB.t12 2077.78
R138 VNB.t14 VNB.t8 2077.78
R139 a_1647_49.n1 a_1647_49.t4 241.534
R140 a_1647_49.n1 a_1647_49.t5 169.234
R141 a_1647_49.n3 a_1647_49.n2 153.417
R142 a_1647_49.n2 a_1647_49.n0 141.613
R143 a_1647_49.n2 a_1647_49.n1 103.366
R144 a_1647_49.t0 a_1647_49.n3 31.66
R145 a_1647_49.n3 a_1647_49.t2 31.66
R146 a_1647_49.n0 a_1647_49.t3 29.062
R147 a_1647_49.n0 a_1647_49.t1 25.312
R148 VPWR.n46 VPWR.n45 314.335
R149 VPWR.n1 VPWR.n0 313.205
R150 VPWR.n25 VPWR.n24 308.015
R151 VPWR.n3 VPWR.n2 175.818
R152 VPWR.n24 VPWR.t7 44.325
R153 VPWR.n45 VPWR.t6 42.355
R154 VPWR.n2 VPWR.t1 26.595
R155 VPWR.n2 VPWR.t2 26.595
R156 VPWR.n0 VPWR.t5 26.595
R157 VPWR.n0 VPWR.t0 26.595
R158 VPWR.n24 VPWR.t3 26.595
R159 VPWR.n45 VPWR.t4 26.595
R160 VPWR.n3 VPWR.n1 9.78
R161 VPWR.n48 VPWR.n47 4.65
R162 VPWR.n5 VPWR.n4 4.65
R163 VPWR.n7 VPWR.n6 4.65
R164 VPWR.n9 VPWR.n8 4.65
R165 VPWR.n11 VPWR.n10 4.65
R166 VPWR.n13 VPWR.n12 4.65
R167 VPWR.n15 VPWR.n14 4.65
R168 VPWR.n17 VPWR.n16 4.65
R169 VPWR.n19 VPWR.n18 4.65
R170 VPWR.n21 VPWR.n20 4.65
R171 VPWR.n23 VPWR.n22 4.65
R172 VPWR.n26 VPWR.n25 4.65
R173 VPWR.n28 VPWR.n27 4.65
R174 VPWR.n30 VPWR.n29 4.65
R175 VPWR.n32 VPWR.n31 4.65
R176 VPWR.n34 VPWR.n33 4.65
R177 VPWR.n36 VPWR.n35 4.65
R178 VPWR.n38 VPWR.n37 4.65
R179 VPWR.n40 VPWR.n39 4.65
R180 VPWR.n42 VPWR.n41 4.65
R181 VPWR.n44 VPWR.n43 4.65
R182 VPWR.n47 VPWR.n46 0.376
R183 VPWR.n5 VPWR.n3 0.141
R184 VPWR.n7 VPWR.n5 0.119
R185 VPWR.n9 VPWR.n7 0.119
R186 VPWR.n11 VPWR.n9 0.119
R187 VPWR.n13 VPWR.n11 0.119
R188 VPWR.n15 VPWR.n13 0.119
R189 VPWR.n17 VPWR.n15 0.119
R190 VPWR.n19 VPWR.n17 0.119
R191 VPWR.n21 VPWR.n19 0.119
R192 VPWR.n23 VPWR.n21 0.119
R193 VPWR.n26 VPWR.n23 0.119
R194 VPWR.n28 VPWR.n26 0.119
R195 VPWR.n30 VPWR.n28 0.119
R196 VPWR.n32 VPWR.n30 0.119
R197 VPWR.n34 VPWR.n32 0.119
R198 VPWR.n36 VPWR.n34 0.119
R199 VPWR.n38 VPWR.n36 0.119
R200 VPWR.n40 VPWR.n38 0.119
R201 VPWR.n42 VPWR.n40 0.119
R202 VPWR.n44 VPWR.n42 0.119
R203 VPWR.n48 VPWR.n44 0.119
R204 VPWR.n49 VPWR.n48 0.119
R205 VPWR VPWR.n49 0.022
R206 SUM.n1 SUM.t1 173.924
R207 SUM.n0 SUM.t0 79.594
R208 SUM  20.723
R209 SUM.n2 SUM 17.066
R210  SUM.n1 9.77
R211  SUM.n0 6.843
R212 SUM.n0  5.57
R213  SUM.n2 3.657
R214 SUM.n1  3.155
R215 SUM.n2  2.258
R216 CIN.n1 CIN.t2 215.73
R217 CIN.n0 CIN.t1 212.079
R218 CIN.n1 CIN.t3 139.779
R219 CIN.n0 CIN.t0 138.172
R220 CIN.n2 CIN.n0 100.051
R221 CIN CIN.n2 77.582
R222 CIN.n2 CIN.n1 37.245
R223 a_1251_49.n0 a_1251_49.t3 294.462
R224 a_1251_49.n0 a_1251_49.t0 232.218
R225 a_1251_49.t2 a_1251_49.n1 169.084
R226 a_1251_49.n1 a_1251_49.t1 136.304
R227 a_1251_49.n1 a_1251_49.n0 12.5
R228 a_67_199.t3 a_67_199.n7 407.384
R229 a_67_199.n1 a_67_199.t6 236.179
R230 a_67_199.n4 a_67_199.t2 217.669
R231 a_67_199.n1 a_67_199.t7 165.486
R232 a_67_199.n8 a_67_199.t3 126.08
R233 a_67_199.n4 a_67_199.n3 92.5
R234 a_67_199.n6 a_67_199.n1 76
R235 a_67_199.n7 a_67_199.n6 69.572
R236 a_67_199.n7 a_67_199.n0 59
R237 a_67_199.n5 a_67_199.n2 48.937
R238 a_67_199.n6 a_67_199.n5 45.347
R239 a_67_199.n5 a_67_199.n4 41.064
R240 a_67_199.n0 a_67_199.t4 37.621
R241 a_67_199.n0 a_67_199.t1 34.448
R242 a_67_199.n3 a_67_199.t5 25.312
R243 a_67_199.n2 a_67_199.t0 14.183
R244 B.n2 B.t0 244.797
R245 B.n1 B.t4 212.079
R246 B.n0 B.t2 186.373
R247 B.n4 B.n0 157.518
R248 B.n1 B.t3 139.779
R249 B.n0 B.t1 138.172
R250 B.n2 B.t5 138.172
R251 B.n3 B.n1 116.848
R252 B B.n3 98.883
R253 B.n3 B.n2 18.987
R254 B B.n4 4.73
R255 B.n4 B 4.65
R256 a_434_49.n5 a_434_49.n4 317.885
R257 a_434_49.n1 a_434_49.t5 244.519
R258 a_434_49.n1 a_434_49.t6 215.312
R259 a_434_49.n0 a_434_49.t7 186.373
R260 a_434_49.n0 a_434_49.t4 146.205
R261 a_434_49.n4 a_434_49.n3 106.09
R262 a_434_49.n2 a_434_49.n0 50.036
R263 a_434_49.t0 a_434_49.n5 32.833
R264 a_434_49.n5 a_434_49.t3 31.66
R265 a_434_49.n3 a_434_49.t1 26.25
R266 a_434_49.n3 a_434_49.t2 25.312
R267 a_434_49.n2 a_434_49.n1 12.359
R268 a_434_49.n4 a_434_49.n2 8.263
R269 COUT COUT.n1 300.796
R270 COUT.n2 COUT.n0 100.405
R271 COUT.n1 COUT.t3 31.66
R272 COUT.n1 COUT.t0 31.66
R273 COUT.n0 COUT.t2 26.25
R274 COUT.n0 COUT.t1 25.312
R275 COUT.n2 COUT 24.651
R276 COUT.n2  10.164
R277  COUT.n2 7.585
R278 A.n0 A.t0 230.361
R279 A.n0 A.t1 158.061
R280 A A.n0 83.04
R281 a_1142_49.n0 a_1142_49.t3 312.713
R282 a_1142_49.n3 a_1142_49.n2 302.963
R283 a_1142_49.n1 a_1142_49.n0 292.5
R284 a_1142_49.n2 a_1142_49.t0 183.901
R285 a_1142_49.n4 a_1142_49.n1 79.738
R286 a_1142_49.n1 a_1142_49.t2 31.66
R287 a_1142_49.n4 a_1142_49.n3 24.827
R288 a_1142_49.n5 a_1142_49.n4 24.818
R289 a_1142_49.n3 a_1142_49.t1 18.62
C0 VPWR SUM 0.17fF
C1 VPB VPWR 0.25fF
C2 SUM VGND 0.10fF
C3 B VGND 0.26fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__fahcon_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__fahcon_1 COUT_N B A SUM CI VPWR VGND VNB VPB
X0 a_1144_49.t2 B.t0 VPWR.t4 VPB.t13 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 VPWR.t6 a_67_199.t6 a_28_47.t4 VPB.t14 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 VGND.t5 B.t1 a_488_21.t1 VNB.t13 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 COUT_N.t1 a_434_49.t4 a_1261_49.t0 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X4 a_1589_49.t0 a_434_49.t5 a_1710_49.t1 VPB.t5 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X5 SUM.t1 a_1710_49.t4 VGND.t3 VNB.t7 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 a_1710_49.t2 a_726_47.t4 a_1634_315.t3 VPB.t8 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X7 a_434_49.t3 B.t2 a_67_199.t4 VNB.t12 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X8 a_434_49.t2 B.t3 a_28_47.t3 VPB.t12 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X9 a_1589_49.t2 CI.t0 VPWR.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 COUT_N.t0 a_434_49.t6 a_1144_49.t0 VPB.t6 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X11 a_1144_49.t1 a_726_47.t5 COUT_N.t2 VNB.t8 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X12 SUM.t0 a_1710_49.t5 VPWR.t3 VPB.t7 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13 a_67_199.t0 A.t0 VPWR.t2 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14 a_28_47.t2 B.t4 a_726_47.t2 VNB.t11 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X15 VPWR.t1 CI.t1 a_1261_49.t2 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16 VGND.t7 a_67_199.t7 a_28_47.t5 VNB.t15 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X17 a_28_47.t0 a_488_21.t2 a_434_49.t0 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X18 a_1144_49.t3 B.t5 VGND.t4 VNB.t10 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X19 a_726_47.t0 a_488_21.t3 a_28_47.t1 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X20 a_67_199.t3 A.t1 VGND.t2 VNB.t6 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X21 VPWR.t7 a_1589_49.t4 a_1634_315.t1 VPB.t15 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X22 a_726_47.t1 a_488_21.t4 a_67_199.t1 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X23 a_1710_49.t3 a_726_47.t6 a_1589_49.t3 VNB.t9 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X24 a_1634_315.t0 a_434_49.t7 a_1710_49.t0 VNB.t5 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X25 a_67_199.t5 B.t6 a_726_47.t3 VPB.t11 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X26 a_1589_49.t1 CI.t2 VGND.t0 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X27 a_67_199.t2 a_488_21.t5 a_434_49.t1 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X28 VPWR.t5 B.t7 a_488_21.t0 VPB.t10 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X29 VGND.t6 a_1589_49.t5 a_1634_315.t2 VNB.t14 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X30 a_1261_49.t3 a_726_47.t7 COUT_N.t3 VPB.t9 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X31 VGND.t1 CI.t3 a_1261_49.t1 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
R0 B.n4 B.t6 246.258
R1 B.n1 B.t0 212.079
R2 B.n3 B.t7 212.079
R3 B.n0 B.t3 186.373
R4 B.n6 B.n0 154.962
R5 B.n2 B.t1 139.779
R6 B.n0 B.t2 138.172
R7 B.n1 B.t5 138.172
R8 B.n4 B.t4 138.172
R9 B.n5 B.n3 114.657
R10 B B.n5 98.905
R11 B.n2 B.n1 71.569
R12 B.n5 B.n4 18.987
R13 B.n6 B 4.65
R14 B B.n6 4.029
R15 B.n3 B.n2 2.921
R16 VPWR.n46 VPWR.n45 314.335
R17 VPWR.n25 VPWR.n24 308.015
R18 VPWR.n1 VPWR.n0 306.255
R19 VPWR.n3 VPWR.n2 175.816
R20 VPWR.n24 VPWR.t5 44.325
R21 VPWR.n45 VPWR.t2 42.355
R22 VPWR.n2 VPWR.t3 26.595
R23 VPWR.n2 VPWR.t1 26.595
R24 VPWR.n0 VPWR.t0 26.595
R25 VPWR.n0 VPWR.t7 26.595
R26 VPWR.n24 VPWR.t4 26.595
R27 VPWR.n45 VPWR.t6 26.595
R28 VPWR.n48 VPWR.n47 4.65
R29 VPWR.n5 VPWR.n4 4.65
R30 VPWR.n7 VPWR.n6 4.65
R31 VPWR.n9 VPWR.n8 4.65
R32 VPWR.n11 VPWR.n10 4.65
R33 VPWR.n13 VPWR.n12 4.65
R34 VPWR.n15 VPWR.n14 4.65
R35 VPWR.n17 VPWR.n16 4.65
R36 VPWR.n19 VPWR.n18 4.65
R37 VPWR.n21 VPWR.n20 4.65
R38 VPWR.n23 VPWR.n22 4.65
R39 VPWR.n26 VPWR.n25 4.65
R40 VPWR.n28 VPWR.n27 4.65
R41 VPWR.n30 VPWR.n29 4.65
R42 VPWR.n32 VPWR.n31 4.65
R43 VPWR.n34 VPWR.n33 4.65
R44 VPWR.n36 VPWR.n35 4.65
R45 VPWR.n38 VPWR.n37 4.65
R46 VPWR.n40 VPWR.n39 4.65
R47 VPWR.n42 VPWR.n41 4.65
R48 VPWR.n44 VPWR.n43 4.65
R49 VPWR.n3 VPWR.n1 4.018
R50 VPWR.n47 VPWR.n46 0.376
R51 VPWR.n5 VPWR.n3 0.145
R52 VPWR.n7 VPWR.n5 0.119
R53 VPWR.n9 VPWR.n7 0.119
R54 VPWR.n11 VPWR.n9 0.119
R55 VPWR.n13 VPWR.n11 0.119
R56 VPWR.n15 VPWR.n13 0.119
R57 VPWR.n17 VPWR.n15 0.119
R58 VPWR.n19 VPWR.n17 0.119
R59 VPWR.n21 VPWR.n19 0.119
R60 VPWR.n23 VPWR.n21 0.119
R61 VPWR.n26 VPWR.n23 0.119
R62 VPWR.n28 VPWR.n26 0.119
R63 VPWR.n30 VPWR.n28 0.119
R64 VPWR.n32 VPWR.n30 0.119
R65 VPWR.n34 VPWR.n32 0.119
R66 VPWR.n36 VPWR.n34 0.119
R67 VPWR.n38 VPWR.n36 0.119
R68 VPWR.n40 VPWR.n38 0.119
R69 VPWR.n42 VPWR.n40 0.119
R70 VPWR.n44 VPWR.n42 0.119
R71 VPWR.n48 VPWR.n44 0.119
R72 VPWR.n49 VPWR.n48 0.119
R73 VPWR VPWR.n49 0.022
R74 a_1144_49.n0 a_1144_49.t1 305.863
R75 a_1144_49.n3 a_1144_49.n2 302.963
R76 a_1144_49.n1 a_1144_49.n0 292.5
R77 a_1144_49.n2 a_1144_49.t3 184.271
R78 a_1144_49.n4 a_1144_49.n1 79.738
R79 a_1144_49.n1 a_1144_49.t0 31.66
R80 a_1144_49.n4 a_1144_49.n3 24.827
R81 a_1144_49.n5 a_1144_49.n4 24.818
R82 a_1144_49.n3 a_1144_49.t2 18.62
R83 VPB.t9 VPB.t8 899.688
R84 VPB.t5 VPB.t15 668.847
R85 VPB.t2 VPB.t12 662.928
R86 VPB.t4 VPB.t3 642.211
R87 VPB.t11 VPB.t10 621.495
R88 VPB.t0 VPB.t1 571.183
R89 VPB.t13 VPB.t6 556.386
R90 VPB.t10 VPB.t13 301.869
R91 VPB.t14 VPB.t2 295.95
R92 VPB.t3 VPB.t11 287.071
R93 VPB.t1 VPB.t7 248.598
R94 VPB.t15 VPB.t0 248.598
R95 VPB.t8 VPB.t5 248.598
R96 VPB.t6 VPB.t9 248.598
R97 VPB.t12 VPB.t4 248.598
R98 VPB VPB.t14 195.327
R99 a_67_199.n0 a_67_199.t2 426.936
R100 a_67_199.t0 a_67_199.n7 413.061
R101 a_67_199.n1 a_67_199.t6 236.179
R102 a_67_199.n4 a_67_199.t1 209.333
R103 a_67_199.n1 a_67_199.t7 165.486
R104 a_67_199.n8 a_67_199.t0 141.84
R105 a_67_199.n4 a_67_199.n3 92.5
R106 a_67_199.n6 a_67_199.n1 76
R107 a_67_199.n7 a_67_199.n6 69.572
R108 a_67_199.n0 a_67_199.t5 52.071
R109 a_67_199.n5 a_67_199.n2 48.937
R110 a_67_199.n6 a_67_199.n5 45.347
R111 a_67_199.n5 a_67_199.n4 41.064
R112 a_67_199.n3 a_67_199.t4 25.312
R113 a_67_199.n7 a_67_199.n0 15.058
R114 a_67_199.n2 a_67_199.t3 14.183
R115 a_28_47.n2 a_28_47.t3 452.585
R116 a_28_47.n1 a_28_47.t1 244.5
R117 a_28_47.n0 a_28_47.t2 223.111
R118 a_28_47.n3 a_28_47.t5 170.375
R119 a_28_47.n0 a_28_47.t0 168.089
R120 a_28_47.n2 a_28_47.n1 138.205
R121 a_28_47.t4 a_28_47.n3 123.83
R122 a_28_47.n3 a_28_47.n2 121.747
R123 a_28_47.n1 a_28_47.n0 74.913
R124 a_488_21.t0 a_488_21.n3 301.63
R125 a_488_21.n0 a_488_21.t3 192.945
R126 a_488_21.n1 a_488_21.t5 186.373
R127 a_488_21.n3 a_488_21.t1 155.381
R128 a_488_21.n0 a_488_21.t4 141.386
R129 a_488_21.n1 a_488_21.t2 138.172
R130 a_488_21.n2 a_488_21.n0 108.815
R131 a_488_21.n3 a_488_21.n2 94.366
R132 a_488_21.n2 a_488_21.n1 43.087
R133 VGND.n2 VGND.n1 116.217
R134 VGND.n46 VGND.n45 114.711
R135 VGND.n3 VGND.n0 113.492
R136 VGND.n25 VGND.n24 64.067
R137 VGND.n24 VGND.t4 38.437
R138 VGND.n0 VGND.t3 32.479
R139 VGND.n1 VGND.t6 30.937
R140 VGND.n45 VGND.t7 30.937
R141 VGND.n1 VGND.t0 26.854
R142 VGND.n45 VGND.t2 26.854
R143 VGND.n0 VGND.t1 25.312
R144 VGND.n24 VGND.t5 22.167
R145 VGND.n3 VGND.n2 9.026
R146 VGND.n47 VGND.n46 6.029
R147 VGND.n5 VGND.n4 4.65
R148 VGND.n7 VGND.n6 4.65
R149 VGND.n9 VGND.n8 4.65
R150 VGND.n11 VGND.n10 4.65
R151 VGND.n13 VGND.n12 4.65
R152 VGND.n15 VGND.n14 4.65
R153 VGND.n17 VGND.n16 4.65
R154 VGND.n19 VGND.n18 4.65
R155 VGND.n21 VGND.n20 4.65
R156 VGND.n23 VGND.n22 4.65
R157 VGND.n26 VGND.n25 4.65
R158 VGND.n28 VGND.n27 4.65
R159 VGND.n30 VGND.n29 4.65
R160 VGND.n32 VGND.n31 4.65
R161 VGND.n34 VGND.n33 4.65
R162 VGND.n36 VGND.n35 4.65
R163 VGND.n38 VGND.n37 4.65
R164 VGND.n40 VGND.n39 4.65
R165 VGND.n42 VGND.n41 4.65
R166 VGND.n44 VGND.n43 4.65
R167 VGND.n5 VGND.n3 0.141
R168 VGND.n47 VGND.n44 0.132
R169 VGND VGND.n47 0.129
R170 VGND.n7 VGND.n5 0.119
R171 VGND.n9 VGND.n7 0.119
R172 VGND.n11 VGND.n9 0.119
R173 VGND.n13 VGND.n11 0.119
R174 VGND.n15 VGND.n13 0.119
R175 VGND.n17 VGND.n15 0.119
R176 VGND.n19 VGND.n17 0.119
R177 VGND.n21 VGND.n19 0.119
R178 VGND.n23 VGND.n21 0.119
R179 VGND.n26 VGND.n23 0.119
R180 VGND.n28 VGND.n26 0.119
R181 VGND.n30 VGND.n28 0.119
R182 VGND.n32 VGND.n30 0.119
R183 VGND.n34 VGND.n32 0.119
R184 VGND.n36 VGND.n34 0.119
R185 VGND.n38 VGND.n36 0.119
R186 VGND.n40 VGND.n38 0.119
R187 VGND.n42 VGND.n40 0.119
R188 VGND.n44 VGND.n42 0.119
R189 VNB.t8 VNB.t9 6893.33
R190 VNB VNB.t15 6115.42
R191 VNB.t6 VNB.t12 5556.41
R192 VNB.t5 VNB.t14 5524.44
R193 VNB.t3 VNB.t2 5058.39
R194 VNB.t10 VNB.t4 4864.44
R195 VNB.t0 VNB.t1 4545.05
R196 VNB.t11 VNB.t13 4520.88
R197 VNB.t2 VNB.t11 3215.38
R198 VNB.t1 VNB.t7 2296.7
R199 VNB.t13 VNB.t10 2285.08
R200 VNB.t14 VNB.t0 2248.62
R201 VNB.t15 VNB.t6 2248.62
R202 VNB.t9 VNB.t5 2151.11
R203 VNB.t4 VNB.t8 2077.78
R204 VNB.t12 VNB.t3 2053.33
R205 a_434_49.n5 a_434_49.n4 303.399
R206 a_434_49.n1 a_434_49.t5 240.144
R207 a_434_49.n0 a_434_49.t6 186.373
R208 a_434_49.n1 a_434_49.t7 165.266
R209 a_434_49.n0 a_434_49.t4 146.205
R210 a_434_49.n4 a_434_49.n3 104.412
R211 a_434_49.n2 a_434_49.n0 50.036
R212 a_434_49.t1 a_434_49.n5 31.66
R213 a_434_49.n5 a_434_49.t2 31.66
R214 a_434_49.n3 a_434_49.t0 25.312
R215 a_434_49.n3 a_434_49.t3 25.312
R216 a_434_49.n2 a_434_49.n1 12.573
R217 a_434_49.n4 a_434_49.n2 8.272
R218 a_1261_49.n0 a_1261_49.t3 295.197
R219 a_1261_49.n0 a_1261_49.t0 233.316
R220 a_1261_49.t2 a_1261_49.n1 169.084
R221 a_1261_49.n1 a_1261_49.t1 136.304
R222 a_1261_49.n1 a_1261_49.n0 12.5
R223 COUT_N COUT_N.n1 300.796
R224 COUT_N.n2 COUT_N.n0 100.405
R225 COUT_N.n1 COUT_N.t3 31.66
R226 COUT_N.n1 COUT_N.t0 31.66
R227 COUT_N.n0 COUT_N.t2 26.25
R228 COUT_N.n0 COUT_N.t1 25.312
R229 COUT_N.n2 COUT_N 24.651
R230 COUT_N.n2  10.164
R231  COUT_N.n2 7.585
R232 a_1710_49.n1 a_1710_49.t5 241.534
R233 a_1710_49.n3 a_1710_49.n2 174.607
R234 a_1710_49.n1 a_1710_49.t4 169.234
R235 a_1710_49.n2 a_1710_49.n0 160.878
R236 a_1710_49.n2 a_1710_49.n1 111.648
R237 a_1710_49.t1 a_1710_49.n3 31.66
R238 a_1710_49.n3 a_1710_49.t2 31.66
R239 a_1710_49.n0 a_1710_49.t3 29.062
R240 a_1710_49.n0 a_1710_49.t0 25.312
R241 a_1589_49.n2 a_1589_49.t3 280.307
R242 a_1589_49.n0 a_1589_49.t4 241.534
R243 a_1589_49.n2 a_1589_49.t0 196.673
R244 a_1589_49.n0 a_1589_49.t5 167.627
R245 a_1589_49.t2 a_1589_49.n3 126.594
R246 a_1589_49.n1 a_1589_49.t1 123.471
R247 a_1589_49.n1 a_1589_49.n0 76
R248 a_1589_49.n3 a_1589_49.n1 21.997
R249 a_1589_49.n3 a_1589_49.n2 14.552
R250 SUM.n1 SUM.t0 173.927
R251 SUM.n0 SUM.t1 80.894
R252 SUM  21.76
R253 SUM.n2 SUM 17.92
R254  SUM.n1 10.069
R255  SUM.n0 6.846
R256 SUM.n0  5.573
R257  SUM.n2 3.84
R258 SUM.n1  3.252
R259 SUM.n2  2.258
R260 a_726_47.n4 a_726_47.n2 531.192
R261 a_726_47.n5 a_726_47.n4 292.5
R262 a_726_47.n1 a_726_47.t7 195.136
R263 a_726_47.n4 a_726_47.n3 166.553
R264 a_726_47.n0 a_726_47.t4 164.841
R265 a_726_47.n0 a_726_47.t6 138.172
R266 a_726_47.n1 a_726_47.t5 138.172
R267 a_726_47.n2 a_726_47.n1 130.724
R268 a_726_47.n3 a_726_47.t1 62.592
R269 a_726_47.n2 a_726_47.n0 51.431
R270 a_726_47.n5 a_726_47.t3 50.66
R271 a_726_47.t0 a_726_47.n5 32.248
R272 a_726_47.n3 a_726_47.t2 20.109
R273 a_1634_315.n1 a_1634_315.t3 310.76
R274 a_1634_315.t1 a_1634_315.n1 173.635
R275 a_1634_315.n0 a_1634_315.t0 156.562
R276 a_1634_315.n1 a_1634_315.n0 128.172
R277 a_1634_315.n0 a_1634_315.t2 27.187
R278 CI.n1 CI.t0 215.73
R279 CI.n0 CI.t1 212.079
R280 CI.n1 CI.t2 139.779
R281 CI.n0 CI.t3 138.172
R282 CI.n2 CI.n0 100.051
R283 CI CI.n2 77.582
R284 CI.n2 CI.n1 37.245
R285 A.n0 A.t0 230.361
R286 A.n0 A.t1 158.061
R287 A A.n0 83.04
C0 VPB VPWR 0.25fF
C1 SUM VGND 0.11fF
C2 B VGND 0.27fF
C3 VPWR SUM 0.17fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__fill_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__fill_1 VPWR VGND VPB VNB
.ends

* NGSPICE file created from sky130_fd_sc_hd__fill_2.ext - technology: sky130A

.subckt sky130_fd_sc_hd__fill_2 VGND VPWR VPB VNB
.ends

* NGSPICE file created from sky130_fd_sc_hd__fill_4.ext - technology: sky130A

.subckt sky130_fd_sc_hd__fill_4 VGND VPWR VPB VNB
.ends

* NGSPICE file created from sky130_fd_sc_hd__fill_8.ext - technology: sky130A

.subckt sky130_fd_sc_hd__fill_8 VGND VPWR VPB VNB
C0 VPWR VGND 0.12fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__ha_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__ha_1 VGND VPWR B A COUT SUM VNB VPB
X0 a_297_47.t2 a_250_199.t3 a_79_21.t2 VNB.t6 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1 a_297_47.t0 A.t0 VGND.t0 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 COUT.t0 a_250_199.t4 VPWR.t5 VPB.t6 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 a_250_199.t1 B.t0 VPWR.t3 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 a_376_413.t0 B.t1 a_79_21.t0 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 a_79_21.t1 a_250_199.t5 VPWR.t4 VPB.t5 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 a_674_47.t0 B.t2 a_250_199.t2 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7 VPWR.t0 A.t1 a_376_413.t1 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 VGND.t3 B.t3 a_297_47.t1 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9 COUT.t1 a_250_199.t6 VGND.t4 VNB.t5 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 VPWR.t2 a_79_21.t3 SUM.t0 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 VPWR.t1 A.t2 a_250_199.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12 VGND.t1 A.t3 a_674_47.t1 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13 VGND.t2 a_79_21.t4 SUM.t1 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
R0 a_250_199.n4 a_250_199.n3 387.844
R1 a_250_199.n1 a_250_199.t5 334.721
R2 a_250_199.n0 a_250_199.t4 241.534
R3 a_250_199.n2 a_250_199.n1 211.905
R4 a_250_199.n1 a_250_199.t3 206.188
R5 a_250_199.n0 a_250_199.t6 169.234
R6 a_250_199.n2 a_250_199.t2 146.506
R7 a_250_199.n3 a_250_199.n2 77.65
R8 a_250_199.n3 a_250_199.n0 76
R9 a_250_199.t0 a_250_199.n4 68.011
R10 a_250_199.n4 a_250_199.t1 68.011
R11 a_79_21.n2 a_79_21.n1 392.263
R12 a_79_21.n0 a_79_21.t3 232.213
R13 a_79_21.n1 a_79_21.t2 167.686
R14 a_79_21.n0 a_79_21.t4 159.913
R15 a_79_21.n1 a_79_21.n0 105.364
R16 a_79_21.t0 a_79_21.n2 63.321
R17 a_79_21.n2 a_79_21.t1 63.321
R18 a_297_47.t0 a_297_47.n0 305.64
R19 a_297_47.n0 a_297_47.t1 38.571
R20 a_297_47.n0 a_297_47.t2 38.571
R21 VNB.t1 VNB.t3 6761.76
R22 VNB VNB.t0 6053.91
R23 VNB.t0 VNB.t6 5321.88
R24 VNB.t4 VNB.t1 2717.65
R25 VNB.t6 VNB.t4 2717.65
R26 VNB.t3 VNB.t2 2329.41
R27 VNB.t2 VNB.t5 2255.35
R28 A.n0 A.t0 405.292
R29 A.n1 A.t2 274.51
R30 A.n0 A.t1 250.548
R31 A.n1 A.t3 248.803
R32 A.n3 A.n0 140.752
R33 A.n2 A.n1 76
R34 A.n2 A 12.231
R35 A.n3 A.n2 4.551
R36 A A.n3 2.56
R37 VGND.n3 VGND.n0 115.917
R38 VGND.n8 VGND.t2 115.886
R39 VGND.n2 VGND.n1 107.239
R40 VGND.n0 VGND.t1 54.285
R41 VGND.n1 VGND.t0 38.571
R42 VGND.n1 VGND.t3 38.571
R43 VGND.n0 VGND.t4 25.934
R44 VGND.n5 VGND.n4 4.65
R45 VGND.n7 VGND.n6 4.65
R46 VGND.n9 VGND.n8 4.05
R47 VGND.n3 VGND.n2 3.983
R48 VGND.n5 VGND.n3 0.139
R49 VGND.n9 VGND.n7 0.134
R50 VGND VGND.n9 0.124
R51 VGND.n7 VGND.n5 0.119
R52 VPWR.n3 VPWR.n2 318.164
R53 VPWR.n5 VPWR.n4 292.5
R54 VPWR.n1 VPWR.n0 292.5
R55 VPWR.n13 VPWR.n12 292.5
R56 VPWR.n19 VPWR.n17 170.062
R57 VPWR.n12 VPWR.t4 100.845
R58 VPWR.n2 VPWR.t1 89.119
R59 VPWR.n0 VPWR.t3 86.773
R60 VPWR.n4 VPWR.t0 86.773
R61 VPWR.n2 VPWR.t5 29.315
R62 VPWR.n17 VPWR.t2 25.61
R63 VPWR.n3 VPWR.n1 4.814
R64 VPWR.n15 VPWR.n14 4.65
R65 VPWR.n7 VPWR.n6 4.65
R66 VPWR.n9 VPWR.n8 4.65
R67 VPWR.n11 VPWR.n10 4.65
R68 VPWR.n20 VPWR.n19 4.65
R69 VPWR.n17 VPWR.n16 2.345
R70 VPWR.n6 VPWR.n5 2.052
R71 VPWR.n14 VPWR.n13 1.328
R72 VPWR.n19 VPWR.n18 0.241
R73 VPWR.n7 VPWR.n3 0.212
R74 VPWR.n9 VPWR.n7 0.119
R75 VPWR.n11 VPWR.n9 0.119
R76 VPWR.n15 VPWR.n11 0.119
R77 VPWR.n20 VPWR.n15 0.119
R78 VPWR.n21 VPWR.n20 0.119
R79 VPWR VPWR.n21 0.02
R80 COUT.n2 COUT.n1 292.5
R81 COUT.n3 COUT.n2 146.895
R82 COUT.n0 COUT.t1 82.802
R83 COUT.n1 COUT.n0 63.47
R84 COUT.n2 COUT.t0 26.595
R85 COUT.n3 COUT 10.204
R86 COUT.n0 COUT 5.593
R87 COUT.n1 COUT 5.082
R88 COUT COUT.n3 2.553
R89 VPB.t2 VPB.t5 541.588
R90 VPB.t1 VPB.t3 509.034
R91 VPB.t4 VPB.t1 325.545
R92 VPB.t0 VPB.t6 281.152
R93 VPB.t3 VPB.t0 260.436
R94 VPB.t5 VPB.t4 248.598
R95 VPB VPB.t2 189.408
R96 B.n0 B.t2 419.874
R97 B.n2 B.t3 360.791
R98 B.n2 B.t1 167.991
R99 B.n0 B.t0 154.226
R100 B.n1 B.n0 139.623
R101 B.n3 B.n2 76
R102 B B.n3 9.022
R103 B.n3 B.n1 3.357
R104 B.n1 B 1.888
R105 a_376_413.t0 a_376_413.t1 187.619
R106 a_674_47.t0 a_674_47.t1 60
R107 SUM.n4 SUM.n3 292.5
R108 SUM.n5 SUM.n4 146.904
R109 SUM.n0 SUM.t1 82.765
R110 SUM.n4 SUM.t0 26.595
R111 SUM SUM.n1 15.582
R112 SUM.n5 SUM 10.356
R113 SUM SUM.n0 6.909
R114 SUM.n2 SUM 6.678
R115 SUM.n0 SUM 5.674
R116 SUM.n3 SUM 5.158
R117 SUM.n2 SUM 4.585
R118 SUM.n1 SUM 3.339
R119 SUM.n3 SUM.n2 3.247
R120 SUM SUM.n5 2.591
R121 SUM.n1 SUM 2.292
C0 VPWR VGND 0.10fF
C1 SUM VGND 0.12fF
C2 SUM VPWR 0.18fF
C3 VPWR B 0.11fF
C4 A B 0.41fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__ha_2.ext - technology: sky130A

.subckt sky130_fd_sc_hd__ha_2 VGND VPWR A COUT SUM B VNB VPB
X0 VPWR.t3 A.t0 a_342_199.t0 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1 a_766_47.t0 B.t0 a_342_199.t1 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 VGND.t0 B.t1 a_389_47.t0 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3 COUT.t3 a_342_199.t3 VGND.t6 VNB.t8 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 VGND.t3 A.t1 a_766_47.t1 VNB.t5 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 a_342_199.t2 B.t2 VPWR.t7 VPB.t8 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X6 a_468_369.t0 B.t3 a_79_21.t0 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X7 a_79_21.t2 a_342_199.t4 VPWR.t4 VPB.t7 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X8 a_389_47.t2 a_342_199.t5 a_79_21.t1 VNB.t7 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9 a_389_47.t1 A.t2 VGND.t4 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10 COUT.t1 a_342_199.t6 VPWR.t6 VPB.t6 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 VPWR.t5 a_342_199.t7 COUT.t0 VPB.t5 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 VGND.t1 a_79_21.t3 SUM.t3 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 VPWR.t0 a_79_21.t4 SUM.t1 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14 VGND.t5 a_342_199.t8 COUT.t2 VNB.t6 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X15 SUM.t0 a_79_21.t5 VPWR.t1 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16 VPWR.t2 A.t3 a_468_369.t1 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X17 SUM.t2 a_79_21.t6 VGND.t2 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
R0 A.n1 A.t3 299.068
R1 A.n0 A.t0 272.745
R2 A.n0 A.t1 224.545
R3 A.n1 A.t2 166.517
R4 A.n2 A.n1 141.129
R5 A.n3 A.n0 76
R6 A A.n3 12.231
R7 A.n3 A.n2 5.12
R8 A.n2 A 1.991
R9 a_342_199.n5 a_342_199.n4 304.923
R10 a_342_199.n3 a_342_199.t4 299.374
R11 a_342_199.n4 a_342_199.n3 282.681
R12 a_342_199.n2 a_342_199.t1 224.156
R13 a_342_199.n0 a_342_199.t7 212.079
R14 a_342_199.n1 a_342_199.t6 212.079
R15 a_342_199.n3 a_342_199.t5 206.188
R16 a_342_199.n0 a_342_199.t8 139.779
R17 a_342_199.n1 a_342_199.t3 139.779
R18 a_342_199.n2 a_342_199.n1 84.033
R19 a_342_199.n4 a_342_199.n2 82.92
R20 a_342_199.n1 a_342_199.n0 67.187
R21 a_342_199.t0 a_342_199.n5 44.632
R22 a_342_199.n5 a_342_199.t2 44.632
R23 VPWR.n1 VPWR.n0 309.178
R24 VPWR.n10 VPWR.n9 292.5
R25 VPWR.n6 VPWR.n5 292.5
R26 VPWR.n19 VPWR.t4 194.287
R27 VPWR.n2 VPWR.t5 157.949
R28 VPWR.n24 VPWR.t1 153.887
R29 VPWR.n20 VPWR.n19 141.423
R30 VPWR.n0 VPWR.t3 58.484
R31 VPWR.n5 VPWR.t7 56.945
R32 VPWR.n9 VPWR.t2 56.945
R33 VPWR.n0 VPWR.t6 31.605
R34 VPWR.n19 VPWR.t0 30.225
R35 VPWR.n4 VPWR.n3 4.65
R36 VPWR.n8 VPWR.n7 4.65
R37 VPWR.n12 VPWR.n11 4.65
R38 VPWR.n14 VPWR.n13 4.65
R39 VPWR.n16 VPWR.n15 4.65
R40 VPWR.n18 VPWR.n17 4.65
R41 VPWR.n21 VPWR.n20 4.65
R42 VPWR.n23 VPWR.n22 4.65
R43 VPWR.n25 VPWR.n24 4.65
R44 VPWR.n2 VPWR.n1 3.814
R45 VPWR.n11 VPWR.n10 1.813
R46 VPWR.n7 VPWR.n6 0.746
R47 VPWR.n4 VPWR.n2 0.241
R48 VPWR.n8 VPWR.n4 0.119
R49 VPWR.n12 VPWR.n8 0.119
R50 VPWR.n14 VPWR.n12 0.119
R51 VPWR.n16 VPWR.n14 0.119
R52 VPWR.n18 VPWR.n16 0.119
R53 VPWR.n21 VPWR.n18 0.119
R54 VPWR.n23 VPWR.n21 0.119
R55 VPWR.n25 VPWR.n23 0.119
R56 VPWR VPWR.n25 0.02
R57 VPB.t0 VPB.t7 541.588
R58 VPB.t3 VPB.t8 509.034
R59 VPB.t2 VPB.t3 325.545
R60 VPB.t4 VPB.t6 281.152
R61 VPB.t6 VPB.t5 272.274
R62 VPB.t1 VPB.t0 272.274
R63 VPB.t8 VPB.t4 260.436
R64 VPB.t7 VPB.t2 248.598
R65 VPB VPB.t1 189.408
R66 B.n0 B.t0 382.385
R67 B.n1 B.t3 261.177
R68 B.n1 B.t1 232.257
R69 B.n0 B.t2 218.505
R70 B B.n0 117.034
R71 B.n2 B.n1 76
R72 B.n2 B 7.763
R73 B B.n2 6.504
R74 a_766_47.t0 a_766_47.t1 60
R75 VNB.t4 VNB.t1 6761.76
R76 VNB VNB.t3 6053.91
R77 VNB.t2 VNB.t7 5321.88
R78 VNB.t0 VNB.t4 2717.65
R79 VNB.t7 VNB.t0 2717.65
R80 VNB.t1 VNB.t5 2329.41
R81 VNB.t5 VNB.t8 2255.35
R82 VNB.t8 VNB.t6 2224.18
R83 VNB.t3 VNB.t2 2224.18
R84 a_389_47.n0 a_389_47.t1 305.64
R85 a_389_47.t0 a_389_47.n0 38.571
R86 a_389_47.n0 a_389_47.t2 38.571
R87 VGND.n16 VGND.t1 115.887
R88 VGND.n2 VGND.t5 114.311
R89 VGND.n1 VGND.n0 111.956
R90 VGND.n20 VGND.t2 110.226
R91 VGND.n10 VGND.n9 107.239
R92 VGND.n0 VGND.t3 54.285
R93 VGND.n9 VGND.t4 38.571
R94 VGND.n9 VGND.t0 38.571
R95 VGND.n0 VGND.t6 25.934
R96 VGND.n21 VGND.n20 4.65
R97 VGND.n4 VGND.n3 4.65
R98 VGND.n6 VGND.n5 4.65
R99 VGND.n8 VGND.n7 4.65
R100 VGND.n11 VGND.n10 4.65
R101 VGND.n13 VGND.n12 4.65
R102 VGND.n15 VGND.n14 4.65
R103 VGND.n17 VGND.n16 4.65
R104 VGND.n19 VGND.n18 4.65
R105 VGND.n2 VGND.n1 3.953
R106 VGND.n4 VGND.n2 0.221
R107 VGND.n6 VGND.n4 0.119
R108 VGND.n8 VGND.n6 0.119
R109 VGND.n11 VGND.n8 0.119
R110 VGND.n13 VGND.n11 0.119
R111 VGND.n15 VGND.n13 0.119
R112 VGND.n17 VGND.n15 0.119
R113 VGND.n19 VGND.n17 0.119
R114 VGND.n21 VGND.n19 0.119
R115 VGND VGND.n21 0.02
R116 COUT.n0 COUT 298.9
R117 COUT.n3 COUT.n0 292.5
R118 COUT COUT.n1 93.469
R119 COUT.n2 COUT.n1 92.5
R120 COUT.n3 COUT.n2 64.406
R121 COUT.n0 COUT.t0 34.475
R122 COUT.n1 COUT.t2 32.307
R123 COUT.n0 COUT.t1 26.595
R124 COUT.n1 COUT.t3 24.923
R125 COUT.n2 COUT 12.218
R126 COUT COUT.n3 3.84
R127 a_79_21.n3 a_79_21.n2 406.193
R128 a_79_21.n1 a_79_21.t4 212.079
R129 a_79_21.n0 a_79_21.t5 212.079
R130 a_79_21.n2 a_79_21.t1 167.686
R131 a_79_21.n1 a_79_21.t3 139.779
R132 a_79_21.n0 a_79_21.t6 139.779
R133 a_79_21.n2 a_79_21.n1 132.385
R134 a_79_21.n1 a_79_21.n0 67.187
R135 a_79_21.t0 a_79_21.n3 41.554
R136 a_79_21.n3 a_79_21.t2 41.554
R137 a_468_369.t0 a_468_369.t1 123.125
R138 SUM.n5 SUM.n4 292.5
R139 SUM.n6 SUM.n5 146.914
R140 SUM.n1 SUM.n0 43.625
R141 SUM.n5 SUM.t0 34.475
R142 SUM.n0 SUM.t2 32.307
R143 SUM.n5 SUM.t1 26.595
R144 SUM.n0 SUM.t3 24.923
R145 SUM SUM.n2 15.928
R146 SUM.n6 SUM 10.512
R147 SUM.n3 SUM 6.826
R148 SUM SUM.n1 6.672
R149 SUM.n1 SUM 5.763
R150 SUM.n4 SUM 5.236
R151 SUM.n3 SUM 4.654
R152 SUM.n2 SUM 3.413
R153 SUM.n4 SUM.n3 3.296
R154 SUM SUM.n6 2.63
R155 SUM.n2 SUM 2.327
C0 SUM VGND 0.20fF
C1 VPWR VGND 0.16fF
C2 VPWR COUT 0.18fF
C3 VPWR SUM 0.26fF
C4 B A 0.40fF
C5 VPB VPWR 0.12fF
C6 COUT VGND 0.14fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__ha_4.ext - technology: sky130A

.subckt sky130_fd_sc_hd__ha_4 VGND VPWR A COUT SUM B VNB VPB
X0 a_467_47.t3 B.t0 VGND.t5 VNB.t9 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 a_1325_47.t0 B.t1 a_514_199.t1 VNB.t8 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 COUT.t3 a_514_199.t6 VGND.t0 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 COUT.t2 a_514_199.t7 VGND.t1 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 a_467_47.t0 a_514_199.t8 a_79_21.t1 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 a_1167_47.t1 A.t0 VGND.t10 VNB.t14 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 a_717_297.t1 A.t1 VPWR.t15 VPB.t17 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 VPWR.t7 B.t2 a_514_199.t3 VPB.t9 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 VPWR.t5 a_514_199.t9 COUT.t7 VPB.t5 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 VPWR.t11 a_79_21.t6 SUM.t7 VPB.t13 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 VGND.t11 A.t2 a_1325_47.t1 VNB.t15 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 a_514_199.t4 A.t3 VPWR.t14 VPB.t16 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 COUT.t6 a_514_199.t10 VPWR.t4 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13 a_79_21.t0 a_514_199.t11 a_467_47.t1 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14 VPWR.t3 a_514_199.t12 COUT.t5 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 SUM.t6 a_79_21.t7 VPWR.t10 VPB.t12 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16 VPWR.t1 a_514_199.t13 a_79_21.t3 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17 VGND.t12 A.t4 a_467_47.t4 VNB.t16 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X18 VPWR.t9 a_79_21.t8 SUM.t5 VPB.t11 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X19 COUT.t4 a_514_199.t14 VPWR.t2 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X20 VGND.t6 a_79_21.t9 SUM.t3 VNB.t10 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X21 VGND.t7 a_79_21.t10 SUM.t2 VNB.t11 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X22 SUM.t1 a_79_21.t11 VGND.t8 VNB.t12 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X23 a_79_21.t2 a_514_199.t15 VPWR.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X24 a_514_199.t0 B.t3 a_1167_47.t0 VNB.t7 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X25 VPWR.t12 A.t5 a_890_297.t1 VPB.t15 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X26 VPWR.t13 A.t6 a_514_199.t5 VPB.t14 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X27 VGND.t4 B.t4 a_467_47.t2 VNB.t6 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X28 VGND.t2 a_514_199.t16 COUT.t1 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X29 VGND.t3 a_514_199.t17 COUT.t0 VNB.t5 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X30 a_890_297.t0 B.t5 a_79_21.t4 VPB.t8 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X31 a_514_199.t2 B.t6 VPWR.t6 VPB.t7 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X32 VGND.t13 A.t7 a_467_47.t5 VNB.t17 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X33 SUM.t4 a_79_21.t12 VPWR.t8 VPB.t10 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X34 a_79_21.t5 B.t7 a_717_297.t0 VPB.t6 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X35 SUM.t0 a_79_21.t13 VGND.t9 VNB.t13 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
R0 B B.n4 374.85
R1 B.n0 B.t6 212.079
R2 B.n1 B.t2 212.079
R3 B.n4 B.t5 212.079
R4 B.n3 B.t7 212.079
R5 B.n0 B.t1 139.779
R6 B.n1 B.t3 139.779
R7 B.n4 B.t4 139.779
R8 B.n3 B.t0 139.779
R9 B B.n2 79.06
R10 B.n4 B.n3 61.345
R11 B.n2 B.n0 46.739
R12 B.n2 B.n1 14.606
R13 VGND.n20 VGND.t4 190.315
R14 VGND.n2 VGND.t3 117.848
R15 VGND.n1 VGND.n0 116.88
R16 VGND.n42 VGND.t9 113.732
R17 VGND.n32 VGND.t7 110.227
R18 VGND.n6 VGND.n5 107.239
R19 VGND.n13 VGND.n12 107.239
R20 VGND.n24 VGND.n23 106.201
R21 VGND.n37 VGND.n36 74.084
R22 VGND.n5 VGND.t0 32.307
R23 VGND.n5 VGND.t11 32.307
R24 VGND.n23 VGND.t5 27.692
R25 VGND.n23 VGND.t12 26.769
R26 VGND.n0 VGND.t1 24.923
R27 VGND.n0 VGND.t2 24.923
R28 VGND.n12 VGND.t10 24.923
R29 VGND.n12 VGND.t13 24.923
R30 VGND.n36 VGND.t8 24.923
R31 VGND.n36 VGND.t6 24.923
R32 VGND.n43 VGND.n42 4.65
R33 VGND.n4 VGND.n3 4.65
R34 VGND.n7 VGND.n6 4.65
R35 VGND.n9 VGND.n8 4.65
R36 VGND.n11 VGND.n10 4.65
R37 VGND.n15 VGND.n14 4.65
R38 VGND.n17 VGND.n16 4.65
R39 VGND.n19 VGND.n18 4.65
R40 VGND.n22 VGND.n21 4.65
R41 VGND.n25 VGND.n24 4.65
R42 VGND.n27 VGND.n26 4.65
R43 VGND.n29 VGND.n28 4.65
R44 VGND.n31 VGND.n30 4.65
R45 VGND.n33 VGND.n32 4.65
R46 VGND.n35 VGND.n34 4.65
R47 VGND.n39 VGND.n38 4.65
R48 VGND.n41 VGND.n40 4.65
R49 VGND.n2 VGND.n1 3.821
R50 VGND.n21 VGND.n20 3.764
R51 VGND.n38 VGND.n37 3.764
R52 VGND.n14 VGND.n13 2.635
R53 VGND.n4 VGND.n2 0.234
R54 VGND.n7 VGND.n4 0.119
R55 VGND.n9 VGND.n7 0.119
R56 VGND.n11 VGND.n9 0.119
R57 VGND.n15 VGND.n11 0.119
R58 VGND.n17 VGND.n15 0.119
R59 VGND.n19 VGND.n17 0.119
R60 VGND.n22 VGND.n19 0.119
R61 VGND.n25 VGND.n22 0.119
R62 VGND.n27 VGND.n25 0.119
R63 VGND.n29 VGND.n27 0.119
R64 VGND.n31 VGND.n29 0.119
R65 VGND.n33 VGND.n31 0.119
R66 VGND.n35 VGND.n33 0.119
R67 VGND.n39 VGND.n35 0.119
R68 VGND.n41 VGND.n39 0.119
R69 VGND.n43 VGND.n41 0.119
R70 VGND VGND.n43 0.02
R71 a_467_47.n1 a_467_47.t1 236.843
R72 a_467_47.n2 a_467_47.t5 196.224
R73 a_467_47.n3 a_467_47.n2 102.664
R74 a_467_47.n1 a_467_47.n0 92.5
R75 a_467_47.n2 a_467_47.n1 75.293
R76 a_467_47.n0 a_467_47.t4 24.923
R77 a_467_47.n0 a_467_47.t0 24.923
R78 a_467_47.n3 a_467_47.t2 24.923
R79 a_467_47.t3 a_467_47.n3 24.923
R80 VNB VNB.t13 6053.91
R81 VNB.t6 VNB.t17 4665.93
R82 VNB.t11 VNB.t3 4545.05
R83 VNB.t15 VNB.t0 2417.58
R84 VNB.t16 VNB.t9 2151.65
R85 VNB.t1 VNB.t5 2030.77
R86 VNB.t4 VNB.t1 2030.77
R87 VNB.t0 VNB.t4 2030.77
R88 VNB.t8 VNB.t15 2030.77
R89 VNB.t7 VNB.t8 2030.77
R90 VNB.t17 VNB.t14 2030.77
R91 VNB.t9 VNB.t6 2030.77
R92 VNB.t2 VNB.t16 2030.77
R93 VNB.t3 VNB.t2 2030.77
R94 VNB.t12 VNB.t11 2030.77
R95 VNB.t10 VNB.t12 2030.77
R96 VNB.t13 VNB.t10 2030.77
R97 VNB.t14 VNB.t7 1789.01
R98 a_514_199.n13 a_514_199.n12 335.009
R99 a_514_199.n13 a_514_199.n9 304.923
R100 a_514_199.n15 a_514_199.n14 304.923
R101 a_514_199.n11 a_514_199.t15 215.73
R102 a_514_199.n10 a_514_199.t13 212.079
R103 a_514_199.n1 a_514_199.t9 212.079
R104 a_514_199.n2 a_514_199.t10 212.079
R105 a_514_199.n4 a_514_199.t12 212.079
R106 a_514_199.n5 a_514_199.t14 212.079
R107 a_514_199.n8 a_514_199.n0 198.662
R108 a_514_199.n10 a_514_199.t8 143.43
R109 a_514_199.n11 a_514_199.t11 139.779
R110 a_514_199.n1 a_514_199.t17 139.779
R111 a_514_199.n2 a_514_199.t7 139.779
R112 a_514_199.n4 a_514_199.t16 139.779
R113 a_514_199.n5 a_514_199.t6 139.779
R114 a_514_199.n7 a_514_199.n3 101.6
R115 a_514_199.n14 a_514_199.n8 87.34
R116 a_514_199.n7 a_514_199.n6 76
R117 a_514_199.n14 a_514_199.n13 63.247
R118 a_514_199.n2 a_514_199.n1 61.345
R119 a_514_199.n12 a_514_199.n11 48.93
R120 a_514_199.n3 a_514_199.n2 36.515
R121 a_514_199.n6 a_514_199.n5 36.515
R122 a_514_199.n8 a_514_199.n7 30.87
R123 a_514_199.n9 a_514_199.t3 26.595
R124 a_514_199.n9 a_514_199.t4 26.595
R125 a_514_199.n15 a_514_199.t5 26.595
R126 a_514_199.t2 a_514_199.n15 26.595
R127 a_514_199.n0 a_514_199.t1 24.923
R128 a_514_199.n0 a_514_199.t0 24.923
R129 a_514_199.n6 a_514_199.n4 24.83
R130 a_514_199.n12 a_514_199.n10 8.763
R131 a_1325_47.t0 a_1325_47.t1 49.846
R132 COUT.n1 COUT 298.214
R133 COUT.n2 COUT.n1 292.5
R134 COUT.n3 COUT.n0 219.754
R135 COUT.n7 COUT.n4 147.464
R136 COUT.n6 COUT.n5 92.5
R137 COUT.n1 COUT.t7 26.595
R138 COUT.n1 COUT.t6 26.595
R139 COUT.n0 COUT.t5 26.595
R140 COUT.n0 COUT.t4 26.595
R141 COUT.n5 COUT.t0 24.923
R142 COUT.n5 COUT.t2 24.923
R143 COUT.n4 COUT.t1 24.923
R144 COUT.n4 COUT.t3 24.923
R145 COUT COUT.n7 13.028
R146 COUT.n3 COUT.n2 9.6
R147 COUT COUT.n6 8.914
R148 COUT.n6 COUT 6.628
R149 COUT.n2 COUT 3.428
R150 COUT COUT.n3 2.514
R151 COUT.n7 COUT 2.514
R152 a_79_21.n2 a_79_21.n0 411.463
R153 a_79_21.n6 a_79_21.t6 212.079
R154 a_79_21.n5 a_79_21.t7 212.079
R155 a_79_21.n4 a_79_21.t8 212.079
R156 a_79_21.n3 a_79_21.t12 212.079
R157 a_79_21.n2 a_79_21.n1 150.897
R158 a_79_21.n6 a_79_21.t10 139.779
R159 a_79_21.n5 a_79_21.t11 139.779
R160 a_79_21.n4 a_79_21.t9 139.779
R161 a_79_21.n3 a_79_21.t13 139.779
R162 a_79_21.n8 a_79_21.n7 128.264
R163 a_79_21.n7 a_79_21.n6 111.947
R164 a_79_21.n6 a_79_21.n5 61.345
R165 a_79_21.n5 a_79_21.n4 61.345
R166 a_79_21.n4 a_79_21.n3 61.345
R167 a_79_21.n7 a_79_21.n2 53.457
R168 a_79_21.n1 a_79_21.t3 26.595
R169 a_79_21.n1 a_79_21.t2 26.595
R170 a_79_21.n0 a_79_21.t4 26.595
R171 a_79_21.n0 a_79_21.t5 26.595
R172 a_79_21.t1 a_79_21.n8 24.923
R173 a_79_21.n8 a_79_21.t0 24.923
R174 A.n0 A.t5 267.289
R175 A.n3 A.n2 261.222
R176 A.n4 A.t6 241.534
R177 A.n2 A.t1 241.534
R178 A.n1 A.t3 212.079
R179 A.n4 A.t2 169.234
R180 A.n2 A.t4 169.234
R181 A.n1 A.t0 147.082
R182 A.n0 A.t7 139.779
R183 A.n3 A.n1 101.976
R184 A.n5 A.n4 86.666
R185 A A.n3 73.574
R186 A.n1 A.n0 54.042
R187 A A.n5 6.678
R188 A.n5 A 4.46
R189 a_1167_47.t0 a_1167_47.t1 40.615
R190 VPWR.n25 VPWR.n24 319.982
R191 VPWR.n16 VPWR.n15 309.178
R192 VPWR.n11 VPWR.n10 309.178
R193 VPWR.n6 VPWR.n5 309.178
R194 VPWR.n1 VPWR.n0 167.515
R195 VPWR.n2 VPWR.t5 162.173
R196 VPWR.n43 VPWR.t8 158.057
R197 VPWR.n38 VPWR.n37 131.359
R198 VPWR.n32 VPWR.t0 90.62
R199 VPWR.n32 VPWR.t11 60.085
R200 VPWR.n15 VPWR.t14 45.31
R201 VPWR.n15 VPWR.t12 45.31
R202 VPWR.n5 VPWR.t2 34.475
R203 VPWR.n5 VPWR.t13 34.475
R204 VPWR.n24 VPWR.t15 31.52
R205 VPWR.n37 VPWR.t10 26.595
R206 VPWR.n37 VPWR.t9 26.595
R207 VPWR.n24 VPWR.t1 26.595
R208 VPWR.n10 VPWR.t6 26.595
R209 VPWR.n10 VPWR.t7 26.595
R210 VPWR.n0 VPWR.t4 26.595
R211 VPWR.n0 VPWR.t3 26.595
R212 VPWR.n33 VPWR.n32 18.07
R213 VPWR.n26 VPWR.n25 13.176
R214 VPWR.n4 VPWR.n3 4.65
R215 VPWR.n7 VPWR.n6 4.65
R216 VPWR.n9 VPWR.n8 4.65
R217 VPWR.n12 VPWR.n11 4.65
R218 VPWR.n14 VPWR.n13 4.65
R219 VPWR.n17 VPWR.n16 4.65
R220 VPWR.n19 VPWR.n18 4.65
R221 VPWR.n21 VPWR.n20 4.65
R222 VPWR.n23 VPWR.n22 4.65
R223 VPWR.n27 VPWR.n26 4.65
R224 VPWR.n29 VPWR.n28 4.65
R225 VPWR.n31 VPWR.n30 4.65
R226 VPWR.n34 VPWR.n33 4.65
R227 VPWR.n36 VPWR.n35 4.65
R228 VPWR.n40 VPWR.n39 4.65
R229 VPWR.n42 VPWR.n41 4.65
R230 VPWR.n44 VPWR.n43 4.65
R231 VPWR.n2 VPWR.n1 3.821
R232 VPWR.n39 VPWR.n38 3.764
R233 VPWR.n4 VPWR.n2 0.234
R234 VPWR.n7 VPWR.n4 0.119
R235 VPWR.n9 VPWR.n7 0.119
R236 VPWR.n12 VPWR.n9 0.119
R237 VPWR.n14 VPWR.n12 0.119
R238 VPWR.n17 VPWR.n14 0.119
R239 VPWR.n19 VPWR.n17 0.119
R240 VPWR.n21 VPWR.n19 0.119
R241 VPWR.n23 VPWR.n21 0.119
R242 VPWR.n27 VPWR.n23 0.119
R243 VPWR.n29 VPWR.n27 0.119
R244 VPWR.n31 VPWR.n29 0.119
R245 VPWR.n34 VPWR.n31 0.119
R246 VPWR.n36 VPWR.n34 0.119
R247 VPWR.n40 VPWR.n36 0.119
R248 VPWR.n42 VPWR.n40 0.119
R249 VPWR.n44 VPWR.n42 0.119
R250 VPWR VPWR.n44 0.02
R251 a_717_297.t0 a_717_297.t1 58.115
R252 VPB.t13 VPB.t0 541.588
R253 VPB.t8 VPB.t15 429.127
R254 VPB.t15 VPB.t16 361.059
R255 VPB.t14 VPB.t1 295.95
R256 VPB.t17 VPB.t6 263.395
R257 VPB.t2 VPB.t17 263.395
R258 VPB.t4 VPB.t5 248.598
R259 VPB.t3 VPB.t4 248.598
R260 VPB.t1 VPB.t3 248.598
R261 VPB.t7 VPB.t14 248.598
R262 VPB.t9 VPB.t7 248.598
R263 VPB.t16 VPB.t9 248.598
R264 VPB.t6 VPB.t8 248.598
R265 VPB.t0 VPB.t2 248.598
R266 VPB.t12 VPB.t13 248.598
R267 VPB.t11 VPB.t12 248.598
R268 VPB.t10 VPB.t11 248.598
R269 VPB VPB.t10 189.408
R270 SUM.n7 SUM.n6 292.5
R271 SUM.n8 SUM.n7 146.914
R272 SUM.n2 SUM.n0 122.925
R273 SUM SUM.n3 93.469
R274 SUM.n4 SUM.n3 92.5
R275 SUM.n2 SUM.n1 68.377
R276 SUM.n5 SUM.n2 28.681
R277 SUM.n7 SUM.t5 26.595
R278 SUM.n7 SUM.t4 26.595
R279 SUM.n0 SUM.t7 26.595
R280 SUM.n0 SUM.t6 26.595
R281 SUM.n3 SUM.t3 24.923
R282 SUM.n3 SUM.t0 24.923
R283 SUM.n1 SUM.t2 24.923
R284 SUM.n1 SUM.t1 24.923
R285 SUM.n4 SUM 12.218
R286 SUM.n8 SUM 10.512
R287 SUM SUM.n5 9.503
R288 SUM.n6 SUM 7.951
R289 SUM.n6 SUM 5.236
R290 SUM.n5 SUM 3.684
R291 SUM SUM.n8 2.63
R292 SUM SUM.n4 0.969
R293 a_890_297.t0 a_890_297.t1 113.275
C0 COUT VPWR 0.46fF
C1 VGND B 0.11fF
C2 COUT VGND 0.32fF
C3 VPB VPWR 0.19fF
C4 A B 0.61fF
C5 VGND VPWR 0.23fF
C6 VPWR SUM 0.56fF
C7 VGND SUM 0.46fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__inv_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__inv_1 Y A VGND VPWR VNB VPB
X0 Y.t0 A.t0 VGND.t0 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 Y.t1 A.t1 VPWR.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
R0 A.n0 A.t1 230.574
R1 A.n0 A.t0 158.274
R2 A A.n0 82.666
R3 VGND VGND.t0 118.397
R4 Y.n0 Y.t1 137.914
R5 Y Y.t0 106.634
R6 Y Y.n0 2.226
R7 Y.n0 Y 1.551
R8 VNB VNB.t0 7390.78
R9 VPWR VPWR.t0 164.986
R10 VPB VPB.t0 350.852
C0 Y VGND 0.17fF
C1 VPWR Y 0.22fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__inv_2.ext - technology: sky130A

.subckt sky130_fd_sc_hd__inv_2 A Y VPWR VGND VNB VPB
X0 Y.t1 A.t0 VPWR.t1 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 VGND.t1 A.t1 Y.t3 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 Y.t2 A.t2 VGND.t0 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 VPWR.t0 A.t3 Y.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
R0 A.n0 A.t3 212.079
R1 A.n1 A.t0 212.079
R2 A.n0 A.t1 139.779
R3 A.n1 A.t2 139.779
R4 A A.n1 113.072
R5 A.n1 A.n0 61.345
R6 VPWR.n0 VPWR.t0 162.171
R7 VPWR.n0 VPWR.t1 159.068
R8 VPWR VPWR.n0 0.126
R9 Y.n2 Y.n1 111.319
R10 Y Y.n0 50.466
R11 Y.n1 Y.t0 26.595
R12 Y.n1 Y.t1 26.595
R13 Y.n0 Y.t3 24.923
R14 Y.n0 Y.t2 24.923
R15 Y.n3 Y 11.264
R16 Y Y.n3 6.144
R17 Y.n3 Y 4.654
R18 Y Y.n2 2.048
R19 Y.n2 Y 1.551
R20 VPB.t1 VPB.t0 248.598
R21 VPB VPB.t1 198.286
R22 VGND.n0 VGND.t1 120.227
R23 VGND.n0 VGND.t0 117.585
R24 VGND VGND.n0 0.126
R25 VNB VNB.t0 6126.44
R26 VNB.t0 VNB.t1 2030.77
C0 Y VGND 0.27fF
C1 VPWR Y 0.38fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__inv_4.ext - technology: sky130A

.subckt sky130_fd_sc_hd__inv_4 Y A VPWR VGND VNB VPB
X0 VPWR.t3 A.t0 Y.t3 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 Y.t2 A.t1 VPWR.t2 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 Y.t7 A.t2 VGND.t3 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 VPWR.t1 A.t3 Y.t1 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 VGND.t2 A.t4 Y.t6 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 Y.t0 A.t5 VPWR.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 VGND.t1 A.t6 Y.t5 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 Y.t4 A.t7 VGND.t0 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
R0 A.n0 A.t0 212.079
R1 A.n1 A.t1 212.079
R2 A.n7 A.t3 212.079
R3 A.n3 A.t5 212.079
R4 A.n0 A.t6 139.779
R5 A.n1 A.t7 139.779
R6 A.n7 A.t4 139.779
R7 A.n3 A.t2 139.779
R8 A.n4 A.n3 112.515
R9 A A.n2 78.304
R10 A.n9 A.n8 76
R11 A.n6 A.n5 76
R12 A.n2 A.n0 30.672
R13 A.n2 A.n1 30.672
R14 A.n8 A.n7 30.672
R15 A.n7 A.n6 30.672
R16 A.n6 A.n3 30.672
R17 A A.n9 19.2
R18 A.n5 A 17.152
R19 A A.n4 17.152
R20 A.n5 A 6.4
R21 A.n4 A 6.4
R22 A.n9 A 4.352
R23 Y.n5 Y.n4 146.422
R24 Y.n2 Y.n0 144.087
R25 Y.n2 Y.n1 107.821
R26 Y.n5 Y.n3 107.247
R27 Y.n3 Y.t3 26.595
R28 Y.n3 Y.t2 26.595
R29 Y.n4 Y.t1 26.595
R30 Y.n4 Y.t0 26.595
R31 Y.n0 Y.t6 24.923
R32 Y.n0 Y.t7 24.923
R33 Y.n1 Y.t5 24.923
R34 Y.n1 Y.t4 24.923
R35 Y Y.n5 18.455
R36 Y.n6 Y 14.007
R37 Y.n6 Y.n2 12.088
R38 Y Y.n6 2.415
R39 VPWR.n2 VPWR.t3 588.709
R40 VPWR.n1 VPWR.n0 174.594
R41 VPWR.n5 VPWR.t0 151.12
R42 VPWR.n0 VPWR.t2 26.595
R43 VPWR.n0 VPWR.t1 26.595
R44 VPWR.n4 VPWR.n3 4.65
R45 VPWR.n6 VPWR.n5 4.65
R46 VPWR.n2 VPWR.n1 4.064
R47 VPWR.n4 VPWR.n2 0.208
R48 VPWR.n6 VPWR.n4 0.119
R49 VPWR VPWR.n6 0.022
R50 VPB.t2 VPB.t3 248.598
R51 VPB.t1 VPB.t2 248.598
R52 VPB.t0 VPB.t1 248.598
R53 VPB VPB.t0 221.962
R54 VGND.n2 VGND.t1 197.049
R55 VGND.n5 VGND.t3 193.93
R56 VGND.n1 VGND.n0 114.711
R57 VGND.n0 VGND.t0 24.923
R58 VGND.n0 VGND.t2 24.923
R59 VGND.n6 VGND.n5 4.65
R60 VGND.n4 VGND.n3 4.65
R61 VGND.n2 VGND.n1 4.064
R62 VGND.n4 VGND.n2 0.208
R63 VGND.n6 VGND.n4 0.119
R64 VGND VGND.n6 0.022
R65 VNB VNB.t3 6319.84
R66 VNB.t0 VNB.t1 2030.77
R67 VNB.t2 VNB.t0 2030.77
R68 VNB.t3 VNB.t2 2030.77
C0 VPWR Y 0.62fF
C1 A Y 0.48fF
C2 Y VGND 0.40fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__inv_6.ext - technology: sky130A

.subckt sky130_fd_sc_hd__inv_6 Y A VPWR VGND VNB VPB
X0 VPWR.t5 A.t0 Y.t5 VPB.t5 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 Y.t4 A.t1 VPWR.t4 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 Y.t11 A.t2 VGND.t5 VNB.t5 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 VPWR.t3 A.t3 Y.t3 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 Y.t2 A.t4 VPWR.t2 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 VPWR.t1 A.t5 Y.t1 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 Y.t10 A.t6 VGND.t4 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 Y.t9 A.t7 VGND.t3 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 Y.t0 A.t8 VPWR.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 VGND.t2 A.t9 Y.t8 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 VGND.t1 A.t10 Y.t7 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 VGND.t0 A.t11 Y.t6 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
R0 A.n0 A.t0 212.079
R1 A.n1 A.t1 212.079
R2 A.n9 A.t3 212.079
R3 A.n3 A.t4 212.079
R4 A.n4 A.t5 212.079
R5 A.n5 A.t8 212.079
R6 A.n0 A.t11 139.779
R7 A.n1 A.t2 139.779
R8 A.n9 A.t10 139.779
R9 A.n3 A.t7 139.779
R10 A.n4 A.t9 139.779
R11 A.n5 A.t6 139.779
R12 A.n6 A.n5 130.042
R13 A A.n2 78.304
R14 A.n11 A.n10 76
R15 A.n8 A.n7 76
R16 A A.n6 62.208
R17 A.n4 A.n3 61.345
R18 A.n5 A.n4 61.345
R19 A.n2 A.n0 42.357
R20 A.n9 A.n8 42.357
R21 A A.n11 19.2
R22 A.n2 A.n1 18.987
R23 A.n10 A.n9 18.987
R24 A.n8 A.n3 18.987
R25 A.n7 A 17.152
R26 A.n7 A 6.4
R27 A.n6 A 6.4
R28 A.n11 A 4.352
R29 Y.n3 Y.n2 175.197
R30 Y.n8 Y.n6 146.035
R31 Y.n3 Y.n1 115.464
R32 Y.n4 Y.n0 115.464
R33 Y.n8 Y.n7 107.635
R34 Y.n9 Y.n5 107.247
R35 Y.n4 Y.n3 59.733
R36 Y.n9 Y.n8 38.787
R37 Y.n5 Y.t5 26.595
R38 Y.n5 Y.t4 26.595
R39 Y.n6 Y.t1 26.595
R40 Y.n6 Y.t0 26.595
R41 Y.n7 Y.t3 26.595
R42 Y.n7 Y.t2 26.595
R43 Y.n2 Y.t8 24.923
R44 Y.n2 Y.t10 24.923
R45 Y.n1 Y.t7 24.923
R46 Y.n1 Y.t9 24.923
R47 Y.n0 Y.t6 24.923
R48 Y.n0 Y.t11 24.923
R49 Y.n10 Y.n4 18.133
R50 Y Y.n9 11.365
R51 Y.n10 Y 10.605
R52 Y Y.n10 1.828
R53 VPWR.n0 VPWR.t5 579.315
R54 VPWR.n13 VPWR.t0 181.903
R55 VPWR.n8 VPWR.n7 174.594
R56 VPWR.n2 VPWR.n1 174.594
R57 VPWR.n7 VPWR.t2 26.595
R58 VPWR.n7 VPWR.t1 26.595
R59 VPWR.n1 VPWR.t4 26.595
R60 VPWR.n1 VPWR.t3 26.595
R61 VPWR.n9 VPWR.n8 9.035
R62 VPWR.n4 VPWR.n3 4.65
R63 VPWR.n6 VPWR.n5 4.65
R64 VPWR.n10 VPWR.n9 4.65
R65 VPWR.n12 VPWR.n11 4.65
R66 VPWR.n14 VPWR.n13 4.65
R67 VPWR.n3 VPWR.n2 3.011
R68 VPWR.n4 VPWR.n0 0.941
R69 VPWR.n6 VPWR.n4 0.119
R70 VPWR.n10 VPWR.n6 0.119
R71 VPWR.n12 VPWR.n10 0.119
R72 VPWR.n14 VPWR.n12 0.119
R73 VPWR VPWR.n14 0.022
R74 VPB VPB.t0 292.99
R75 VPB.t4 VPB.t5 248.598
R76 VPB.t3 VPB.t4 248.598
R77 VPB.t2 VPB.t3 248.598
R78 VPB.t1 VPB.t2 248.598
R79 VPB.t0 VPB.t1 248.598
R80 VGND.n0 VGND.t0 193.19
R81 VGND.n13 VGND.t4 157.93
R82 VGND.n2 VGND.n1 114.711
R83 VGND.n8 VGND.n7 114.711
R84 VGND.n1 VGND.t5 24.923
R85 VGND.n1 VGND.t1 24.923
R86 VGND.n7 VGND.t3 24.923
R87 VGND.n7 VGND.t2 24.923
R88 VGND.n9 VGND.n8 9.035
R89 VGND.n14 VGND.n13 4.65
R90 VGND.n4 VGND.n3 4.65
R91 VGND.n6 VGND.n5 4.65
R92 VGND.n10 VGND.n9 4.65
R93 VGND.n12 VGND.n11 4.65
R94 VGND.n3 VGND.n2 3.011
R95 VGND.n4 VGND.n0 0.895
R96 VGND.n6 VGND.n4 0.119
R97 VGND.n10 VGND.n6 0.119
R98 VGND.n12 VGND.n10 0.119
R99 VGND.n14 VGND.n12 0.119
R100 VGND VGND.n14 0.022
R101 VNB VNB.t4 6900.06
R102 VNB.t5 VNB.t0 2030.77
R103 VNB.t1 VNB.t5 2030.77
R104 VNB.t3 VNB.t1 2030.77
R105 VNB.t2 VNB.t3 2030.77
R106 VNB.t4 VNB.t2 2030.77
C0 Y VGND 0.46fF
C1 VPWR Y 0.89fF
C2 A Y 0.73fF
C3 A VPWR 0.12fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__inv_8.ext - technology: sky130A

.subckt sky130_fd_sc_hd__inv_8 A Y VGND VPWR VNB VPB
X0 VPWR.t7 A.t0 Y.t15 VPB.t7 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 Y.t14 A.t1 VPWR.t6 VPB.t6 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 Y.t7 A.t2 VGND.t7 VNB.t7 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 Y.t6 A.t3 VGND.t6 VNB.t6 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 VPWR.t5 A.t4 Y.t13 VPB.t5 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 Y.t12 A.t5 VPWR.t4 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 Y.t5 A.t6 VGND.t5 VNB.t5 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 VPWR.t3 A.t7 Y.t11 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 Y.t4 A.t8 VGND.t4 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 Y.t10 A.t9 VPWR.t2 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 VPWR.t1 A.t10 Y.t9 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 VGND.t3 A.t11 Y.t3 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 VGND.t2 A.t12 Y.t2 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 VGND.t1 A.t13 Y.t1 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14 Y.t8 A.t14 VPWR.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 VGND.t0 A.t15 Y.t0 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
R0 A.n0 A.t7 212.079
R1 A.n1 A.t9 212.079
R2 A.n17 A.t10 212.079
R3 A.n3 A.t14 212.079
R4 A.n12 A.t0 212.079
R5 A.n4 A.t1 212.079
R6 A.n7 A.t4 212.079
R7 A.n5 A.t5 212.079
R8 A.n0 A.t15 139.779
R9 A.n1 A.t3 139.779
R10 A.n17 A.t13 139.779
R11 A.n3 A.t2 139.779
R12 A.n12 A.t12 139.779
R13 A.n4 A.t8 139.779
R14 A.n7 A.t11 139.779
R15 A.n5 A.t6 139.779
R16 A.n6 A 87.264
R17 A A.n2 76
R18 A.n19 A.n18 76
R19 A.n16 A.n15 76
R20 A.n14 A.n13 76
R21 A.n11 A.n10 76
R22 A.n9 A.n8 76
R23 A.n2 A.n0 30.672
R24 A.n2 A.n1 30.672
R25 A.n18 A.n17 30.672
R26 A.n17 A.n16 30.672
R27 A.n16 A.n3 30.672
R28 A.n13 A.n3 30.672
R29 A.n13 A.n12 30.672
R30 A.n12 A.n11 30.672
R31 A.n11 A.n4 30.672
R32 A.n8 A.n4 30.672
R33 A.n8 A.n7 30.672
R34 A.n7 A.n6 30.672
R35 A.n6 A.n5 30.672
R36 A A.n19 21.504
R37 A.n15 A 19.456
R38 A A.n14 17.408
R39 A.n10 A 15.36
R40 A A.n9 13.312
R41 A.n9 A 10.24
R42 A.n10 A 8.192
R43 A.n14 A 6.144
R44 A.n15 A 4.096
R45 A.n19 A 2.048
R46 Y.n1 Y.n0 107.635
R47 Y.n3 Y.n2 107.635
R48 Y.n5 Y.n4 107.635
R49 Y.n7 Y.n6 107.635
R50 Y.n9 Y.n8 52.818
R51 Y.n11 Y.n10 52.818
R52 Y.n13 Y.n12 52.818
R53 Y.n15 Y.n14 52.818
R54 Y.n3 Y.n1 38.4
R55 Y.n5 Y.n3 38.4
R56 Y.n7 Y.n5 38.4
R57 Y Y.n1 36.446
R58 Y Y.n7 34.435
R59 Y.n11 Y.n9 34.357
R60 Y.n13 Y.n11 34.357
R61 Y.n15 Y.n13 34.357
R62 Y Y.n15 27.786
R63 Y.n0 Y.t13 26.595
R64 Y.n0 Y.t12 26.595
R65 Y.n2 Y.t15 26.595
R66 Y.n2 Y.t14 26.595
R67 Y.n4 Y.t9 26.595
R68 Y.n4 Y.t8 26.595
R69 Y.n6 Y.t11 26.595
R70 Y.n6 Y.t10 26.595
R71 Y.n9 Y 25.61
R72 Y.n8 Y.t0 24.923
R73 Y.n8 Y.t6 24.923
R74 Y.n10 Y.t1 24.923
R75 Y.n10 Y.t7 24.923
R76 Y.n12 Y.t2 24.923
R77 Y.n12 Y.t4 24.923
R78 Y.n14 Y.t3 24.923
R79 Y.n14 Y.t5 24.923
R80 VPWR.n2 VPWR.t3 196.567
R81 VPWR.n17 VPWR.t4 196.066
R82 VPWR.n12 VPWR.n11 174.594
R83 VPWR.n6 VPWR.n5 174.594
R84 VPWR.n1 VPWR.n0 174.594
R85 VPWR.n11 VPWR.t6 26.595
R86 VPWR.n11 VPWR.t5 26.595
R87 VPWR.n5 VPWR.t0 26.595
R88 VPWR.n5 VPWR.t7 26.595
R89 VPWR.n0 VPWR.t2 26.595
R90 VPWR.n0 VPWR.t1 26.595
R91 VPWR.n13 VPWR.n12 8.658
R92 VPWR.n2 VPWR.n1 7.442
R93 VPWR.n18 VPWR.n17 6.532
R94 VPWR.n4 VPWR.n3 4.65
R95 VPWR.n8 VPWR.n7 4.65
R96 VPWR.n10 VPWR.n9 4.65
R97 VPWR.n14 VPWR.n13 4.65
R98 VPWR.n16 VPWR.n15 4.65
R99 VPWR.n7 VPWR.n6 2.635
R100 VPWR.n4 VPWR.n2 0.217
R101 VPWR.n8 VPWR.n4 0.119
R102 VPWR.n10 VPWR.n8 0.119
R103 VPWR.n14 VPWR.n10 0.119
R104 VPWR.n16 VPWR.n14 0.119
R105 VPWR.n18 VPWR.n16 0.119
R106 VPWR VPWR.n18 0.022
R107 VPB VPB.t4 290.031
R108 VPB.t2 VPB.t3 248.598
R109 VPB.t1 VPB.t2 248.598
R110 VPB.t0 VPB.t1 248.598
R111 VPB.t7 VPB.t0 248.598
R112 VPB.t6 VPB.t7 248.598
R113 VPB.t5 VPB.t6 248.598
R114 VPB.t4 VPB.t5 248.598
R115 VGND.n2 VGND.t0 195.492
R116 VGND.n17 VGND.t5 194.65
R117 VGND.n1 VGND.n0 114.711
R118 VGND.n6 VGND.n5 114.711
R119 VGND.n12 VGND.n11 114.711
R120 VGND.n0 VGND.t6 24.923
R121 VGND.n0 VGND.t1 24.923
R122 VGND.n5 VGND.t7 24.923
R123 VGND.n5 VGND.t2 24.923
R124 VGND.n11 VGND.t4 24.923
R125 VGND.n11 VGND.t3 24.923
R126 VGND.n13 VGND.n12 8.658
R127 VGND.n2 VGND.n1 7.442
R128 VGND.n18 VGND.n17 6.532
R129 VGND.n4 VGND.n3 4.65
R130 VGND.n8 VGND.n7 4.65
R131 VGND.n10 VGND.n9 4.65
R132 VGND.n14 VGND.n13 4.65
R133 VGND.n16 VGND.n15 4.65
R134 VGND.n7 VGND.n6 2.635
R135 VGND.n4 VGND.n2 0.217
R136 VGND.n8 VGND.n4 0.119
R137 VGND.n10 VGND.n8 0.119
R138 VGND.n14 VGND.n10 0.119
R139 VGND.n16 VGND.n14 0.119
R140 VGND.n18 VGND.n16 0.119
R141 VGND VGND.n18 0.022
R142 VNB VNB.t5 6916.79
R143 VNB.t6 VNB.t0 2030.77
R144 VNB.t1 VNB.t6 2030.77
R145 VNB.t7 VNB.t1 2030.77
R146 VNB.t2 VNB.t7 2030.77
R147 VNB.t4 VNB.t2 2030.77
R148 VNB.t3 VNB.t4 2030.77
R149 VNB.t5 VNB.t3 2030.77
C0 Y VGND 0.98fF
C1 VPWR Y 1.40fF
C2 A Y 1.35fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__inv_12.ext - technology: sky130A

.subckt sky130_fd_sc_hd__inv_12 A Y VGND VPWR VNB VPB
X0 VPWR.t11 A.t0 Y.t10 VPB.t11 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 Y.t9 A.t1 VPWR.t10 VPB.t10 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 Y.t8 A.t2 VPWR.t9 VPB.t9 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 VPWR.t8 A.t3 Y.t7 VPB.t8 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 Y.t22 A.t4 VGND.t11 VNB.t11 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 Y.t21 A.t5 VGND.t10 VNB.t10 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 VPWR.t7 A.t6 Y.t6 VPB.t7 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 VPWR.t6 A.t7 Y.t5 VPB.t6 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 Y.t20 A.t8 VGND.t9 VNB.t9 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 Y.t19 A.t9 VGND.t8 VNB.t8 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 Y.t4 A.t10 VPWR.t5 VPB.t5 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 VGND.t7 A.t11 Y.t18 VNB.t7 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 VGND.t6 A.t12 Y.t17 VNB.t6 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 Y.t3 A.t13 VPWR.t4 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14 Y.t16 A.t14 VGND.t5 VNB.t5 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X15 VPWR.t3 A.t15 Y.t2 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16 Y.t15 A.t16 VGND.t4 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X17 Y.t1 A.t17 VPWR.t2 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X18 VPWR.t1 A.t18 Y.t0 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X19 VGND.t3 A.t19 Y.t14 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X20 VGND.t2 A.t20 Y.t13 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X21 VGND.t1 A.t21 Y.t12 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X22 Y.t23 A.t22 VPWR.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X23 VGND.t0 A.t23 Y.t11 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
R0 A.n23 A.t3 212.079
R1 A.n22 A.t2 212.079
R2 A.n27 A.t7 212.079
R3 A.n28 A.t10 212.079
R4 A.n19 A.t15 212.079
R5 A.n0 A.t17 212.079
R6 A.n15 A.t18 212.079
R7 A.n1 A.t22 212.079
R8 A.n10 A.t0 212.079
R9 A.n2 A.t1 212.079
R10 A.n5 A.t6 212.079
R11 A.n3 A.t13 212.079
R12 A.n23 A.t11 139.779
R13 A.n22 A.t9 139.779
R14 A.n27 A.t12 139.779
R15 A.n28 A.t8 139.779
R16 A.n19 A.t23 139.779
R17 A.n0 A.t5 139.779
R18 A.n15 A.t21 139.779
R19 A.n1 A.t4 139.779
R20 A.n10 A.t20 139.779
R21 A.n2 A.t16 139.779
R22 A.n5 A.t19 139.779
R23 A.n3 A.t14 139.779
R24 A.n4 A 87.264
R25 A A.n24 78.048
R26 A.n26 A.n25 76
R27 A A.n29 76
R28 A.n21 A.n20 76
R29 A.n18 A 76
R30 A.n17 A.n16 76
R31 A.n14 A.n13 76
R32 A.n12 A.n11 76
R33 A.n9 A.n8 76
R34 A.n7 A.n6 76
R35 A.n24 A.n23 30.672
R36 A.n24 A.n22 30.672
R37 A.n26 A.n22 30.672
R38 A.n27 A.n26 30.672
R39 A.n29 A.n27 30.672
R40 A.n29 A.n28 30.672
R41 A.n20 A.n19 30.672
R42 A.n19 A.n18 30.672
R43 A.n18 A.n0 30.672
R44 A.n16 A.n0 30.672
R45 A.n16 A.n15 30.672
R46 A.n15 A.n14 30.672
R47 A.n14 A.n1 30.672
R48 A.n11 A.n1 30.672
R49 A.n11 A.n10 30.672
R50 A.n10 A.n9 30.672
R51 A.n9 A.n2 30.672
R52 A.n6 A.n2 30.672
R53 A.n6 A.n5 30.672
R54 A.n5 A.n4 30.672
R55 A.n4 A.n3 30.672
R56 A A.n21 21.504
R57 A A.n17 21.504
R58 A.n25 A 19.456
R59 A.n13 A 19.456
R60 A A.n12 17.408
R61 A.n8 A 15.36
R62 A A.n7 13.312
R63 A.n7 A 10.24
R64 A.n8 A 8.192
R65 A.n12 A 6.144
R66 A.n13 A 4.096
R67 A.n25 A 2.048
R68 A.n21 A 2.048
R69 A.n17 A 2.048
R70 Y.n1 Y.n0 107.635
R71 Y.n3 Y.n2 107.635
R72 Y.n5 Y.n4 107.635
R73 Y.n7 Y.n6 107.635
R74 Y.n9 Y.n8 107.635
R75 Y.n11 Y.n10 107.635
R76 Y.n13 Y.n12 52.818
R77 Y.n15 Y.n14 52.818
R78 Y.n17 Y.n16 52.818
R79 Y.n19 Y.n18 52.818
R80 Y.n21 Y.n20 52.818
R81 Y.n23 Y.n22 52.818
R82 Y Y.n11 42.594
R83 Y.n3 Y.n1 38.4
R84 Y.n5 Y.n3 38.4
R85 Y.n7 Y.n5 38.4
R86 Y.n9 Y.n7 38.4
R87 Y.n11 Y.n9 38.4
R88 Y.n15 Y.n13 34.357
R89 Y.n17 Y.n15 34.357
R90 Y.n19 Y.n17 34.357
R91 Y.n21 Y.n19 34.357
R92 Y.n23 Y.n21 34.357
R93 Y.n13 Y 33.356
R94 Y Y.n1 27.105
R95 Y.n0 Y.t6 26.595
R96 Y.n0 Y.t3 26.595
R97 Y.n2 Y.t10 26.595
R98 Y.n2 Y.t9 26.595
R99 Y.n4 Y.t0 26.595
R100 Y.n4 Y.t23 26.595
R101 Y.n6 Y.t2 26.595
R102 Y.n6 Y.t1 26.595
R103 Y.n8 Y.t5 26.595
R104 Y.n8 Y.t4 26.595
R105 Y.n10 Y.t7 26.595
R106 Y.n10 Y.t8 26.595
R107 Y.n12 Y.t18 24.923
R108 Y.n12 Y.t19 24.923
R109 Y.n14 Y.t17 24.923
R110 Y.n14 Y.t20 24.923
R111 Y.n16 Y.t11 24.923
R112 Y.n16 Y.t21 24.923
R113 Y.n18 Y.t12 24.923
R114 Y.n18 Y.t22 24.923
R115 Y.n20 Y.t13 24.923
R116 Y.n20 Y.t15 24.923
R117 Y.n22 Y.t14 24.923
R118 Y.n22 Y.t16 24.923
R119 Y Y.n23 20.336
R120 VPWR.n2 VPWR.t8 244.522
R121 VPWR.n29 VPWR.t4 196.066
R122 VPWR.n24 VPWR.n23 174.594
R123 VPWR.n18 VPWR.n17 174.594
R124 VPWR.n12 VPWR.n11 174.594
R125 VPWR.n6 VPWR.n5 174.594
R126 VPWR.n1 VPWR.n0 174.594
R127 VPWR.n23 VPWR.t10 26.595
R128 VPWR.n23 VPWR.t7 26.595
R129 VPWR.n17 VPWR.t0 26.595
R130 VPWR.n17 VPWR.t11 26.595
R131 VPWR.n11 VPWR.t2 26.595
R132 VPWR.n11 VPWR.t1 26.595
R133 VPWR.n5 VPWR.t5 26.595
R134 VPWR.n5 VPWR.t3 26.595
R135 VPWR.n0 VPWR.t9 26.595
R136 VPWR.n0 VPWR.t6 26.595
R137 VPWR.n2 VPWR.n1 19.493
R138 VPWR.n7 VPWR.n6 9.411
R139 VPWR.n25 VPWR.n24 8.658
R140 VPWR.n30 VPWR.n29 6.532
R141 VPWR.n4 VPWR.n3 4.65
R142 VPWR.n8 VPWR.n7 4.65
R143 VPWR.n10 VPWR.n9 4.65
R144 VPWR.n14 VPWR.n13 4.65
R145 VPWR.n16 VPWR.n15 4.65
R146 VPWR.n20 VPWR.n19 4.65
R147 VPWR.n22 VPWR.n21 4.65
R148 VPWR.n26 VPWR.n25 4.65
R149 VPWR.n28 VPWR.n27 4.65
R150 VPWR.n13 VPWR.n12 3.388
R151 VPWR.n19 VPWR.n18 2.635
R152 VPWR.n4 VPWR.n2 0.213
R153 VPWR.n8 VPWR.n4 0.119
R154 VPWR.n10 VPWR.n8 0.119
R155 VPWR.n14 VPWR.n10 0.119
R156 VPWR.n16 VPWR.n14 0.119
R157 VPWR.n20 VPWR.n16 0.119
R158 VPWR.n22 VPWR.n20 0.119
R159 VPWR.n26 VPWR.n22 0.119
R160 VPWR.n28 VPWR.n26 0.119
R161 VPWR.n30 VPWR.n28 0.119
R162 VPWR VPWR.n30 0.022
R163 VPB VPB.t4 290.031
R164 VPB.t9 VPB.t8 248.598
R165 VPB.t6 VPB.t9 248.598
R166 VPB.t5 VPB.t6 248.598
R167 VPB.t3 VPB.t5 248.598
R168 VPB.t2 VPB.t3 248.598
R169 VPB.t1 VPB.t2 248.598
R170 VPB.t0 VPB.t1 248.598
R171 VPB.t11 VPB.t0 248.598
R172 VPB.t10 VPB.t11 248.598
R173 VPB.t7 VPB.t10 248.598
R174 VPB.t4 VPB.t7 248.598
R175 VGND.n29 VGND.t5 194.65
R176 VGND.n2 VGND.t7 182.809
R177 VGND.n1 VGND.n0 114.711
R178 VGND.n6 VGND.n5 114.711
R179 VGND.n12 VGND.n11 114.711
R180 VGND.n18 VGND.n17 114.711
R181 VGND.n24 VGND.n23 114.711
R182 VGND.n0 VGND.t8 24.923
R183 VGND.n0 VGND.t6 24.923
R184 VGND.n5 VGND.t9 24.923
R185 VGND.n5 VGND.t0 24.923
R186 VGND.n11 VGND.t10 24.923
R187 VGND.n11 VGND.t1 24.923
R188 VGND.n17 VGND.t11 24.923
R189 VGND.n17 VGND.t2 24.923
R190 VGND.n23 VGND.t4 24.923
R191 VGND.n23 VGND.t3 24.923
R192 VGND.n2 VGND.n1 19.493
R193 VGND.n7 VGND.n6 9.411
R194 VGND.n25 VGND.n24 8.658
R195 VGND.n30 VGND.n29 6.532
R196 VGND.n4 VGND.n3 4.65
R197 VGND.n8 VGND.n7 4.65
R198 VGND.n10 VGND.n9 4.65
R199 VGND.n14 VGND.n13 4.65
R200 VGND.n16 VGND.n15 4.65
R201 VGND.n20 VGND.n19 4.65
R202 VGND.n22 VGND.n21 4.65
R203 VGND.n26 VGND.n25 4.65
R204 VGND.n28 VGND.n27 4.65
R205 VGND.n13 VGND.n12 3.388
R206 VGND.n19 VGND.n18 2.635
R207 VGND.n4 VGND.n2 0.213
R208 VGND.n8 VGND.n4 0.119
R209 VGND.n10 VGND.n8 0.119
R210 VGND.n14 VGND.n10 0.119
R211 VGND.n16 VGND.n14 0.119
R212 VGND.n20 VGND.n16 0.119
R213 VGND.n22 VGND.n20 0.119
R214 VGND.n26 VGND.n22 0.119
R215 VGND.n28 VGND.n26 0.119
R216 VGND.n30 VGND.n28 0.119
R217 VGND VGND.n30 0.022
R218 VNB VNB.t5 6916.79
R219 VNB.t8 VNB.t7 2030.77
R220 VNB.t6 VNB.t8 2030.77
R221 VNB.t9 VNB.t6 2030.77
R222 VNB.t0 VNB.t9 2030.77
R223 VNB.t10 VNB.t0 2030.77
R224 VNB.t1 VNB.t10 2030.77
R225 VNB.t11 VNB.t1 2030.77
R226 VNB.t2 VNB.t11 2030.77
R227 VNB.t4 VNB.t2 2030.77
R228 VNB.t3 VNB.t4 2030.77
R229 VNB.t5 VNB.t3 2030.77
C0 Y VGND 1.38fF
C1 A Y 2.14fF
C2 VPB A 0.15fF
C3 VPWR Y 1.99fF
C4 VPB VPWR 0.12fF
C5 VPWR VGND 0.14fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__inv_16.ext - technology: sky130A

.subckt sky130_fd_sc_hd__inv_16 Y A VGND VPWR VNB VPB
X0 Y.t31 A.t0 VPWR.t1 VPB.t15 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 VPWR.t0 A.t1 Y.t30 VPB.t14 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 VGND.t15 A.t2 Y.t15 VNB.t15 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 Y.t29 A.t3 VPWR.t15 VPB.t13 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 VGND.t14 A.t4 Y.t14 VNB.t14 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 VGND.t13 A.t5 Y.t13 VNB.t13 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 Y.t28 A.t6 VPWR.t14 VPB.t12 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 VGND.t12 A.t7 Y.t12 VNB.t12 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 VPWR.t13 A.t8 Y.t27 VPB.t11 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 Y.t11 A.t9 VGND.t11 VNB.t11 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 VPWR.t12 A.t10 Y.t26 VPB.t10 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 Y.t10 A.t11 VGND.t10 VNB.t10 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 Y.t25 A.t12 VPWR.t11 VPB.t9 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13 VPWR.t10 A.t13 Y.t24 VPB.t8 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14 Y.t23 A.t14 VPWR.t9 VPB.t7 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 VGND.t9 A.t15 Y.t9 VNB.t9 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X16 Y.t8 A.t16 VGND.t8 VNB.t8 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X17 VGND.t7 A.t17 Y.t7 VNB.t7 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X18 VGND.t6 A.t18 Y.t6 VNB.t6 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X19 Y.t22 A.t19 VPWR.t8 VPB.t6 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X20 VGND.t5 A.t20 Y.t5 VNB.t5 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X21 Y.t21 A.t21 VPWR.t7 VPB.t5 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X22 VPWR.t6 A.t22 Y.t20 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X23 VPWR.t5 A.t23 Y.t19 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X24 VPWR.t4 A.t24 Y.t18 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X25 Y.t4 A.t25 VGND.t4 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X26 Y.t17 A.t26 VPWR.t3 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X27 Y.t3 A.t27 VGND.t3 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X28 Y.t2 A.t28 VGND.t2 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X29 Y.t1 A.t29 VGND.t1 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X30 VPWR.t2 A.t30 Y.t16 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X31 Y.t0 A.t31 VGND.t0 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
R0 A.n0 A.t1 212.079
R1 A.n1 A.t3 212.079
R2 A.n2 A.t8 212.079
R3 A.n3 A.t14 212.079
R4 A.n5 A.t22 212.079
R5 A.n6 A.t21 212.079
R6 A.n9 A.t24 212.079
R7 A.n10 A.t26 212.079
R8 A.n25 A.t30 212.079
R9 A.n24 A.t0 212.079
R10 A.n11 A.t10 212.079
R11 A.n12 A.t12 212.079
R12 A.n14 A.t13 212.079
R13 A.n15 A.t19 212.079
R14 A.n18 A.t23 212.079
R15 A.n17 A.t6 212.079
R16 A.n0 A.t7 139.779
R17 A.n1 A.t11 139.779
R18 A.n2 A.t5 139.779
R19 A.n3 A.t27 139.779
R20 A.n5 A.t2 139.779
R21 A.n6 A.t31 139.779
R22 A.n9 A.t4 139.779
R23 A.n10 A.t29 139.779
R24 A.n25 A.t20 139.779
R25 A.n24 A.t28 139.779
R26 A.n11 A.t18 139.779
R27 A.n12 A.t25 139.779
R28 A.n14 A.t17 139.779
R29 A.n15 A.t9 139.779
R30 A.n18 A.t15 139.779
R31 A.n17 A.t16 139.779
R32 A.n17 A.n16 111.054
R33 A.n8 A.n7 76
R34 A.n27 A.n26 76
R35 A.n23 A.n22 76
R36 A.n20 A.n19 76
R37 A.n1 A.n0 61.345
R38 A.n2 A.n1 61.345
R39 A.n3 A.n2 61.345
R40 A.n6 A.n5 61.345
R41 A.n10 A.n9 61.345
R42 A.n25 A.n24 61.345
R43 A.n12 A.n11 61.345
R44 A.n15 A.n14 61.345
R45 A.n18 A.n17 61.345
R46 A.n22 A.n21 45.066
R47 A A.n20 43.733
R48 A.n27  41.6
R49 A.n16  41.066
R50 A.n4 A.n3 31.403
R51 A.n23 A.n11 31.403
R52 A.n8 A.n6 30.672
R53 A.n9 A.n8 30.672
R54 A.n26 A.n10 30.672
R55 A.n26 A.n25 30.672
R56 A.n13 A.n12 30.672
R57 A.n14 A.n13 30.672
R58 A.n19 A.n15 30.672
R59 A.n19 A.n18 30.672
R60 A.n5 A.n4 29.942
R61 A.n24 A.n23 29.942
R62 A.n7 A 12.8
R63 A.n16 A 8
R64 A A.n27 7.466
R65 A.n20  5.333
R66 A.n22  2.933
R67 A.n21 A 1.066
R68 VPWR.n2 VPWR.t0 205.068
R69 VPWR.n34 VPWR.n33 174.594
R70 VPWR.n28 VPWR.n27 174.594
R71 VPWR.n22 VPWR.n21 174.594
R72 VPWR.n16 VPWR.n15 174.594
R73 VPWR.n12 VPWR.n11 174.594
R74 VPWR.n6 VPWR.n5 174.594
R75 VPWR.n1 VPWR.n0 174.594
R76 VPWR.n39 VPWR.t14 158.114
R77 VPWR.n33 VPWR.t8 26.595
R78 VPWR.n33 VPWR.t5 26.595
R79 VPWR.n27 VPWR.t11 26.595
R80 VPWR.n27 VPWR.t10 26.595
R81 VPWR.n21 VPWR.t1 26.595
R82 VPWR.n21 VPWR.t12 26.595
R83 VPWR.n15 VPWR.t3 26.595
R84 VPWR.n15 VPWR.t2 26.595
R85 VPWR.n11 VPWR.t7 26.595
R86 VPWR.n11 VPWR.t4 26.595
R87 VPWR.n5 VPWR.t9 26.595
R88 VPWR.n5 VPWR.t6 26.595
R89 VPWR.n0 VPWR.t15 26.595
R90 VPWR.n0 VPWR.t13 26.595
R91 VPWR.n17 VPWR.n16 16.941
R92 VPWR.n13 VPWR.n12 11.67
R93 VPWR.n23 VPWR.n22 10.917
R94 VPWR.n7 VPWR.n6 5.647
R95 VPWR.n29 VPWR.n28 4.894
R96 VPWR.n4 VPWR.n3 4.65
R97 VPWR.n8 VPWR.n7 4.65
R98 VPWR.n10 VPWR.n9 4.65
R99 VPWR.n14 VPWR.n13 4.65
R100 VPWR.n18 VPWR.n17 4.65
R101 VPWR.n20 VPWR.n19 4.65
R102 VPWR.n24 VPWR.n23 4.65
R103 VPWR.n26 VPWR.n25 4.65
R104 VPWR.n30 VPWR.n29 4.65
R105 VPWR.n32 VPWR.n31 4.65
R106 VPWR.n36 VPWR.n35 4.65
R107 VPWR.n38 VPWR.n37 4.65
R108 VPWR.n40 VPWR.n39 4.65
R109 VPWR.n2 VPWR.n1 4.439
R110 VPWR.n35 VPWR.n34 1.129
R111 VPWR.n4 VPWR.n2 0.208
R112 VPWR.n8 VPWR.n4 0.119
R113 VPWR.n10 VPWR.n8 0.119
R114 VPWR.n14 VPWR.n10 0.119
R115 VPWR.n18 VPWR.n14 0.119
R116 VPWR.n20 VPWR.n18 0.119
R117 VPWR.n24 VPWR.n20 0.119
R118 VPWR.n26 VPWR.n24 0.119
R119 VPWR.n30 VPWR.n26 0.119
R120 VPWR.n32 VPWR.n30 0.119
R121 VPWR.n36 VPWR.n32 0.119
R122 VPWR.n38 VPWR.n36 0.119
R123 VPWR.n40 VPWR.n38 0.119
R124 VPWR VPWR.n40 0.022
R125 Y.n15 Y.n13 145.807
R126 Y.n15 Y.n14 107.407
R127 Y.n17 Y.n16 107.407
R128 Y.n19 Y.n18 107.407
R129 Y.n21 Y.n20 107.407
R130 Y.n23 Y.n22 107.407
R131 Y.n25 Y.n24 107.407
R132 Y.n27 Y.n26 107.407
R133 Y.n2 Y.n0 87.175
R134 Y.n2 Y.n1 52.818
R135 Y.n4 Y.n3 52.818
R136 Y.n6 Y.n5 52.818
R137 Y.n8 Y.n7 52.818
R138 Y.n10 Y.n9 52.818
R139 Y.n12 Y.n11 52.818
R140 Y Y.n29 51.073
R141 Y.n17 Y.n15 38.4
R142 Y.n19 Y.n17 38.4
R143 Y.n21 Y.n19 38.4
R144 Y.n23 Y.n21 38.4
R145 Y.n25 Y.n23 38.4
R146 Y.n27 Y.n25 38.4
R147 Y.n4 Y.n2 34.357
R148 Y.n6 Y.n4 34.357
R149 Y.n8 Y.n6 34.357
R150 Y.n10 Y.n8 34.357
R151 Y.n12 Y.n10 34.357
R152 Y.n28 Y.n12 34.357
R153 Y.n26 Y.t30 26.595
R154 Y.n26 Y.t29 26.595
R155 Y.n13 Y.t19 26.595
R156 Y.n13 Y.t28 26.595
R157 Y.n14 Y.t24 26.595
R158 Y.n14 Y.t22 26.595
R159 Y.n16 Y.t26 26.595
R160 Y.n16 Y.t25 26.595
R161 Y.n18 Y.t16 26.595
R162 Y.n18 Y.t31 26.595
R163 Y.n20 Y.t18 26.595
R164 Y.n20 Y.t17 26.595
R165 Y.n22 Y.t20 26.595
R166 Y.n22 Y.t21 26.595
R167 Y.n24 Y.t27 26.595
R168 Y.n24 Y.t23 26.595
R169 Y.n29 Y.t12 24.923
R170 Y.n29 Y.t10 24.923
R171 Y.n0 Y.t9 24.923
R172 Y.n0 Y.t8 24.923
R173 Y.n1 Y.t7 24.923
R174 Y.n1 Y.t11 24.923
R175 Y.n3 Y.t6 24.923
R176 Y.n3 Y.t4 24.923
R177 Y.n5 Y.t5 24.923
R178 Y.n5 Y.t2 24.923
R179 Y.n7 Y.t14 24.923
R180 Y.n7 Y.t1 24.923
R181 Y.n9 Y.t15 24.923
R182 Y.n9 Y.t0 24.923
R183 Y.n11 Y.t13 24.923
R184 Y.n11 Y.t3 24.923
R185 Y Y.n27 18.424
R186 Y.n28 Y 11.442
R187 Y Y.n28 1.745
R188 VPB.t13 VPB.t14 248.598
R189 VPB.t11 VPB.t13 248.598
R190 VPB.t7 VPB.t11 248.598
R191 VPB.t4 VPB.t7 248.598
R192 VPB.t5 VPB.t4 248.598
R193 VPB.t2 VPB.t5 248.598
R194 VPB.t1 VPB.t2 248.598
R195 VPB.t0 VPB.t1 248.598
R196 VPB.t15 VPB.t0 248.598
R197 VPB.t10 VPB.t15 248.598
R198 VPB.t9 VPB.t10 248.598
R199 VPB.t8 VPB.t9 248.598
R200 VPB.t6 VPB.t8 248.598
R201 VPB.t3 VPB.t6 248.598
R202 VPB.t12 VPB.t3 248.598
R203 VPB VPB.t12 230.841
R204 VGND.n2 VGND.t12 117.791
R205 VGND.n1 VGND.n0 114.711
R206 VGND.n6 VGND.n5 114.711
R207 VGND.n12 VGND.n11 114.711
R208 VGND.n16 VGND.n15 114.711
R209 VGND.n22 VGND.n21 114.711
R210 VGND.n28 VGND.n27 114.711
R211 VGND.n34 VGND.n33 114.711
R212 VGND.n39 VGND.t8 111.294
R213 VGND.n0 VGND.t10 24.923
R214 VGND.n0 VGND.t13 24.923
R215 VGND.n5 VGND.t3 24.923
R216 VGND.n5 VGND.t15 24.923
R217 VGND.n11 VGND.t0 24.923
R218 VGND.n11 VGND.t14 24.923
R219 VGND.n15 VGND.t1 24.923
R220 VGND.n15 VGND.t5 24.923
R221 VGND.n21 VGND.t2 24.923
R222 VGND.n21 VGND.t6 24.923
R223 VGND.n27 VGND.t4 24.923
R224 VGND.n27 VGND.t7 24.923
R225 VGND.n33 VGND.t11 24.923
R226 VGND.n33 VGND.t9 24.923
R227 VGND.n17 VGND.n16 16.941
R228 VGND.n13 VGND.n12 11.67
R229 VGND.n23 VGND.n22 10.917
R230 VGND.n7 VGND.n6 5.647
R231 VGND.n29 VGND.n28 4.894
R232 VGND.n40 VGND.n39 4.65
R233 VGND.n4 VGND.n3 4.65
R234 VGND.n8 VGND.n7 4.65
R235 VGND.n10 VGND.n9 4.65
R236 VGND.n14 VGND.n13 4.65
R237 VGND.n18 VGND.n17 4.65
R238 VGND.n20 VGND.n19 4.65
R239 VGND.n24 VGND.n23 4.65
R240 VGND.n26 VGND.n25 4.65
R241 VGND.n30 VGND.n29 4.65
R242 VGND.n32 VGND.n31 4.65
R243 VGND.n36 VGND.n35 4.65
R244 VGND.n38 VGND.n37 4.65
R245 VGND.n2 VGND.n1 4.439
R246 VGND.n35 VGND.n34 1.129
R247 VGND.n4 VGND.n2 0.208
R248 VGND.n8 VGND.n4 0.119
R249 VGND.n10 VGND.n8 0.119
R250 VGND.n14 VGND.n10 0.119
R251 VGND.n18 VGND.n14 0.119
R252 VGND.n20 VGND.n18 0.119
R253 VGND.n24 VGND.n20 0.119
R254 VGND.n26 VGND.n24 0.119
R255 VGND.n30 VGND.n26 0.119
R256 VGND.n32 VGND.n30 0.119
R257 VGND.n36 VGND.n32 0.119
R258 VGND.n38 VGND.n36 0.119
R259 VGND.n40 VGND.n38 0.119
R260 VGND VGND.n40 0.022
R261 VNB VNB.t8 6392.37
R262 VNB.t10 VNB.t12 2030.77
R263 VNB.t13 VNB.t10 2030.77
R264 VNB.t3 VNB.t13 2030.77
R265 VNB.t15 VNB.t3 2030.77
R266 VNB.t0 VNB.t15 2030.77
R267 VNB.t14 VNB.t0 2030.77
R268 VNB.t1 VNB.t14 2030.77
R269 VNB.t5 VNB.t1 2030.77
R270 VNB.t2 VNB.t5 2030.77
R271 VNB.t6 VNB.t2 2030.77
R272 VNB.t4 VNB.t6 2030.77
R273 VNB.t7 VNB.t4 2030.77
R274 VNB.t11 VNB.t7 2030.77
R275 VNB.t9 VNB.t11 2030.77
R276 VNB.t8 VNB.t9 2030.77
C0 VGND A 0.14fF
C1 VPB VPWR 0.15fF
C2 VGND VPWR 0.18fF
C3 A VPWR 0.17fF
C4 VGND Y 1.78fF
C5 A Y 1.82fF
C6 VPB A 0.22fF
C7 VPWR Y 2.60fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__lpflow_bleeder_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__lpflow_bleeder_1 VPB SHORT VPWR VGND VNB
X0 a_363_105.t0 SHORT.t0 a_291_105.t0 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X1 a_291_105.t1 SHORT.t1 a_219_105.t0 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X2 a_219_105.t1 SHORT.t2 a_147_105.t0 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X3 a_147_105.t1 SHORT.t3 VGND.t0 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X4 VPWR.t0 SHORT.t4 a_363_105.t1 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
R0 SHORT.n0 SHORT.t4 145.767
R1 SHORT.n6 SHORT.t3 101.949
R2 SHORT.n0 SHORT.t0 93.186
R3 SHORT.n3 SHORT.t2 93.186
R4 SHORT.n1 SHORT.t1 93.186
R5 SHORT.n5 SHORT.n4 76
R6 SHORT.n7 SHORT.n6 76
R7 SHORT.n5 SHORT.n2 36.386
R8 SHORT.n2 SHORT.n1 21.07
R9 SHORT.n2 SHORT.n0 19.655
R10 SHORT.n7 SHORT.n5 6.307
R11 SHORT.n4 SHORT.n3 5.842
R12 SHORT SHORT.n7 5.286
R13 a_291_105.t0 a_291_105.t1 70
R14 a_363_105.t0 a_363_105.t1 70
R15 VNB VNB.t1 18640.9
R16 VNB.t4 VNB.t0 2554.84
R17 VNB.t3 VNB.t4 2554.84
R18 VNB.t2 VNB.t3 2554.84
R19 VNB.t1 VNB.t2 2554.84
R20 a_219_105.t0 a_219_105.t1 70
R21 a_147_105.t0 a_147_105.t1 70
R22 VGND VGND.t0 169.529
R23 VPWR VPWR.t0 220.813
C0 SHORT VPWR 0.14fF
C1 SHORT VGND 0.14fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__lpflow_clkbufkapwr_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__lpflow_clkbufkapwr_1 KAPWR VGND VPWR X A VNB VPB
X0 KAPWR.t0 a_75_212.t2 X.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X1 a_75_212.t0 A.t0 VGND.t1 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X2 a_75_212.t1 A.t1 KAPWR.t1 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X3 VGND.t0 a_75_212.t3 X.t1 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
R0 a_75_212.t1 a_75_212.n1 260.844
R1 a_75_212.n0 a_75_212.t2 254.387
R2 a_75_212.n0 a_75_212.t3 211.007
R3 a_75_212.n1 a_75_212.t0 201.838
R4 a_75_212.n1 a_75_212.n0 76
R5 X.n1 X.t0 222.242
R6 X.n0 X.t1 123.653
R7 X X.n0 82.224
R8 X.n1 X 10.483
R9 X X.n1 5.504
R10 X.n0 X 5.169
R11 KAPWR.n0 KAPWR.t1 36.46
R12 KAPWR.n0 KAPWR.t0 35.128
R13 KAPWR KAPWR.n0 11.198
R14 VPB.t1 VPB.t0 260.436
R15 VPB VPB.t1 91.744
R16 A.n0 A.t1 260.32
R17 A.n0 A.t0 175.167
R18 A A.n0 78.133
R19 VGND VGND.n0 110.77
R20 VGND.n0 VGND.t1 33.461
R21 VGND.n0 VGND.t0 33.461
R22 VNB VNB.t1 6271.49
R23 VNB.t1 VNB.t0 2482.05
C0 VPWR KAPWR 0.55fF
C1 X KAPWR 0.10fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__lpflow_clkbufkapwr_2.ext - technology: sky130A

.subckt sky130_fd_sc_hd__lpflow_clkbufkapwr_2 A X KAPWR VGND VPWR VNB VPB
X0 KAPWR.t2 A.t0 a_27_47.t1 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 KAPWR.t1 a_27_47.t2 X.t3 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 VGND.t2 A.t1 a_27_47.t0 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3 X.t2 a_27_47.t3 KAPWR.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 X.t1 a_27_47.t4 VGND.t1 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 VGND.t0 a_27_47.t5 X.t0 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
R0 A.n0 A.t0 239.292
R1 A.n0 A.t1 171.059
R2 A A.n0 86.666
R3 a_27_47.t1 a_27_47.n3 261.044
R4 a_27_47.n3 a_27_47.t0 206.769
R5 a_27_47.n0 a_27_47.t3 189.586
R6 a_27_47.n0 a_27_47.t2 189.586
R7 a_27_47.n3 a_27_47.n2 139.081
R8 a_27_47.n1 a_27_47.t5 96.4
R9 a_27_47.n1 a_27_47.t4 96.4
R10 a_27_47.n2 a_27_47.n1 35.092
R11 a_27_47.n2 a_27_47.n0 19.871
R12 KAPWR.n0 KAPWR.t1 221.681
R13 KAPWR.n1 KAPWR.t0 36.445
R14 KAPWR.n2 KAPWR.t2 26.875
R15 KAPWR.n3 KAPWR.n2 8.636
R16 KAPWR.n5 KAPWR.n4 4.212
R17 KAPWR.n4 KAPWR.n3 2.235
R18 KAPWR KAPWR.n6 0.317
R19 KAPWR.n2 KAPWR.n1 0.248
R20 KAPWR.n5 KAPWR.n0 0.038
R21 KAPWR.n6 KAPWR.n5 0.002
R22 VPB.t2 VPB.t0 281.152
R23 VPB.t0 VPB.t1 248.598
R24 VPB VPB.t2 195.327
R25 X X.n0 342.551
R26 X X.n1 123.962
R27 X.n1 X.t0 38.571
R28 X.n1 X.t1 38.571
R29 X.n0 X.t3 26.595
R30 X.n0 X.t2 26.595
R31 VGND.n1 VGND.t0 150.351
R32 VGND.n1 VGND.n0 114.507
R33 VGND.n0 VGND.t1 52.857
R34 VGND.n0 VGND.t2 40
R35 VGND VGND.n1 0.214
R36 VNB VNB.t2 6502.94
R37 VNB.t2 VNB.t1 3073.53
R38 VNB.t1 VNB.t0 2717.65
C0 X VGND 0.17fF
C1 KAPWR VPWR 0.79fF
C2 KAPWR X 0.16fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__lpflow_clkbufkapwr_4.ext - technology: sky130A

.subckt sky130_fd_sc_hd__lpflow_clkbufkapwr_4 X A KAPWR VGND VPWR VNB VPB
X0 KAPWR.t4 A.t0 a_27_47.t1 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 VGND.t3 a_27_47.t2 X.t3 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 VGND.t2 a_27_47.t3 X.t2 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3 X.t7 a_27_47.t4 KAPWR.t3 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 X.t1 a_27_47.t5 VGND.t1 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 VGND.t4 A.t1 a_27_47.t0 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 KAPWR.t2 a_27_47.t6 X.t6 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 X.t0 a_27_47.t7 VGND.t0 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 X.t5 a_27_47.t8 KAPWR.t1 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 KAPWR.t0 a_27_47.t9 X.t4 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
R0 A.n0 A.t0 238.589
R1 A.n0 A.t1 203.243
R2 A A.n0 78.011
R3 a_27_47.t1 a_27_47.n11 271.613
R4 a_27_47.n8 a_27_47.t8 223.188
R5 a_27_47.n0 a_27_47.t6 221.719
R6 a_27_47.n3 a_27_47.t4 221.719
R7 a_27_47.n7 a_27_47.t9 221.719
R8 a_27_47.n11 a_27_47.t0 212.086
R9 a_27_47.n0 a_27_47.t2 185.378
R10 a_27_47.n8 a_27_47.t7 184.766
R11 a_27_47.n6 a_27_47.t3 184.766
R12 a_27_47.n2 a_27_47.t5 184.766
R13 a_27_47.n5 a_27_47.n1 101.6
R14 a_27_47.n11 a_27_47.n10 85.457
R15 a_27_47.n5 a_27_47.n4 76
R16 a_27_47.n10 a_27_47.n9 76
R17 a_27_47.n1 a_27_47.n0 56.963
R18 a_27_47.n9 a_27_47.n8 49.076
R19 a_27_47.n4 a_27_47.n3 41.189
R20 a_27_47.n10 a_27_47.n5 25.6
R21 a_27_47.n9 a_27_47.n7 25.414
R22 a_27_47.n3 a_27_47.n2 0.876
R23 a_27_47.n7 a_27_47.n6 0.876
R24 KAPWR.n1 KAPWR.t2 40.604
R25 KAPWR.n3 KAPWR.t1 37.43
R26 KAPWR.n0 KAPWR.t3 28.783
R27 KAPWR.n4 KAPWR.t4 26.875
R28 KAPWR.n0 KAPWR.t0 25.914
R29 KAPWR.n1 KAPWR.n0 11.256
R30 KAPWR.n5 KAPWR.n4 8.637
R31 KAPWR.n7 KAPWR.n6 4.465
R32 KAPWR.n6 KAPWR.n5 2.894
R33 KAPWR.n2 KAPWR.n1 0.466
R34 KAPWR KAPWR.n8 0.301
R35 KAPWR.n4 KAPWR.n3 0.248
R36 KAPWR.n7 KAPWR.n2 0.038
R37 KAPWR.n8 KAPWR.n7 0.002
R38 VPB.t4 VPB.t1 284.112
R39 VPB.t3 VPB.t2 254.517
R40 VPB.t0 VPB.t3 254.517
R41 VPB.t1 VPB.t0 254.517
R42 VPB VPB.t4 195.327
R43 X.n5 X.n3 400.623
R44 X.n2 X.n0 151.126
R45 X.n2 X.n1 107.761
R46 X.n5 X.n4 99.179
R47 X.n0 X.t2 40
R48 X.n0 X.t0 40
R49 X.n1 X.t3 40
R50 X.n1 X.t1 40
R51 X.n3 X.t4 27.58
R52 X.n3 X.t5 27.58
R53 X.n4 X.t6 27.58
R54 X.n4 X.t7 27.58
R55 X X.n6 19.259
R56 X.n6 X.n5 13.263
R57 X.n7 X 9.007
R58 X.n7 X.n2 6.776
R59 X.n6 X 2.707
R60 X X.n7 1.738
R61 VGND.n2 VGND.t3 154.76
R62 VGND.n1 VGND.n0 112.578
R63 VGND.n6 VGND.n5 111.118
R64 VGND.n5 VGND.t0 55.714
R65 VGND.n0 VGND.t1 40
R66 VGND.n0 VGND.t2 40
R67 VGND.n5 VGND.t4 40
R68 VGND.n4 VGND.n3 4.65
R69 VGND.n7 VGND.n6 3.996
R70 VGND.n2 VGND.n1 3.901
R71 VGND.n4 VGND.n2 0.238
R72 VGND.n7 VGND.n4 0.136
R73 VGND VGND.n7 0.125
R74 VNB VNB.t4 6502.94
R75 VNB.t4 VNB.t0 3138.24
R76 VNB.t1 VNB.t3 2782.35
R77 VNB.t2 VNB.t1 2782.35
R78 VNB.t0 VNB.t2 2782.35
C0 X VPWR 0.11fF
C1 X VGND 0.35fF
C2 KAPWR VPWR 1.20fF
C3 KAPWR X 0.39fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__lpflow_clkbufkapwr_8.ext - technology: sky130A

.subckt sky130_fd_sc_hd__lpflow_clkbufkapwr_8 X A KAPWR VGND VPWR VNB VPB
X0 KAPWR.t9 A.t0 a_110_47.t3 VPB.t9 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 KAPWR.t7 a_110_47.t4 X.t15 VPB.t7 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 X.t14 a_110_47.t5 KAPWR.t6 VPB.t6 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 a_110_47.t2 A.t1 KAPWR.t8 VPB.t8 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 X.t7 a_110_47.t6 VGND.t7 VNB.t7 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 X.t13 a_110_47.t7 KAPWR.t5 VPB.t5 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 VGND.t6 a_110_47.t8 X.t6 VNB.t6 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7 KAPWR.t4 a_110_47.t9 X.t12 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 VGND.t9 A.t2 a_110_47.t1 VNB.t9 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9 VGND.t5 a_110_47.t10 X.t5 VNB.t5 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10 a_110_47.t0 A.t3 VGND.t8 VNB.t8 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11 KAPWR.t3 a_110_47.t11 X.t11 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 X.t10 a_110_47.t12 KAPWR.t2 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13 VGND.t4 a_110_47.t13 X.t4 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14 VGND.t3 a_110_47.t14 X.t3 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15 X.t9 a_110_47.t15 KAPWR.t1 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16 X.t2 a_110_47.t16 VGND.t2 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17 KAPWR.t0 a_110_47.t17 X.t8 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X18 X.t1 a_110_47.t18 VGND.t1 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19 X.t0 a_110_47.t19 VGND.t0 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
R0 A.n0 A.t0 184.766
R1 A.n1 A.t1 184.766
R2 A.n0 A.t2 146.206
R3 A.n1 A.t3 146.206
R4 A A.n1 97.608
R5 A.n1 A.n0 40.639
R6 a_110_47.n1 a_110_47.t17 212.079
R7 a_110_47.n2 a_110_47.t12 212.079
R8 a_110_47.n3 a_110_47.t9 212.079
R9 a_110_47.n5 a_110_47.t5 212.079
R10 a_110_47.n8 a_110_47.t4 212.079
R11 a_110_47.n11 a_110_47.t15 212.079
R12 a_110_47.n16 a_110_47.t11 212.079
R13 a_110_47.n17 a_110_47.t7 212.079
R14 a_110_47.n21 a_110_47.n20 170.244
R15 a_110_47.n1 a_110_47.t10 162.273
R16 a_110_47.n2 a_110_47.t16 162.273
R17 a_110_47.n3 a_110_47.t13 162.273
R18 a_110_47.n5 a_110_47.t18 162.273
R19 a_110_47.n8 a_110_47.t14 162.273
R20 a_110_47.n11 a_110_47.t19 162.273
R21 a_110_47.n16 a_110_47.t8 162.273
R22 a_110_47.n17 a_110_47.t6 162.273
R23 a_110_47.n20 a_110_47.n0 124.756
R24 a_110_47.n7 a_110_47.n4 93.408
R25 a_110_47.n19 a_110_47.n18 76
R26 a_110_47.n7 a_110_47.n6 76
R27 a_110_47.n10 a_110_47.n9 76
R28 a_110_47.n13 a_110_47.n12 76
R29 a_110_47.n15 a_110_47.n14 76
R30 a_110_47.n2 a_110_47.n1 55.269
R31 a_110_47.n3 a_110_47.n2 55.269
R32 a_110_47.n20 a_110_47.n19 43.52
R33 a_110_47.n0 a_110_47.t1 40
R34 a_110_47.n0 a_110_47.t0 40
R35 a_110_47.n4 a_110_47.n3 30.848
R36 a_110_47.n18 a_110_47.n16 28.277
R37 a_110_47.n21 a_110_47.t3 27.58
R38 a_110_47.t2 a_110_47.n21 27.58
R39 a_110_47.n18 a_110_47.n17 26.992
R40 a_110_47.n6 a_110_47.n5 19.28
R41 a_110_47.n10 a_110_47.n7 17.408
R42 a_110_47.n13 a_110_47.n10 17.408
R43 a_110_47.n15 a_110_47.n13 17.408
R44 a_110_47.n19 a_110_47.n15 17.408
R45 a_110_47.n9 a_110_47.n8 7.712
R46 a_110_47.n12 a_110_47.n11 3.856
R47 KAPWR.n1 KAPWR.t0 182.85
R48 KAPWR.n8 KAPWR.t8 40.344
R49 KAPWR.n2 KAPWR.t6 28.781
R50 KAPWR.n4 KAPWR.t1 27.832
R51 KAPWR.n0 KAPWR.t2 27.827
R52 KAPWR.n6 KAPWR.t5 27.58
R53 KAPWR.n6 KAPWR.t9 27.58
R54 KAPWR.n0 KAPWR.t4 26.878
R55 KAPWR.n4 KAPWR.t3 26.871
R56 KAPWR.n2 KAPWR.t7 25.914
R57 KAPWR.n7 KAPWR.n6 12.867
R58 KAPWR.n1 KAPWR.n0 11.115
R59 KAPWR.n3 KAPWR.n2 11.062
R60 KAPWR.n5 KAPWR.n4 11.032
R61 KAPWR.n3 KAPWR.n1 0.523
R62 KAPWR.n8 KAPWR.n7 0.494
R63 KAPWR.n5 KAPWR.n3 0.491
R64 KAPWR.n7 KAPWR.n5 0.482
R65 KAPWR KAPWR.n8 0.055
R66 VPB.t2 VPB.t0 254.517
R67 VPB.t4 VPB.t2 254.517
R68 VPB.t6 VPB.t4 254.517
R69 VPB.t7 VPB.t6 254.517
R70 VPB.t1 VPB.t7 254.517
R71 VPB.t3 VPB.t1 254.517
R72 VPB.t5 VPB.t3 254.517
R73 VPB.t9 VPB.t5 254.517
R74 VPB.t8 VPB.t9 254.517
R75 VPB VPB.t8 195.327
R76 X.n7 X.n5 187.05
R77 X.n2 X.n0 156.137
R78 X.n7 X.n6 155.05
R79 X.n9 X.n8 155.05
R80 X.n11 X.n10 151.969
R81 X.n2 X.n1 110.961
R82 X.n4 X.n3 110.961
R83 X X.n13 107.171
R84 X.n4 X.n2 45.176
R85 X.n0 X.t6 40
R86 X.n0 X.t7 40
R87 X.n1 X.t3 40
R88 X.n1 X.t0 40
R89 X.n3 X.t4 40
R90 X.n3 X.t1 40
R91 X.n13 X.t5 40
R92 X.n13 X.t2 40
R93 X.n9 X.n7 32
R94 X.n5 X.t11 27.58
R95 X.n5 X.t13 27.58
R96 X.n6 X.t15 27.58
R97 X.n6 X.t9 27.58
R98 X.n8 X.t12 27.58
R99 X.n8 X.t14 27.58
R100 X.n10 X.t8 27.58
R101 X.n10 X.t10 27.58
R102 X.n12 X.n4 27.105
R103 X.n11 X.n9 19.2
R104 X.n12 X 3.76
R105 X X.n11 2.243
R106 X X.n12 0.725
R107 VGND.n2 VGND.t5 155.887
R108 VGND.n21 VGND.t8 152.353
R109 VGND.n17 VGND.n16 114.407
R110 VGND.n1 VGND.n0 112.192
R111 VGND.n6 VGND.n5 112.192
R112 VGND.n12 VGND.n11 112.192
R113 VGND.n0 VGND.t2 40
R114 VGND.n0 VGND.t4 40
R115 VGND.n5 VGND.t1 40
R116 VGND.n5 VGND.t3 40
R117 VGND.n11 VGND.t0 40
R118 VGND.n11 VGND.t6 40
R119 VGND.n16 VGND.t7 40
R120 VGND.n16 VGND.t9 40
R121 VGND.n2 VGND.n1 9.871
R122 VGND.n22 VGND.n21 4.65
R123 VGND.n4 VGND.n3 4.65
R124 VGND.n8 VGND.n7 4.65
R125 VGND.n10 VGND.n9 4.65
R126 VGND.n13 VGND.n12 4.65
R127 VGND.n15 VGND.n14 4.65
R128 VGND.n18 VGND.n17 4.65
R129 VGND.n20 VGND.n19 4.65
R130 VGND.n7 VGND.n6 1.505
R131 VGND.n4 VGND.n2 0.42
R132 VGND.n8 VGND.n4 0.119
R133 VGND.n10 VGND.n8 0.119
R134 VGND.n13 VGND.n10 0.119
R135 VGND.n15 VGND.n13 0.119
R136 VGND.n18 VGND.n15 0.119
R137 VGND.n20 VGND.n18 0.119
R138 VGND.n22 VGND.n20 0.119
R139 VGND VGND.n22 0.022
R140 VNB VNB.t8 6502.94
R141 VNB.t2 VNB.t5 2782.35
R142 VNB.t4 VNB.t2 2782.35
R143 VNB.t1 VNB.t4 2782.35
R144 VNB.t3 VNB.t1 2782.35
R145 VNB.t0 VNB.t3 2782.35
R146 VNB.t6 VNB.t0 2782.35
R147 VNB.t7 VNB.t6 2782.35
R148 VNB.t9 VNB.t7 2782.35
R149 VNB.t8 VNB.t9 2782.35
C0 X VPWR 0.25fF
C1 KAPWR X 0.99fF
C2 KAPWR VGND 0.13fF
C3 KAPWR VPWR 2.23fF
C4 X VGND 0.80fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__lpflow_clkbufkapwr_16.ext - technology: sky130A

.subckt sky130_fd_sc_hd__lpflow_clkbufkapwr_16 X A KAPWR VGND VPWR VNB VPB
X0 KAPWR.t3 A.t0 a_110_47.t3 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 KAPWR.t13 a_110_47.t8 X.t15 VPB.t19 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 X.t14 a_110_47.t9 KAPWR.t12 VPB.t18 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 X.t13 a_110_47.t10 KAPWR.t11 VPB.t17 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 KAPWR.t10 a_110_47.t11 X.t12 VPB.t16 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 KAPWR.t9 a_110_47.t12 X.t11 VPB.t15 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 a_110_47.t2 A.t1 KAPWR.t2 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 a_110_47.t7 A.t2 VGND.t3 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 VGND.t19 a_110_47.t13 X.t21 VNB.t19 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9 X.t20 a_110_47.t14 VGND.t18 VNB.t18 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10 VGND.t17 a_110_47.t15 X.t19 VNB.t17 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11 a_110_47.t1 A.t3 KAPWR.t1 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 VGND.t2 A.t4 a_110_47.t6 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13 VGND.t16 a_110_47.t16 X.t18 VNB.t16 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14 KAPWR.t8 a_110_47.t17 X.t10 VPB.t14 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 X.t9 a_110_47.t18 KAPWR.t7 VPB.t13 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16 VGND.t1 A.t5 a_110_47.t5 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17 VGND.t15 a_110_47.t19 X.t17 VNB.t15 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18 KAPWR.t6 a_110_47.t20 X.t8 VPB.t12 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X19 VGND.t14 a_110_47.t21 X.t16 VNB.t14 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20 X.t7 a_110_47.t22 KAPWR.t5 VPB.t11 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X21 a_110_47.t4 A.t6 VGND.t0 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22 KAPWR.t0 A.t7 a_110_47.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X23 KAPWR.t4 a_110_47.t23 X.t6 VPB.t10 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X24 KAPWR.t19 a_110_47.t24 X.t5 VPB.t9 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X25 VGND.t13 a_110_47.t25 X.t31 VNB.t13 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X26 X.t4 a_110_47.t26 KAPWR.t18 VPB.t8 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X27 VGND.t12 a_110_47.t27 X.t30 VNB.t12 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X28 VGND.t11 a_110_47.t28 X.t29 VNB.t11 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X29 X.t28 a_110_47.t29 VGND.t10 VNB.t10 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X30 X.t3 a_110_47.t30 KAPWR.t17 VPB.t7 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X31 X.t2 a_110_47.t31 KAPWR.t16 VPB.t6 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X32 X.t27 a_110_47.t32 VGND.t9 VNB.t9 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X33 KAPWR.t15 a_110_47.t33 X.t1 VPB.t5 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X34 X.t0 a_110_47.t34 KAPWR.t14 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X35 X.t26 a_110_47.t35 VGND.t8 VNB.t8 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X36 X.t25 a_110_47.t36 VGND.t7 VNB.t7 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X37 X.t24 a_110_47.t37 VGND.t6 VNB.t6 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X38 X.t23 a_110_47.t38 VGND.t5 VNB.t5 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X39 X.t22 a_110_47.t39 VGND.t4 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
R0 A.n0 A.t7 184.766
R1 A.n1 A.t3 184.766
R2 A.n2 A.t0 184.766
R3 A.n3 A.t1 184.766
R4 A.n0 A.t4 146.206
R5 A.n1 A.t2 146.206
R6 A.n2 A.t5 146.206
R7 A.n3 A.t6 146.206
R8 A A.n3 97.608
R9 A.n1 A.n0 40.639
R10 A.n2 A.n1 40.639
R11 A.n3 A.n2 40.639
R12 a_110_47.n1 a_110_47.t12 212.079
R13 a_110_47.n2 a_110_47.t34 212.079
R14 a_110_47.n3 a_110_47.t24 212.079
R15 a_110_47.n5 a_110_47.t18 212.079
R16 a_110_47.n8 a_110_47.t11 212.079
R17 a_110_47.n11 a_110_47.t30 212.079
R18 a_110_47.n14 a_110_47.t23 212.079
R19 a_110_47.n19 a_110_47.t22 212.079
R20 a_110_47.n22 a_110_47.t20 212.079
R21 a_110_47.n25 a_110_47.t10 212.079
R22 a_110_47.n28 a_110_47.t33 212.079
R23 a_110_47.n33 a_110_47.t26 212.079
R24 a_110_47.n36 a_110_47.t17 212.079
R25 a_110_47.n39 a_110_47.t9 212.079
R26 a_110_47.n44 a_110_47.t8 212.079
R27 a_110_47.n45 a_110_47.t31 212.079
R28 a_110_47.n1 a_110_47.t19 162.273
R29 a_110_47.n2 a_110_47.t29 162.273
R30 a_110_47.n3 a_110_47.t25 162.273
R31 a_110_47.n5 a_110_47.t35 162.273
R32 a_110_47.n8 a_110_47.t13 162.273
R33 a_110_47.n11 a_110_47.t37 162.273
R34 a_110_47.n14 a_110_47.t15 162.273
R35 a_110_47.n19 a_110_47.t39 162.273
R36 a_110_47.n22 a_110_47.t16 162.273
R37 a_110_47.n25 a_110_47.t14 162.273
R38 a_110_47.n28 a_110_47.t21 162.273
R39 a_110_47.n33 a_110_47.t32 162.273
R40 a_110_47.n36 a_110_47.t27 162.273
R41 a_110_47.n39 a_110_47.t36 162.273
R42 a_110_47.n44 a_110_47.t28 162.273
R43 a_110_47.n45 a_110_47.t38 162.273
R44 a_110_47.n51 a_110_47.n50 129.666
R45 a_110_47.n53 a_110_47.n52 128.898
R46 a_110_47.n51 a_110_47.n49 128.34
R47 a_110_47.n48 a_110_47.n0 124.756
R48 a_110_47.n7 a_110_47.n4 93.408
R49 a_110_47.n47 a_110_47.n46 76
R50 a_110_47.n7 a_110_47.n6 76
R51 a_110_47.n10 a_110_47.n9 76
R52 a_110_47.n13 a_110_47.n12 76
R53 a_110_47.n16 a_110_47.n15 76
R54 a_110_47.n18 a_110_47.n17 76
R55 a_110_47.n21 a_110_47.n20 76
R56 a_110_47.n24 a_110_47.n23 76
R57 a_110_47.n27 a_110_47.n26 76
R58 a_110_47.n30 a_110_47.n29 76
R59 a_110_47.n32 a_110_47.n31 76
R60 a_110_47.n35 a_110_47.n34 76
R61 a_110_47.n38 a_110_47.n37 76
R62 a_110_47.n41 a_110_47.n40 76
R63 a_110_47.n43 a_110_47.n42 76
R64 a_110_47.n2 a_110_47.n1 55.269
R65 a_110_47.n3 a_110_47.n2 55.269
R66 a_110_47.n48 a_110_47.n47 43.52
R67 a_110_47.n52 a_110_47.n51 43.264
R68 a_110_47.n49 a_110_47.t5 40
R69 a_110_47.n49 a_110_47.t4 40
R70 a_110_47.n0 a_110_47.t6 40
R71 a_110_47.n0 a_110_47.t7 40
R72 a_110_47.n4 a_110_47.n3 35.346
R73 a_110_47.n46 a_110_47.n44 28.277
R74 a_110_47.n50 a_110_47.t3 27.58
R75 a_110_47.n50 a_110_47.t2 27.58
R76 a_110_47.t0 a_110_47.n53 27.58
R77 a_110_47.n53 a_110_47.t1 27.58
R78 a_110_47.n46 a_110_47.n45 26.992
R79 a_110_47.n6 a_110_47.n5 23.778
R80 a_110_47.n20 a_110_47.n19 21.208
R81 a_110_47.n34 a_110_47.n33 19.28
R82 a_110_47.n10 a_110_47.n7 17.408
R83 a_110_47.n13 a_110_47.n10 17.408
R84 a_110_47.n16 a_110_47.n13 17.408
R85 a_110_47.n18 a_110_47.n16 17.408
R86 a_110_47.n21 a_110_47.n18 17.408
R87 a_110_47.n24 a_110_47.n21 17.408
R88 a_110_47.n27 a_110_47.n24 17.408
R89 a_110_47.n30 a_110_47.n27 17.408
R90 a_110_47.n32 a_110_47.n30 17.408
R91 a_110_47.n35 a_110_47.n32 17.408
R92 a_110_47.n38 a_110_47.n35 17.408
R93 a_110_47.n41 a_110_47.n38 17.408
R94 a_110_47.n43 a_110_47.n41 17.408
R95 a_110_47.n47 a_110_47.n43 17.408
R96 a_110_47.n29 a_110_47.n28 12.853
R97 a_110_47.n9 a_110_47.n8 12.21
R98 a_110_47.n15 a_110_47.n14 10.925
R99 a_110_47.n23 a_110_47.n22 10.282
R100 a_110_47.n37 a_110_47.n36 7.712
R101 a_110_47.n40 a_110_47.n39 3.856
R102 a_110_47.n26 a_110_47.n25 1.285
R103 a_110_47.n12 a_110_47.n11 0.642
R104 a_110_47.n52 a_110_47.n48 0.256
R105 KAPWR.n1 KAPWR.t9 182.874
R106 KAPWR.n23 KAPWR.t2 40.036
R107 KAPWR.n12 KAPWR.t12 28.781
R108 KAPWR.n0 KAPWR.t14 27.832
R109 KAPWR.n10 KAPWR.t18 27.827
R110 KAPWR.n8 KAPWR.t11 27.827
R111 KAPWR.n4 KAPWR.t17 27.827
R112 KAPWR.n21 KAPWR.t1 27.58
R113 KAPWR.n21 KAPWR.t3 27.58
R114 KAPWR.n6 KAPWR.t6 27.58
R115 KAPWR.n2 KAPWR.t7 27.58
R116 KAPWR.n2 KAPWR.t10 27.58
R117 KAPWR.n10 KAPWR.t8 26.878
R118 KAPWR.n8 KAPWR.t15 26.878
R119 KAPWR.n4 KAPWR.t4 26.878
R120 KAPWR.n0 KAPWR.t19 26.871
R121 KAPWR.n18 KAPWR.t0 26.595
R122 KAPWR.n6 KAPWR.t5 26.595
R123 KAPWR.n12 KAPWR.t13 25.914
R124 KAPWR.n16 KAPWR.t16 22.111
R125 KAPWR.n3 KAPWR.n2 12.576
R126 KAPWR.n7 KAPWR.n6 12.576
R127 KAPWR.n22 KAPWR.n21 12.457
R128 KAPWR.n11 KAPWR.n10 11.115
R129 KAPWR.n9 KAPWR.n8 11.115
R130 KAPWR.n5 KAPWR.n4 11.115
R131 KAPWR.n1 KAPWR.n0 11.088
R132 KAPWR.n13 KAPWR.n12 11.062
R133 KAPWR.n19 KAPWR.n18 9.3
R134 KAPWR.n17 KAPWR.n16 5.193
R135 KAPWR.n20 KAPWR.n19 4.641
R136 KAPWR.n15 KAPWR.n14 4.465
R137 KAPWR.n18 KAPWR.n17 0.985
R138 KAPWR.n13 KAPWR.n11 0.523
R139 KAPWR.n7 KAPWR.n5 0.503
R140 KAPWR.n11 KAPWR.n9 0.496
R141 KAPWR.n23 KAPWR.n22 0.494
R142 KAPWR.n5 KAPWR.n3 0.484
R143 KAPWR.n9 KAPWR.n7 0.484
R144 KAPWR.n3 KAPWR.n1 0.481
R145 KAPWR.n15 KAPWR.n13 0.481
R146 KAPWR.n22 KAPWR.n20 0.47
R147 KAPWR KAPWR.n23 0.057
R148 KAPWR.n20 KAPWR.n15 0.02
R149 VPB.t4 VPB.t15 254.517
R150 VPB.t9 VPB.t4 254.517
R151 VPB.t13 VPB.t9 254.517
R152 VPB.t16 VPB.t13 254.517
R153 VPB.t7 VPB.t16 254.517
R154 VPB.t10 VPB.t7 254.517
R155 VPB.t11 VPB.t10 254.517
R156 VPB.t17 VPB.t12 254.517
R157 VPB.t5 VPB.t17 254.517
R158 VPB.t8 VPB.t5 254.517
R159 VPB.t14 VPB.t8 254.517
R160 VPB.t18 VPB.t14 254.517
R161 VPB.t19 VPB.t18 254.517
R162 VPB.t6 VPB.t19 254.517
R163 VPB.t0 VPB.t6 254.517
R164 VPB.t1 VPB.t0 254.517
R165 VPB.t3 VPB.t1 254.517
R166 VPB.t2 VPB.t3 254.517
R167 VPB.t12 VPB.t11 251.557
R168 VPB VPB.t2 145.015
R169 X.n15 X.n13 192.158
R170 X.n2 X.n0 156.137
R171 X.n15 X.n14 155.885
R172 X.n17 X.n16 155.885
R173 X.n19 X.n18 155.885
R174 X.n21 X.n20 155.885
R175 X.n23 X.n22 155.885
R176 X.n25 X.n24 155.885
R177 X.n27 X.n26 153.087
R178 X.n2 X.n1 110.961
R179 X.n4 X.n3 110.961
R180 X.n8 X.n7 110.961
R181 X.n10 X.n9 110.961
R182 X.n12 X.n11 110.961
R183 X.n6 X.n5 109.954
R184 X X.n29 107.105
R185 X.n4 X.n2 45.176
R186 X.n10 X.n8 45.176
R187 X.n12 X.n10 45.176
R188 X.n6 X.n4 44.047
R189 X.n8 X.n6 44.047
R190 X.n0 X.t29 40
R191 X.n0 X.t23 40
R192 X.n1 X.t30 40
R193 X.n1 X.t25 40
R194 X.n3 X.t16 40
R195 X.n3 X.t27 40
R196 X.n5 X.t18 40
R197 X.n5 X.t20 40
R198 X.n7 X.t19 40
R199 X.n7 X.t22 40
R200 X.n9 X.t21 40
R201 X.n9 X.t24 40
R202 X.n11 X.t31 40
R203 X.n11 X.t26 40
R204 X.n29 X.t17 40
R205 X.n29 X.t28 40
R206 X.n17 X.n15 32
R207 X.n19 X.n17 32
R208 X.n23 X.n21 32
R209 X.n25 X.n23 32
R210 X.n21 X.n19 31.2
R211 X.n24 X.t5 27.58
R212 X.n24 X.t9 27.58
R213 X.n13 X.t15 27.58
R214 X.n13 X.t2 27.58
R215 X.n14 X.t10 27.58
R216 X.n14 X.t14 27.58
R217 X.n16 X.t1 27.58
R218 X.n16 X.t4 27.58
R219 X.n18 X.t8 27.58
R220 X.n18 X.t13 27.58
R221 X.n20 X.t6 27.58
R222 X.n20 X.t7 27.58
R223 X.n22 X.t12 27.58
R224 X.n22 X.t3 27.58
R225 X.n26 X.t11 27.58
R226 X.n26 X.t0 27.58
R227 X.n28 X.n12 13.176
R228 X.n27 X.n25 10.447
R229 X.n28 X 3.131
R230 X X.n27 1.757
R231 X X.n28 0.604
R232 VGND.n2 VGND.t15 153.42
R233 VGND.n46 VGND.t0 148.447
R234 VGND.n37 VGND.n36 114.407
R235 VGND.n42 VGND.n41 114.407
R236 VGND.n16 VGND.n15 113.397
R237 VGND.n21 VGND.n20 113.397
R238 VGND.n6 VGND.n5 112.98
R239 VGND.n11 VGND.n10 112.98
R240 VGND.n1 VGND.n0 112.192
R241 VGND.n25 VGND.n24 112.192
R242 VGND.n31 VGND.n30 112.192
R243 VGND.n0 VGND.t10 40
R244 VGND.n0 VGND.t13 40
R245 VGND.n5 VGND.t8 40
R246 VGND.n5 VGND.t19 40
R247 VGND.n10 VGND.t6 40
R248 VGND.n10 VGND.t17 40
R249 VGND.n15 VGND.t16 40
R250 VGND.n20 VGND.t18 40
R251 VGND.n20 VGND.t14 40
R252 VGND.n24 VGND.t9 40
R253 VGND.n24 VGND.t12 40
R254 VGND.n30 VGND.t7 40
R255 VGND.n30 VGND.t11 40
R256 VGND.n36 VGND.t5 40
R257 VGND.n36 VGND.t2 40
R258 VGND.n41 VGND.t3 40
R259 VGND.n41 VGND.t1 40
R260 VGND.n15 VGND.t4 38.571
R261 VGND.n26 VGND.n25 6.023
R262 VGND.n47 VGND.n46 4.65
R263 VGND.n4 VGND.n3 4.65
R264 VGND.n7 VGND.n6 4.65
R265 VGND.n9 VGND.n8 4.65
R266 VGND.n12 VGND.n11 4.65
R267 VGND.n14 VGND.n13 4.65
R268 VGND.n17 VGND.n16 4.65
R269 VGND.n19 VGND.n18 4.65
R270 VGND.n23 VGND.n22 4.65
R271 VGND.n27 VGND.n26 4.65
R272 VGND.n29 VGND.n28 4.65
R273 VGND.n33 VGND.n32 4.65
R274 VGND.n35 VGND.n34 4.65
R275 VGND.n38 VGND.n37 4.65
R276 VGND.n40 VGND.n39 4.65
R277 VGND.n43 VGND.n42 4.65
R278 VGND.n45 VGND.n44 4.65
R279 VGND.n22 VGND.n21 4.517
R280 VGND.n2 VGND.n1 3.953
R281 VGND.n32 VGND.n31 1.505
R282 VGND.n4 VGND.n2 0.242
R283 VGND.n7 VGND.n4 0.119
R284 VGND.n9 VGND.n7 0.119
R285 VGND.n12 VGND.n9 0.119
R286 VGND.n14 VGND.n12 0.119
R287 VGND.n17 VGND.n14 0.119
R288 VGND.n19 VGND.n17 0.119
R289 VGND.n23 VGND.n19 0.119
R290 VGND.n27 VGND.n23 0.119
R291 VGND.n29 VGND.n27 0.119
R292 VGND.n33 VGND.n29 0.119
R293 VGND.n35 VGND.n33 0.119
R294 VGND.n38 VGND.n35 0.119
R295 VGND.n40 VGND.n38 0.119
R296 VGND.n43 VGND.n40 0.119
R297 VGND.n45 VGND.n43 0.119
R298 VGND.n47 VGND.n45 0.119
R299 VGND VGND.n47 0.022
R300 VNB VNB.t0 4302.94
R301 VNB.t10 VNB.t15 2782.35
R302 VNB.t13 VNB.t10 2782.35
R303 VNB.t8 VNB.t13 2782.35
R304 VNB.t19 VNB.t8 2782.35
R305 VNB.t6 VNB.t19 2782.35
R306 VNB.t17 VNB.t6 2782.35
R307 VNB.t4 VNB.t17 2782.35
R308 VNB.t18 VNB.t16 2782.35
R309 VNB.t14 VNB.t18 2782.35
R310 VNB.t9 VNB.t14 2782.35
R311 VNB.t12 VNB.t9 2782.35
R312 VNB.t7 VNB.t12 2782.35
R313 VNB.t11 VNB.t7 2782.35
R314 VNB.t5 VNB.t11 2782.35
R315 VNB.t2 VNB.t5 2782.35
R316 VNB.t3 VNB.t2 2782.35
R317 VNB.t1 VNB.t3 2782.35
R318 VNB.t0 VNB.t1 2782.35
R319 VNB.t16 VNB.t4 2750
C0 KAPWR X 1.87fF
C1 VPB VPWR 0.17fF
C2 KAPWR VGND 0.25fF
C3 X VGND 1.57fF
C4 KAPWR VPWR 4.11fF
C5 X VPWR 0.49fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__lpflow_clkinvkapwr_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__lpflow_clkinvkapwr_1 Y A KAPWR VGND VPWR VNB VPB
X0 Y.t2 A.t0 KAPWR.t1 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X1 VGND.t0 A.t1 Y.t0 VNB sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 KAPWR.t0 A.t2 Y.t1 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
R0 A.n0 A.t2 231.907
R1 A.n1 A.t0 231.36
R2 A A.n1 207.012
R3 A.n0 A.t1 170.306
R4 A.n1 A.n0 54.062
R5 KAPWR.n2 KAPWR.t1 124.228
R6 KAPWR.n0 KAPWR.t0 120.497
R7 KAPWR.n3 KAPWR.n2 6.547
R8 KAPWR.n2 KAPWR.n1 0.721
R9 KAPWR.n4 KAPWR.n3 0.036
R10 KAPWR KAPWR.n4 0.024
R11 KAPWR.n3 KAPWR.n0 0.004
R12 Y Y.n0 198.633
R13 Y.n1 Y.t0 147.918
R14 Y.n0 Y.t1 31.66
R15 Y.n0 Y.t2 31.66
R16 Y Y.n1 6.191
R17 Y.n1 Y 0.024
R18 VPB.t1 VPB.t0 248.598
R19 VPB VPB.t1 192.367
R20 VGND VGND.t0 154.376
C0 KAPWR Y 0.27fF
C1 A Y 0.11fF
C2 KAPWR VPWR 0.61fF
C3 Y VGND 0.14fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__lpflow_clkinvkapwr_2.ext - technology: sky130A

.subckt sky130_fd_sc_hd__lpflow_clkinvkapwr_2 Y A KAPWR VPWR VGND VNB VPB
X0 Y.t2 A.t0 VGND.t1 VNB sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1 Y.t4 A.t1 KAPWR.t2 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 KAPWR.t1 A.t2 Y.t3 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 VGND.t0 A.t3 Y.t1 VNB sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 KAPWR.t0 A.t4 Y.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
R0 A.n0 A.t4 221.719
R1 A.n3 A.t1 221.719
R2 A.n7 A.t2 218.506
R3 A.n0 A.t3 189.05
R4 A.n2 A.t0 183.16
R5 A.n8 A.n7 105.086
R6 A.n6 A.n5 76
R7 A.n1 A.n0 63.278
R8 A.n6 A.n3 45.617
R9 A.n7 A.n6 27.957
R10 A.n5 A.n4 19.342
R11 A.n8 A 16.213
R12 A.n2 A.n1 10.328
R13 A A.n8 9.955
R14 A.n4 A 3.697
R15 A.n5 A 3.128
R16 A.n3 A.n2 2.582
R17 VGND.n0 VGND.t1 155.166
R18 VGND.n0 VGND.t0 150.198
R19 VGND VGND.n0 0.242
R20 Y.n2 Y.t3 297.468
R21 Y.n2 Y.n1 172.504
R22 Y.n3 Y.n0 130.205
R23 Y.n0 Y.t1 40
R24 Y.n0 Y.t2 40
R25 Y.n1 Y.t0 27.58
R26 Y.n1 Y.t4 27.58
R27 Y Y.n2 22.641
R28 Y.n3 Y 13.485
R29 Y Y.n3 2.057
R30 KAPWR.n0 KAPWR.t0 39.355
R31 KAPWR.n3 KAPWR.t1 24.625
R32 KAPWR.n1 KAPWR.t2 22.819
R33 KAPWR.n4 KAPWR.n3 9.3
R34 KAPWR.n2 KAPWR.n1 4.55
R35 KAPWR.n6 KAPWR.n5 4.293
R36 KAPWR.n3 KAPWR.n2 2.955
R37 KAPWR.n5 KAPWR.n4 2.461
R38 KAPWR KAPWR.n7 0.279
R39 KAPWR.n7 KAPWR.n6 0.036
R40 KAPWR.n6 KAPWR.n0 0.004
R41 VPB.t2 VPB.t0 254.517
R42 VPB.t1 VPB.t2 254.517
R43 VPB VPB.t1 207.165
C0 Y VGND 0.22fF
C1 Y KAPWR 0.43fF
C2 A Y 0.28fF
C3 KAPWR VPWR 0.79fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__lpflow_clkinvkapwr_4.ext - technology: sky130A

.subckt sky130_fd_sc_hd__lpflow_clkinvkapwr_4 A Y KAPWR VPWR VGND VNB VPB
X0 Y.t9 A.t0 KAPWR.t2 VPB.t5 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 VGND.t3 A.t1 Y.t3 VNB sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 VGND.t2 A.t2 Y.t2 VNB sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3 KAPWR.t1 A.t3 Y.t8 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 KAPWR.t0 A.t4 Y.t7 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 Y.t1 A.t5 VGND.t1 VNB sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 Y.t6 A.t6 KAPWR.t5 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 Y.t0 A.t7 VGND.t0 VNB sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 Y.t5 A.t8 KAPWR.t4 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 KAPWR.t3 A.t9 Y.t4 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
R0 A.n0 A.t4 276.167
R1 A.n6 A.t6 247.604
R2 A.n2 A.t0 221.719
R3 A.n5 A.t9 221.719
R4 A.n13 A.t8 221.719
R5 A.n7 A.t3 221.719
R6 A.n2 A.t1 186.373
R7 A.n5 A.t5 186.373
R8 A.n13 A.t2 186.373
R9 A.n7 A.t7 186.373
R10 A.n1 A.n0 76
R11 A.n4 A.n3 76
R12 A.n15 A.n14 76
R13 A.n12 A.n11 76
R14 A.n10 A.n8 76
R15 A.n12 A.n8 60.696
R16 A.n14 A.n13 54.448
R17 A.n7 A.n6 50.877
R18 A.n3 A.n2 38.381
R19 A.n14 A.n5 22.314
R20 A.n4 A.n1 19.342
R21 A.n10 A.n9 19.342
R22 A A.n15 17.351
R23 A.n11 A 15.644
R24 A.n11 A 10.524
R25 A.n8 A.n7 9.818
R26 A.n15 A 8.817
R27 A.n13 A.n12 6.248
R28 A.n1 A 4.835
R29 A A.n10 3.697
R30 A.n9 A 3.128
R31 A A.n4 1.991
R32 KAPWR.n0 KAPWR.t0 41.866
R33 KAPWR.n18 KAPWR.t5 36.936
R34 KAPWR.n3 KAPWR.t2 25.67
R35 KAPWR.n11 KAPWR.t1 25.61
R36 KAPWR.n9 KAPWR.t4 22.468
R37 KAPWR.n2 KAPWR.n1 14.775
R38 KAPWR.n1 KAPWR.t3 12.805
R39 KAPWR.n12 KAPWR.n11 9.3
R40 KAPWR.n4 KAPWR.n3 8.958
R41 KAPWR.n19 KAPWR.n18 6.654
R42 KAPWR.n10 KAPWR.n9 4.869
R43 KAPWR.n6 KAPWR.n5 4.293
R44 KAPWR.n14 KAPWR.n13 4.293
R45 KAPWR.n13 KAPWR.n12 2.461
R46 KAPWR.n5 KAPWR.n4 2.461
R47 KAPWR.n11 KAPWR.n10 1.97
R48 KAPWR.n3 KAPWR.n2 1.898
R49 KAPWR.n8 KAPWR.n7 0.509
R50 KAPWR.n16 KAPWR.n15 0.453
R51 KAPWR.n18 KAPWR.n17 0.082
R52 KAPWR.n6 KAPWR.n0 0.036
R53 KAPWR.n15 KAPWR.n14 0.036
R54 KAPWR.n20 KAPWR.n19 0.036
R55 KAPWR KAPWR.n20 0.019
R56 KAPWR.n7 KAPWR.n6 0.004
R57 KAPWR.n14 KAPWR.n8 0.004
R58 KAPWR.n19 KAPWR.n16 0.004
R59 Y.n9 Y.n2 169.147
R60 Y.n8 Y.n3 169.147
R61 Y.n7 Y.n4 169.147
R62 Y.n7 Y.n6 146.446
R63 Y.n1 Y.n0 110.821
R64 Y.n6 Y.n5 110.469
R65 Y.n9 Y.n8 64.752
R66 Y.n8 Y.n7 64.752
R67 Y.n10 Y.n1 51.952
R68 Y.n6 Y.n1 45.176
R69 Y.n0 Y.t3 40
R70 Y.n0 Y.t1 40
R71 Y.n5 Y.t2 40
R72 Y.n5 Y.t0 40
R73 Y Y.n9 33.254
R74 Y.n2 Y.t7 27.58
R75 Y.n2 Y.t9 27.58
R76 Y.n3 Y.t4 27.58
R77 Y.n3 Y.t5 27.58
R78 Y.n4 Y.t8 27.58
R79 Y.n4 Y.t6 27.58
R80 Y.n10 Y 12.586
R81 Y Y.n10 1.92
R82 VPB.t5 VPB.t3 254.517
R83 VPB.t0 VPB.t5 254.517
R84 VPB.t1 VPB.t0 254.517
R85 VPB.t4 VPB.t1 254.517
R86 VPB.t2 VPB.t4 254.517
R87 VPB VPB.t2 219.003
R88 VGND.n2 VGND.t3 152.681
R89 VGND.n5 VGND.t0 149.422
R90 VGND.n1 VGND.n0 111.7
R91 VGND.n0 VGND.t1 40
R92 VGND.n0 VGND.t2 40
R93 VGND.n4 VGND.n3 4.65
R94 VGND.n6 VGND.n5 4.01
R95 VGND.n2 VGND.n1 3.921
R96 VGND.n4 VGND.n2 0.23
R97 VGND.n6 VGND.n4 0.135
R98 VGND VGND.n6 0.125
C0 Y VPWR 0.12fF
C1 KAPWR Y 0.83fF
C2 A Y 1.20fF
C3 KAPWR VPWR 1.45fF
C4 Y VGND 0.52fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__lpflow_clkinvkapwr_8.ext - technology: sky130A

.subckt sky130_fd_sc_hd__lpflow_clkinvkapwr_8 Y A KAPWR VGND VPWR VNB VPB
X0 Y.t17 A.t0 VGND.t5 VNB sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1 KAPWR.t11 A.t1 Y.t9 VPB.t11 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 Y.t16 A.t2 VGND.t4 VNB sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3 Y.t15 A.t3 VGND.t3 VNB sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 Y.t8 A.t4 KAPWR.t10 VPB.t10 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 KAPWR.t9 A.t5 Y.t7 VPB.t9 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 KAPWR.t8 A.t6 Y.t6 VPB.t8 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 Y.t14 A.t7 VGND.t2 VNB sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 Y.t5 A.t8 KAPWR.t7 VPB.t7 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 VGND.t1 A.t9 Y.t13 VNB sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10 Y.t4 A.t10 KAPWR.t6 VPB.t6 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 KAPWR.t5 A.t11 Y.t3 VPB.t5 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 VGND.t0 A.t12 Y.t12 VNB sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13 KAPWR.t4 A.t13 Y.t2 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14 Y.t1 A.t14 KAPWR.t3 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 VGND.t7 A.t15 Y.t11 VNB sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16 KAPWR.t2 A.t16 Y.t0 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17 Y.t19 A.t17 KAPWR.t1 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X18 Y.t18 A.t18 KAPWR.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X19 VGND.t6 A.t19 Y.t10 VNB sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
R0 A.n5 A.t11 225.91
R1 A.n41 A.t18 205.372
R2 A.n6 A.t8 192.799
R3 A.n4 A.t13 192.799
R4 A.n13 A.t14 192.799
R5 A.n15 A.t16 192.799
R6 A.n22 A.t17 192.799
R7 A.n2 A.t1 192.799
R8 A.n29 A.t4 192.799
R9 A.n32 A.t6 192.799
R10 A.n0 A.t10 192.799
R11 A.n40 A.t5 192.799
R12 A.n33 A.t0 117.286
R13 A.n31 A.t15 117.286
R14 A.n28 A.t7 117.286
R15 A.n23 A.t12 117.286
R16 A.n3 A.t3 117.286
R17 A.n16 A.t9 117.286
R18 A.n12 A.t2 117.286
R19 A.n7 A.t19 117.286
R20 A.n9 A.n8 76
R21 A.n11 A.n10 76
R22 A.n18 A.n17 76
R23 A.n21 A.n20 76
R24 A.n25 A.n24 76
R25 A.n27 A.n26 76
R26 A.n35 A.n34 76
R27 A.n37 A.n36 76
R28 A.n39 A.n38 76
R29 A.n42 A.n41 76
R30 A.n38 A.n37 28.5
R31 A.n23 A.n22 24.309
R32 A.n41 A.n40 22.633
R33 A.n27 A.n2 21.375
R34 A.n7 A.n6 20.956
R35 A.n11 A.n4 19.699
R36 A.n34 A.n33 18.86
R37 A.n14 A.n3 17.184
R38 A.n20 A.n19 17.066
R39 A.n35 A.n1 17.066
R40 A.n42 A.n39 17.066
R41 A.n26 A 16.564
R42 A A.n18 15.56
R43 A.n30 A.n29 14.669
R44 A.n10 A 13.552
R45 A.n13 A.n12 13.412
R46 A.n17 A.n13 12.993
R47 A.n16 A.n15 12.573
R48 A.n25 A 12.549
R49 A.n36 A 11.545
R50 A.n36 A 11.545
R51 A.n21 A.n3 11.316
R52 A.n31 A.n30 11.316
R53 A A.n25 10.541
R54 A.n29 A.n28 10.059
R55 A.n17 A.n16 9.64
R56 A.n10 A 9.537
R57 A.n32 A.n31 9.22
R58 A.n8 A.n4 8.801
R59 A.n33 A.n0 8.382
R60 A.n34 A.n32 7.963
R61 A.n18 A 7.529
R62 A.n24 A.n2 7.125
R63 A.n26 A 6.525
R64 A.n15 A.n14 6.286
R65 A A.n35 5.521
R66 A.n39 A 5.521
R67 A.n8 A.n7 5.448
R68 A.n20 A 4.517
R69 A.n24 A.n23 3.772
R70 A.n28 A.n27 3.772
R71 A A.n9 3.513
R72 A.n6 A.n5 2.095
R73 A.n12 A.n11 2.095
R74 A.n19 A 1.505
R75 A.n37 A.n0 1.257
R76 A A.n1 0.501
R77 A A.n42 0.501
R78 A.n22 A.n21 0.419
R79 VGND.n3 VGND.t6 151.62
R80 VGND.n0 VGND.t5 147.627
R81 VGND.n2 VGND.n1 107.627
R82 VGND.n7 VGND.n6 107.627
R83 VGND.n12 VGND.n11 107.627
R84 VGND.n1 VGND.t4 40
R85 VGND.n1 VGND.t1 40
R86 VGND.n6 VGND.t3 40
R87 VGND.n6 VGND.t0 40
R88 VGND.n11 VGND.t2 40
R89 VGND.n11 VGND.t7 40
R90 VGND.n5 VGND.n4 4.65
R91 VGND.n8 VGND.n7 4.65
R92 VGND.n10 VGND.n9 4.65
R93 VGND.n13 VGND.n12 4.65
R94 VGND.n15 VGND.n14 4.65
R95 VGND.n16 VGND.n0 4.013
R96 VGND.n3 VGND.n2 3.923
R97 VGND.n5 VGND.n3 0.31
R98 VGND VGND.n16 0.241
R99 VGND.n16 VGND.n15 0.137
R100 VGND.n8 VGND.n5 0.119
R101 VGND.n10 VGND.n8 0.119
R102 VGND.n13 VGND.n10 0.119
R103 VGND.n15 VGND.n13 0.119
R104 Y.n14 Y.n13 181.458
R105 Y.n14 Y.n7 174.971
R106 Y.n19 Y.n2 169.147
R107 Y.n18 Y.n3 169.147
R108 Y.n17 Y.n4 169.147
R109 Y.n16 Y.n5 169.147
R110 Y.n15 Y.n6 169.147
R111 Y.n1 Y.n0 115.068
R112 Y.n9 Y.n8 115.068
R113 Y.n11 Y.n10 115.068
R114 Y.n13 Y.n12 115.068
R115 Y.n20 Y.n1 65.129
R116 Y.n15 Y.n14 63.623
R117 Y.n19 Y.n18 63.247
R118 Y.n18 Y.n17 63.247
R119 Y.n17 Y.n16 63.247
R120 Y.n16 Y.n15 63.247
R121 Y.n9 Y.n1 50.447
R122 Y.n11 Y.n9 50.447
R123 Y.n13 Y.n11 50.447
R124 Y.n0 Y.t10 40
R125 Y.n0 Y.t16 40
R126 Y.n8 Y.t13 40
R127 Y.n8 Y.t15 40
R128 Y.n10 Y.t12 40
R129 Y.n10 Y.t14 40
R130 Y.n12 Y.t11 40
R131 Y.n12 Y.t17 40
R132 Y.n2 Y.t3 26.595
R133 Y.n2 Y.t5 26.595
R134 Y.n3 Y.t2 26.595
R135 Y.n3 Y.t1 26.595
R136 Y.n4 Y.t0 26.595
R137 Y.n4 Y.t19 26.595
R138 Y.n5 Y.t9 26.595
R139 Y.n5 Y.t8 26.595
R140 Y.n6 Y.t6 26.595
R141 Y.n6 Y.t4 26.595
R142 Y.n7 Y.t7 26.595
R143 Y.n7 Y.t18 26.595
R144 Y Y.n19 26.198
R145 Y.n20 Y 15.407
R146 Y Y.n20 0.711
R147 KAPWR.n0 KAPWR.t5 40.083
R148 KAPWR.n42 KAPWR.t0 38.477
R149 KAPWR.n35 KAPWR.t9 24.625
R150 KAPWR.n27 KAPWR.t10 23.73
R151 KAPWR.n3 KAPWR.t4 23.64
R152 KAPWR.n9 KAPWR.t3 22.531
R153 KAPWR.n33 KAPWR.t6 21.834
R154 KAPWR.n1 KAPWR.t7 21.834
R155 KAPWR.n11 KAPWR.t2 21.67
R156 KAPWR.n19 KAPWR.t1 19.907
R157 KAPWR.n17 KAPWR.t11 16.745
R158 KAPWR.n26 KAPWR.n25 13.79
R159 KAPWR.n25 KAPWR.t8 12.805
R160 KAPWR.n18 KAPWR.n17 9.85
R161 KAPWR.n4 KAPWR.n3 9.3
R162 KAPWR.n12 KAPWR.n11 9.3
R163 KAPWR.n36 KAPWR.n35 9.3
R164 KAPWR.n28 KAPWR.n27 8.929
R165 KAPWR.n20 KAPWR.n19 8.816
R166 KAPWR.n43 KAPWR.n42 6.634
R167 KAPWR.n19 KAPWR.n18 6.536
R168 KAPWR.n11 KAPWR.n10 4.925
R169 KAPWR.n34 KAPWR.n33 4.55
R170 KAPWR.n2 KAPWR.n1 4.55
R171 KAPWR.n6 KAPWR.n5 4.293
R172 KAPWR.n14 KAPWR.n13 4.293
R173 KAPWR.n22 KAPWR.n21 4.293
R174 KAPWR.n30 KAPWR.n29 4.293
R175 KAPWR.n38 KAPWR.n37 4.293
R176 KAPWR.n10 KAPWR.n9 3.908
R177 KAPWR.n35 KAPWR.n34 2.955
R178 KAPWR.n3 KAPWR.n2 2.955
R179 KAPWR.n27 KAPWR.n26 2.838
R180 KAPWR.n37 KAPWR.n36 2.461
R181 KAPWR.n29 KAPWR.n28 2.461
R182 KAPWR.n21 KAPWR.n20 2.461
R183 KAPWR.n13 KAPWR.n12 2.461
R184 KAPWR.n5 KAPWR.n4 2.461
R185 KAPWR.n32 KAPWR.n31 0.505
R186 KAPWR.n24 KAPWR.n23 0.456
R187 KAPWR.n40 KAPWR.n39 0.452
R188 KAPWR.n8 KAPWR.n7 0.449
R189 KAPWR.n16 KAPWR.n15 0.354
R190 KAPWR.n42 KAPWR.n41 0.102
R191 KAPWR.n7 KAPWR.n6 0.036
R192 KAPWR.n30 KAPWR.n24 0.033
R193 KAPWR.n39 KAPWR.n38 0.033
R194 KAPWR.n15 KAPWR.n14 0.031
R195 KAPWR.n22 KAPWR.n16 0.024
R196 KAPWR KAPWR.n43 0.021
R197 KAPWR.n23 KAPWR.n22 0.016
R198 KAPWR.n14 KAPWR.n8 0.009
R199 KAPWR.n43 KAPWR.n40 0.009
R200 KAPWR.n31 KAPWR.n30 0.007
R201 KAPWR.n38 KAPWR.n32 0.007
R202 KAPWR.n6 KAPWR.n0 0.004
R203 VPB.t9 VPB.t6 251.557
R204 VPB.t7 VPB.t5 248.598
R205 VPB.t4 VPB.t7 248.598
R206 VPB.t3 VPB.t4 248.598
R207 VPB.t2 VPB.t3 248.598
R208 VPB.t1 VPB.t2 248.598
R209 VPB.t11 VPB.t1 248.598
R210 VPB.t10 VPB.t11 248.598
R211 VPB.t8 VPB.t10 248.598
R212 VPB.t6 VPB.t8 248.598
R213 VPB.t0 VPB.t9 248.598
R214 VPB VPB.t0 189.408
C0 KAPWR VGND 0.16fF
C1 VPWR KAPWR 2.71fF
C2 Y VGND 0.93fF
C3 VPWR Y 0.24fF
C4 A Y 2.37fF
C5 VPWR VPB 0.11fF
C6 VPB A 0.14fF
C7 KAPWR Y 1.55fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__lpflow_clkinvkapwr_16.ext - technology: sky130A

.subckt sky130_fd_sc_hd__lpflow_clkinvkapwr_16 Y A KAPWR VGND VPWR VNB VPB
X0 VGND.t15 A.t0 Y.t39 VNB sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1 Y.t20 A.t1 KAPWR.t23 VPB.t23 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 KAPWR.t22 A.t2 Y.t19 VPB.t22 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 Y.t18 A.t3 KAPWR.t21 VPB.t21 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 VGND.t14 A.t4 Y.t38 VNB sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 KAPWR.t20 A.t5 Y.t17 VPB.t20 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 Y.t37 A.t6 VGND.t13 VNB sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7 VGND.t12 A.t7 Y.t36 VNB sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 KAPWR.t19 A.t8 Y.t16 VPB.t19 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 KAPWR.t18 A.t9 Y.t15 VPB.t18 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 Y.t35 A.t10 VGND.t11 VNB sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11 Y.t14 A.t11 KAPWR.t17 VPB.t17 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 KAPWR.t16 A.t12 Y.t13 VPB.t16 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13 VGND.t10 A.t13 Y.t34 VNB sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14 Y.t12 A.t14 KAPWR.t15 VPB.t15 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 KAPWR.t14 A.t15 Y.t11 VPB.t14 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16 Y.t10 A.t16 KAPWR.t13 VPB.t13 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17 Y.t9 A.t17 KAPWR.t12 VPB.t12 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X18 Y.t33 A.t18 VGND.t9 VNB sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19 VGND.t8 A.t19 Y.t8 VNB sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20 Y.t7 A.t20 VGND.t7 VNB sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21 VGND.t6 A.t21 Y.t6 VNB sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22 Y.t32 A.t22 KAPWR.t11 VPB.t11 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X23 KAPWR.t10 A.t23 Y.t31 VPB.t10 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X24 Y.t30 A.t24 KAPWR.t9 VPB.t9 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X25 Y.t29 A.t25 KAPWR.t8 VPB.t8 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X26 KAPWR.t7 A.t26 Y.t28 VPB.t7 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X27 Y.t5 A.t27 VGND.t5 VNB sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X28 Y.t27 A.t28 KAPWR.t6 VPB.t6 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X29 KAPWR.t5 A.t29 Y.t26 VPB.t5 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X30 KAPWR.t4 A.t30 Y.t25 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X31 Y.t4 A.t31 VGND.t4 VNB sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X32 VGND.t3 A.t32 Y.t3 VNB sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X33 KAPWR.t3 A.t33 Y.t24 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X34 Y.t2 A.t34 VGND.t2 VNB sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X35 Y.t23 A.t35 KAPWR.t2 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X36 Y.t1 A.t36 VGND.t1 VNB sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X37 KAPWR.t1 A.t37 Y.t22 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X38 Y.t21 A.t38 KAPWR.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X39 VGND.t0 A.t39 Y.t0 VNB sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
R0 A.n3 A.t30 218.104
R1 A.n33 A.t14 218.104
R2 A.n4 A.t28 204.046
R3 A.n6 A.t29 204.046
R4 A.n26 A.t17 204.046
R5 A.n24 A.t5 204.046
R6 A.n23 A.t38 204.046
R7 A.n22 A.t26 204.046
R8 A.n21 A.t16 204.046
R9 A.n20 A.t15 204.046
R10 A.n19 A.t3 204.046
R11 A.n18 A.t37 204.046
R12 A.n17 A.t25 204.046
R13 A.n44 A.t12 204.046
R14 A.n45 A.t24 204.046
R15 A.n46 A.t2 204.046
R16 A.n47 A.t35 204.046
R17 A.n48 A.t23 204.046
R18 A.n49 A.t11 204.046
R19 A.n50 A.t9 204.046
R20 A.n51 A.t1 204.046
R21 A.n38 A.t33 204.046
R22 A.n40 A.t22 204.046
R23 A.n34 A.t8 204.046
R24 A.n24 A.t0 175.126
R25 A.n23 A.t10 175.126
R26 A.n22 A.t4 175.126
R27 A.n21 A.t18 175.126
R28 A.n20 A.t7 175.126
R29 A.n19 A.t20 175.126
R30 A.n18 A.t32 175.126
R31 A.n17 A.t27 175.126
R32 A.n44 A.t39 175.126
R33 A.n45 A.t34 175.126
R34 A.n46 A.t13 175.126
R35 A.n47 A.t6 175.126
R36 A.n48 A.t19 175.126
R37 A.n49 A.t31 175.126
R38 A.n50 A.t21 175.126
R39 A.n51 A.t36 175.126
R40 A.n36 A.n33 87.452
R41 A.n45 A.n44 78.325
R42 A.n36 A.n35 76
R43 A.n46 A.n45 62.258
R44 A.n24 A.n23 57.572
R45 A.n23 A.n22 57.572
R46 A.n22 A.n21 57.572
R47 A.n21 A.n20 57.572
R48 A.n20 A.n19 57.572
R49 A.n19 A.n18 57.572
R50 A.n18 A.n17 57.572
R51 A.n47 A.n46 57.572
R52 A.n48 A.n47 57.572
R53 A.n49 A.n48 57.572
R54 A.n50 A.n49 57.572
R55 A.n51 A.n50 57.572
R56 A.n4 A.n3 43.513
R57 A.n9 A.n5 38.158
R58 A.n41 A.n40 35.48
R59 A.n25 A.n24 34.141
R60 A.n54 A.n51 26.108
R61 A.n26 A.n25 23.43
R62 A.n41 A.n38 22.091
R63 A.n27 A.n26 21.422
R64 A.n42 A.n37 11.452
R65 A.n37 A.n36 11.452
R66 A.n16 A.n15 10.711
R67 A.n40 A.n39 10.041
R68 A.n10 A.n9 9.3
R69 A.n28 A.n27 9.3
R70 A.n55 A.n54 9.3
R71 A.n42 A.n41 8.286
R72 A.n54 A.n53 8.033
R73 A.n11 A.n0 7.806
R74 A.n9 A.n8 7.363
R75 A.n43 A.n32 6.435
R76 A.n7 A.n6 6.025
R77 A.n31 A.n30 4.65
R78 A.n8 A.n7 4.016
R79 A.n53 A.n52 3.347
R80 A.n43 A.n42 3.341
R81 A.n55 A.n43 3.33
R82 A.n14 A.n13 2.694
R83 A.n30 A.n29 2.694
R84 A.n12 A.n11 2.106
R85 A.n5 A.n4 2.008
R86 A.n35 A.n34 2.008
R87 A.n10 A.n2 1.852
R88 A.n11 A.n10 1.401
R89 A A.n57 1.178
R90 A.n2 A.n1 1.01
R91 A A.n55 0.842
R92 A.n57 A.n56 0.842
R93 A.n27 A.n16 0.669
R94 A.n28 A.n14 0.168
R95 A.n30 A.n28 0.168
R96 A.n32 A.n31 0.043
R97 A.n31 A.n12 0.002
R98 Y.n20 Y.n18 209.477
R99 Y.n6 Y.n5 161.753
R100 Y.n11 Y.n9 161.556
R101 Y.n31 Y.n29 160.336
R102 Y.n20 Y.n19 157.058
R103 Y.n6 Y.n4 157.058
R104 Y.n7 Y.n3 157.058
R105 Y.n13 Y.n0 157.058
R106 Y.n22 Y.n21 157.058
R107 Y.n24 Y.n23 157.058
R108 Y.n26 Y.n25 157.058
R109 Y.n28 Y.n27 157.058
R110 Y.n8 Y.n2 147.682
R111 Y.n11 Y.n10 147.464
R112 Y.n12 Y.n1 144.233
R113 Y.n28 Y.n14 142.164
R114 Y.n26 Y.n15 142.164
R115 Y.n24 Y.n16 142.164
R116 Y.n22 Y.n17 142.164
R117 Y Y.n30 129.071
R118 Y.n30 Y.t0 75.714
R119 Y.n29 Y.t30 53.19
R120 Y.n7 Y.n6 51.492
R121 Y.n22 Y.n20 51.2
R122 Y.n30 Y.t2 48.571
R123 Y.n24 Y.n22 44.032
R124 Y.n26 Y.n24 44.032
R125 Y.n28 Y.n26 44.032
R126 Y.n31 Y.n28 40.704
R127 Y.n14 Y.t3 40
R128 Y.n14 Y.t5 40
R129 Y.n15 Y.t36 40
R130 Y.n15 Y.t7 40
R131 Y.n16 Y.t38 40
R132 Y.n16 Y.t33 40
R133 Y.n17 Y.t39 40
R134 Y.n17 Y.t35 40
R135 Y.n2 Y.t6 40
R136 Y.n2 Y.t1 40
R137 Y.n10 Y.t8 40
R138 Y.n10 Y.t4 40
R139 Y.n1 Y.t34 40
R140 Y.n1 Y.t37 40
R141 Y.n31 Y.n13 39.168
R142 Y.n12 Y.n11 37.12
R143 Y.n11 Y.n8 36.864
R144 Y.n29 Y.t13 32.505
R145 Y.n27 Y.t22 27.58
R146 Y.n27 Y.t29 27.58
R147 Y.n25 Y.t11 27.58
R148 Y.n25 Y.t18 27.58
R149 Y.n23 Y.t28 27.58
R150 Y.n23 Y.t10 27.58
R151 Y.n21 Y.t17 27.58
R152 Y.n21 Y.t21 27.58
R153 Y.n19 Y.t26 27.58
R154 Y.n19 Y.t9 27.58
R155 Y.n18 Y.t25 27.58
R156 Y.n18 Y.t27 27.58
R157 Y.n0 Y.t19 27.58
R158 Y.n0 Y.t23 27.58
R159 Y.n3 Y.t15 27.58
R160 Y.n3 Y.t20 27.58
R161 Y.n5 Y.t16 27.58
R162 Y.n5 Y.t12 27.58
R163 Y.n4 Y.t24 27.58
R164 Y.n4 Y.t32 27.58
R165 Y.n9 Y.t31 27.58
R166 Y.n9 Y.t14 27.58
R167 Y.n31 Y 3.474
R168 Y Y.n31 2.56
R169 Y.n8 Y.n7 0.768
R170 Y.n13 Y.n12 0.256
R171 VGND.n1 VGND.t15 157.105
R172 VGND.n0 VGND.t1 153.596
R173 VGND.n13 VGND.n12 117.815
R174 VGND.n3 VGND.n2 113.994
R175 VGND.n9 VGND.n8 113.994
R176 VGND.n19 VGND.n18 113.994
R177 VGND.n26 VGND.n25 113.994
R178 VGND.n30 VGND.n29 113.994
R179 VGND.n36 VGND.n35 113.994
R180 VGND.n25 VGND.t10 47.142
R181 VGND.n25 VGND.t2 42.857
R182 VGND.n2 VGND.t11 40
R183 VGND.n2 VGND.t14 40
R184 VGND.n8 VGND.t9 40
R185 VGND.n8 VGND.t12 40
R186 VGND.n12 VGND.t7 40
R187 VGND.n12 VGND.t3 40
R188 VGND.n18 VGND.t5 40
R189 VGND.n18 VGND.t0 40
R190 VGND.n29 VGND.t13 40
R191 VGND.n29 VGND.t8 40
R192 VGND.n35 VGND.t4 40
R193 VGND.n35 VGND.t6 40
R194 VGND.n14 VGND.n13 7.152
R195 VGND.n27 VGND.n26 7.152
R196 VGND.n10 VGND.n9 6.023
R197 VGND.n31 VGND.n30 4.894
R198 VGND.n5 VGND.n4 4.65
R199 VGND.n7 VGND.n6 4.65
R200 VGND.n11 VGND.n10 4.65
R201 VGND.n15 VGND.n14 4.65
R202 VGND.n17 VGND.n16 4.65
R203 VGND.n20 VGND.n19 4.65
R204 VGND.n22 VGND.n21 4.65
R205 VGND.n24 VGND.n23 4.65
R206 VGND.n28 VGND.n27 4.65
R207 VGND.n32 VGND.n31 4.65
R208 VGND.n34 VGND.n33 4.65
R209 VGND.n38 VGND.n37 4.65
R210 VGND.n40 VGND.n39 4.65
R211 VGND.n41 VGND.n0 3.838
R212 VGND.n4 VGND.n3 1.505
R213 VGND.n5 VGND.n1 0.577
R214 VGND VGND.n41 0.477
R215 VGND.n37 VGND.n36 0.376
R216 VGND.n41 VGND.n40 0.142
R217 VGND.n7 VGND.n5 0.119
R218 VGND.n11 VGND.n7 0.119
R219 VGND.n15 VGND.n11 0.119
R220 VGND.n17 VGND.n15 0.119
R221 VGND.n20 VGND.n17 0.119
R222 VGND.n22 VGND.n20 0.119
R223 VGND.n24 VGND.n22 0.119
R224 VGND.n28 VGND.n24 0.119
R225 VGND.n32 VGND.n28 0.119
R226 VGND.n34 VGND.n32 0.119
R227 VGND.n38 VGND.n34 0.119
R228 VGND.n40 VGND.n38 0.119
R229 KAPWR.n0 KAPWR.t4 40.173
R230 KAPWR.n89 KAPWR.t15 38.68
R231 KAPWR.n65 KAPWR.t17 27.58
R232 KAPWR.n66 KAPWR.t18 26.875
R233 KAPWR.n51 KAPWR.t9 26.714
R234 KAPWR.n19 KAPWR.t0 26.626
R235 KAPWR.n74 KAPWR.t3 25.61
R236 KAPWR.n11 KAPWR.t20 25.61
R237 KAPWR.n3 KAPWR.t5 25.61
R238 KAPWR.n41 KAPWR.t8 25.534
R239 KAPWR.n35 KAPWR.t1 24.625
R240 KAPWR.n27 KAPWR.t14 24.625
R241 KAPWR.n80 KAPWR.t11 23.859
R242 KAPWR.n33 KAPWR.t21 22.814
R243 KAPWR.n25 KAPWR.t13 22.814
R244 KAPWR.n72 KAPWR.t23 22.463
R245 KAPWR.n9 KAPWR.t12 22.463
R246 KAPWR.n1 KAPWR.t6 22.463
R247 KAPWR.n59 KAPWR.t2 21.848
R248 KAPWR.n82 KAPWR.t19 21.67
R249 KAPWR.n49 KAPWR.t22 18.715
R250 KAPWR.n43 KAPWR.t16 18.715
R251 KAPWR.n57 KAPWR.t10 16.745
R252 KAPWR.n18 KAPWR.n17 15.76
R253 KAPWR.n50 KAPWR.n49 12.805
R254 KAPWR.n17 KAPWR.t7 11.82
R255 KAPWR.n58 KAPWR.n57 10.835
R256 KAPWR.n4 KAPWR.n3 9.3
R257 KAPWR.n12 KAPWR.n11 9.3
R258 KAPWR.n28 KAPWR.n27 9.3
R259 KAPWR.n36 KAPWR.n35 9.3
R260 KAPWR.n44 KAPWR.n43 9.3
R261 KAPWR.n75 KAPWR.n74 9.3
R262 KAPWR.n83 KAPWR.n82 9.3
R263 KAPWR.n20 KAPWR.n19 8.987
R264 KAPWR.n52 KAPWR.n51 8.901
R265 KAPWR.n60 KAPWR.n59 8.845
R266 KAPWR.n67 KAPWR.n66 8.637
R267 KAPWR.n43 KAPWR.n42 7.88
R268 KAPWR.n90 KAPWR.n89 7.08
R269 KAPWR.n82 KAPWR.n81 5.91
R270 KAPWR.n59 KAPWR.n58 5.621
R271 KAPWR.n73 KAPWR.n72 4.874
R272 KAPWR.n10 KAPWR.n9 4.874
R273 KAPWR.n2 KAPWR.n1 4.874
R274 KAPWR.n34 KAPWR.n33 4.554
R275 KAPWR.n26 KAPWR.n25 4.554
R276 KAPWR.n6 KAPWR.n5 4.465
R277 KAPWR.n14 KAPWR.n13 4.465
R278 KAPWR.n22 KAPWR.n21 4.465
R279 KAPWR.n30 KAPWR.n29 4.465
R280 KAPWR.n38 KAPWR.n37 4.465
R281 KAPWR.n46 KAPWR.n45 4.465
R282 KAPWR.n54 KAPWR.n53 4.465
R283 KAPWR.n62 KAPWR.n61 4.465
R284 KAPWR.n69 KAPWR.n68 4.465
R285 KAPWR.n77 KAPWR.n76 4.465
R286 KAPWR.n85 KAPWR.n84 4.465
R287 KAPWR.n51 KAPWR.n50 3.771
R288 KAPWR.n81 KAPWR.n80 3.59
R289 KAPWR.n35 KAPWR.n34 2.955
R290 KAPWR.n27 KAPWR.n26 2.955
R291 KAPWR.n42 KAPWR.n41 2.944
R292 KAPWR.n84 KAPWR.n83 2.894
R293 KAPWR.n76 KAPWR.n75 2.894
R294 KAPWR.n68 KAPWR.n67 2.894
R295 KAPWR.n61 KAPWR.n60 2.894
R296 KAPWR.n53 KAPWR.n52 2.894
R297 KAPWR.n45 KAPWR.n44 2.894
R298 KAPWR.n37 KAPWR.n36 2.894
R299 KAPWR.n29 KAPWR.n28 2.894
R300 KAPWR.n21 KAPWR.n20 2.894
R301 KAPWR.n13 KAPWR.n12 2.894
R302 KAPWR.n5 KAPWR.n4 2.894
R303 KAPWR.n74 KAPWR.n73 1.97
R304 KAPWR.n11 KAPWR.n10 1.97
R305 KAPWR.n3 KAPWR.n2 1.97
R306 KAPWR.n19 KAPWR.n18 0.952
R307 KAPWR.n24 KAPWR.n23 0.509
R308 KAPWR.n71 KAPWR.n70 0.502
R309 KAPWR.n40 KAPWR.n39 0.476
R310 KAPWR.n64 KAPWR.n63 0.476
R311 KAPWR.n48 KAPWR.n47 0.469
R312 KAPWR.n79 KAPWR.n78 0.469
R313 KAPWR.n56 KAPWR.n55 0.458
R314 KAPWR.n8 KAPWR.n7 0.454
R315 KAPWR.n32 KAPWR.n31 0.453
R316 KAPWR.n87 KAPWR.n86 0.451
R317 KAPWR.n16 KAPWR.n15 0.401
R318 KAPWR.n66 KAPWR.n65 0.248
R319 KAPWR.n89 KAPWR.n88 0.231
R320 KAPWR.n7 KAPWR.n6 0.038
R321 KAPWR.n15 KAPWR.n14 0.038
R322 KAPWR.n69 KAPWR.n64 0.038
R323 KAPWR.n78 KAPWR.n77 0.038
R324 KAPWR.n22 KAPWR.n16 0.036
R325 KAPWR.n31 KAPWR.n30 0.036
R326 KAPWR.n39 KAPWR.n38 0.036
R327 KAPWR.n54 KAPWR.n48 0.028
R328 KAPWR.n86 KAPWR.n85 0.028
R329 KAPWR.n91 KAPWR.n90 0.026
R330 KAPWR.n62 KAPWR.n56 0.024
R331 KAPWR.n47 KAPWR.n46 0.021
R332 KAPWR.n46 KAPWR.n40 0.019
R333 KAPWR.n63 KAPWR.n62 0.016
R334 KAPWR.n90 KAPWR.n87 0.014
R335 KAPWR.n55 KAPWR.n54 0.012
R336 KAPWR.n85 KAPWR.n79 0.012
R337 KAPWR.n23 KAPWR.n22 0.004
R338 KAPWR.n30 KAPWR.n24 0.004
R339 KAPWR.n38 KAPWR.n32 0.004
R340 KAPWR.n6 KAPWR.n0 0.002
R341 KAPWR.n14 KAPWR.n8 0.002
R342 KAPWR.n70 KAPWR.n69 0.002
R343 KAPWR.n77 KAPWR.n71 0.002
R344 KAPWR KAPWR.n91 0.002
R345 VPB.t9 VPB.t16 346.261
R346 VPB.t22 VPB.t9 275.233
R347 VPB.t6 VPB.t4 254.517
R348 VPB.t5 VPB.t6 254.517
R349 VPB.t12 VPB.t5 254.517
R350 VPB.t20 VPB.t12 254.517
R351 VPB.t0 VPB.t20 254.517
R352 VPB.t7 VPB.t0 254.517
R353 VPB.t13 VPB.t7 254.517
R354 VPB.t14 VPB.t13 254.517
R355 VPB.t21 VPB.t14 254.517
R356 VPB.t1 VPB.t21 254.517
R357 VPB.t8 VPB.t1 254.517
R358 VPB.t16 VPB.t8 254.517
R359 VPB.t2 VPB.t22 254.517
R360 VPB.t10 VPB.t2 254.517
R361 VPB.t17 VPB.t10 254.517
R362 VPB.t18 VPB.t17 254.517
R363 VPB.t23 VPB.t18 254.517
R364 VPB.t3 VPB.t23 254.517
R365 VPB.t11 VPB.t3 254.517
R366 VPB.t19 VPB.t11 254.517
R367 VPB.t15 VPB.t19 254.517
R368 VPB VPB.t15 201.246
C0 A VPWR 0.14fF
C1 KAPWR VGND 0.11fF
C2 A KAPWR 0.58fF
C3 KAPWR VPWR 5.05fF
C4 Y VGND 1.37fF
C5 A Y 0.94fF
C6 VPB A 0.32fF
C7 Y VPWR 0.56fF
C8 A VGND 0.71fF
C9 VPB VPWR 0.20fF
C10 KAPWR Y 2.85fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__lpflow_decapkapwr_3.ext - technology: sky130A

.subckt sky130_fd_sc_hd__lpflow_decapkapwr_3 VPWR VGND KAPWR VNB VPB
X0 KAPWR.t1 VGND.t2 KAPWR.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=870000u l=590000u
X1 VGND.t1 KAPWR.t2 VGND.t0 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=550000u l=590000u
R0 VGND.n1 VGND.t2 183.08
R1 VGND.n0 VGND.t0 123.916
R2 VGND.n2 VGND.t1 121.954
R3 VGND.n3 VGND.n2 5.067
R4 VGND.n3 VGND.n0 1.644
R5 VGND.n2 VGND.n1 1.182
R6 VGND VGND.n3 0.022
R7 KAPWR.n4 KAPWR.t0 170.48
R8 KAPWR.n2 KAPWR.t1 170.48
R9 KAPWR.n5 KAPWR.t2 166.281
R10 KAPWR.n3 KAPWR.n2 9.051
R11 KAPWR.n8 KAPWR.n4 9.051
R12 KAPWR.n10 KAPWR.n9 4.65
R13 KAPWR.n10 KAPWR.n8 2.72
R14 KAPWR.n11 KAPWR.n3 2.495
R15 KAPWR.n7 KAPWR.n6 0.973
R16 KAPWR.n1 KAPWR.n0 0.973
R17 KAPWR.n11 KAPWR.n10 0.226
R18 KAPWR.n6 KAPWR.n5 0.208
R19 KAPWR.n8 KAPWR.n7 0.203
R20 KAPWR.n3 KAPWR.n1 0.203
R21 KAPWR KAPWR.n11 0.027
R22 VPB VPB.t0 315.767
R23 VNB VNB.t0 7416.41
C0 KAPWR VPWR 0.70fF
C1 VGND KAPWR 0.44fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__lpflow_decapkapwr_4.ext - technology: sky130A

.subckt sky130_fd_sc_hd__lpflow_decapkapwr_4 VGND VPWR KAPWR VNB VPB
X0 KAPWR.t1 VGND.t2 KAPWR.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X1 VGND.t1 KAPWR.t2 VGND.t0 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
R0 VGND.n0 VGND.t2 142.306
R1 VGND.n1 VGND.t0 124.813
R2 VGND.n2 VGND.t1 121.954
R3 VGND.n1 VGND.n0 5.732
R4 VGND.n3 VGND.n2 5.058
R5 VGND.n3 VGND.n1 0.657
R6 VGND VGND.n3 0.022
R7 KAPWR.n4 KAPWR.t0 170.48
R8 KAPWR.n2 KAPWR.t1 170.48
R9 KAPWR.n5 KAPWR.t2 134.961
R10 KAPWR.n3 KAPWR.n2 9.051
R11 KAPWR.n8 KAPWR.n4 9.051
R12 KAPWR.n10 KAPWR.n9 4.65
R13 KAPWR.n12 KAPWR.n11 4.65
R14 KAPWR.n10 KAPWR.n8 2.72
R15 KAPWR.n13 KAPWR.n3 2.495
R16 KAPWR.n6 KAPWR.n5 1.808
R17 KAPWR.n7 KAPWR.n6 0.973
R18 KAPWR.n1 KAPWR.n0 0.973
R19 KAPWR.n13 KAPWR.n12 0.226
R20 KAPWR.n12 KAPWR.n10 0.221
R21 KAPWR.n8 KAPWR.n7 0.203
R22 KAPWR.n3 KAPWR.n1 0.203
R23 KAPWR KAPWR.n13 0.027
R24 VPB VPB.t0 458.722
R25 VNB VNB.t0 8665.79
C0 KAPWR VPWR 0.97fF
C1 VGND KAPWR 0.66fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__lpflow_decapkapwr_6.ext - technology: sky130A

.subckt sky130_fd_sc_hd__lpflow_decapkapwr_6 VPWR VGND KAPWR VNB VPB
X0 KAPWR.t1 VGND.t2 KAPWR.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.97e+06u
X1 VGND.t1 KAPWR.t2 VGND.t0 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=550000u l=1.97e+06u
R0 VGND.n1 VGND.t0 125.217
R1 VGND.n0 VGND.t1 121.954
R2 VGND.n0 VGND.t2 83.894
R3 VGND.n1 VGND.n0 3.853
R4 VGND VGND.n1 0.465
R5 KAPWR.n5 KAPWR.t0 179.4
R6 KAPWR.n2 KAPWR.t1 170.48
R7 KAPWR.n6 KAPWR.t2 95.458
R8 KAPWR.n3 KAPWR.n2 9.051
R9 KAPWR.n12 KAPWR.n11 4.65
R10 KAPWR.n14 KAPWR.n13 4.65
R11 KAPWR.n15 KAPWR.n3 2.495
R12 KAPWR.n10 KAPWR.n9 2.272
R13 KAPWR.n8 KAPWR.n7 2.062
R14 KAPWR.n7 KAPWR.n6 1.851
R15 KAPWR.n1 KAPWR.n0 0.973
R16 KAPWR.n9 KAPWR.n5 0.687
R17 KAPWR.n12 KAPWR.n10 0.33
R18 KAPWR.n10 KAPWR.n4 0.326
R19 KAPWR.n15 KAPWR.n14 0.226
R20 KAPWR.n14 KAPWR.n12 0.221
R21 KAPWR.n3 KAPWR.n1 0.203
R22 KAPWR.n9 KAPWR.n8 0.105
R23 KAPWR KAPWR.n15 0.027
R24 VPB VPB.t0 730.996
R25 VNB VNB.t0 11164.6
C0 KAPWR VPWR 1.49fF
C1 VGND KAPWR 1.10fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__lpflow_decapkapwr_8.ext - technology: sky130A

.subckt sky130_fd_sc_hd__lpflow_decapkapwr_8 VPWR VGND KAPWR VNB VPB
X0 KAPWR.t1 VGND.t2 KAPWR.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=870000u l=2.89e+06u
X1 VGND.t1 KAPWR.t2 VGND.t0 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=550000u l=2.89e+06u
R0 VGND.n1 VGND.t0 125.437
R1 VGND.n10 VGND.t1 121.954
R2 VGND.n4 VGND.n3 76
R3 VGND.n2 VGND.t2 34.296
R4 VGND.n11 VGND.n10 4.913
R5 VGND.n3 VGND.n2 4.857
R6 VGND.n6 VGND.n5 4.65
R7 VGND.n9 VGND.n8 4.65
R8 VGND.n1 VGND.n0 3.466
R9 VGND.n8 VGND.n7 1.139
R10 VGND.n5 VGND.n4 0.832
R11 VGND.n6 VGND.n1 0.235
R12 VGND.n9 VGND.n6 0.119
R13 VGND.n11 VGND.n9 0.119
R14 VGND VGND.n11 0.022
R15 KAPWR.n2 KAPWR.t1 170.48
R16 KAPWR.n4 KAPWR.t0 170.48
R17 KAPWR.n13 KAPWR.n12 76
R18 KAPWR.n11 KAPWR.t2 50.505
R19 KAPWR.n8 KAPWR.n4 9.053
R20 KAPWR.n3 KAPWR.n2 9.051
R21 KAPWR.n12 KAPWR.n11 7.118
R22 KAPWR.n10 KAPWR.n9 4.65
R23 KAPWR.n15 KAPWR.n14 4.65
R24 KAPWR.n18 KAPWR.n17 4.65
R25 KAPWR.n20 KAPWR.n19 4.65
R26 KAPWR.n22 KAPWR.n21 4.65
R27 KAPWR.n24 KAPWR.n23 4.65
R28 KAPWR.n10 KAPWR.n8 2.659
R29 KAPWR.n25 KAPWR.n3 2.495
R30 KAPWR.n6 KAPWR.n5 2.044
R31 KAPWR.n1 KAPWR.n0 0.973
R32 KAPWR.n14 KAPWR.n13 0.666
R33 KAPWR.n7 KAPWR.n6 0.622
R34 KAPWR.n25 KAPWR.n24 0.226
R35 KAPWR.n15 KAPWR.n10 0.221
R36 KAPWR.n18 KAPWR.n15 0.221
R37 KAPWR.n20 KAPWR.n18 0.221
R38 KAPWR.n22 KAPWR.n20 0.221
R39 KAPWR.n24 KAPWR.n22 0.221
R40 KAPWR.n3 KAPWR.n1 0.203
R41 KAPWR.n17 KAPWR.n16 0.177
R42 KAPWR.n8 KAPWR.n7 0.13
R43 KAPWR KAPWR.n25 0.027
R44 VPB VPB.t0 1003.27
R45 VNB VNB.t0 13663.3
C0 KAPWR VPWR 2.02fF
C1 KAPWR VGND 1.55fF
C2 VPB VGND 0.12fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__lpflow_decapkapwr_12.ext - technology: sky130A

.subckt sky130_fd_sc_hd__lpflow_decapkapwr_12 VGND VPWR KAPWR VNB VPB
X0 KAPWR.t1 VGND.t2 KAPWR.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=870000u l=4.73e+06u
X1 VGND.t1 KAPWR.t2 VGND.t0 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=550000u l=4.73e+06u
R0 VGND.n2 VGND.t0 125.719
R1 VGND.n17 VGND.t1 121.954
R2 VGND.n1 VGND.n0 76
R3 VGND.n6 VGND.n5 76
R4 VGND.n11 VGND.n10 76
R5 VGND.n9 VGND.t2 68.698
R6 VGND.n10 VGND.n9 31.477
R7 VGND.n18 VGND.n17 4.913
R8 VGND.n4 VGND.n3 4.65
R9 VGND.n8 VGND.n7 4.65
R10 VGND.n13 VGND.n12 4.65
R11 VGND.n16 VGND.n15 4.65
R12 VGND.n2 VGND.n1 3.42
R13 VGND.n7 VGND.n6 2.016
R14 VGND.n15 VGND.n14 1.139
R15 VGND.n12 VGND.n11 0.438
R16 VGND.n4 VGND.n2 0.187
R17 VGND.n8 VGND.n4 0.119
R18 VGND.n13 VGND.n8 0.119
R19 VGND.n16 VGND.n13 0.119
R20 VGND.n18 VGND.n16 0.119
R21 VGND VGND.n18 0.022
R22 KAPWR.n2 KAPWR.t1 170.48
R23 KAPWR.n4 KAPWR.t0 170.48
R24 KAPWR.n11 KAPWR.t2 107.792
R25 KAPWR.n23 KAPWR.n22 76
R26 KAPWR.n13 KAPWR.n12 76
R27 KAPWR.n19 KAPWR.n18 76
R28 KAPWR.n12 KAPWR.n11 30.493
R29 KAPWR.n7 KAPWR.n4 9.053
R30 KAPWR.n3 KAPWR.n2 9.051
R31 KAPWR.n10 KAPWR.n9 4.65
R32 KAPWR.n15 KAPWR.n14 4.65
R33 KAPWR.n17 KAPWR.n16 4.65
R34 KAPWR.n21 KAPWR.n20 4.65
R35 KAPWR.n25 KAPWR.n24 4.65
R36 KAPWR.n27 KAPWR.n26 4.65
R37 KAPWR.n29 KAPWR.n28 4.65
R38 KAPWR.n31 KAPWR.n30 4.65
R39 KAPWR.n33 KAPWR.n32 4.65
R40 KAPWR.n35 KAPWR.n34 4.65
R41 KAPWR.n10 KAPWR.n7 2.659
R42 KAPWR.n36 KAPWR.n3 2.495
R43 KAPWR.n20 KAPWR.n19 1.866
R44 KAPWR.n9 KAPWR.n8 0.977
R45 KAPWR.n1 KAPWR.n0 0.973
R46 KAPWR.n6 KAPWR.n5 0.622
R47 KAPWR.n14 KAPWR.n13 0.622
R48 KAPWR.n24 KAPWR.n23 0.266
R49 KAPWR.n36 KAPWR.n35 0.226
R50 KAPWR.n15 KAPWR.n10 0.221
R51 KAPWR.n17 KAPWR.n15 0.221
R52 KAPWR.n21 KAPWR.n17 0.221
R53 KAPWR.n25 KAPWR.n21 0.221
R54 KAPWR.n27 KAPWR.n25 0.221
R55 KAPWR.n29 KAPWR.n27 0.221
R56 KAPWR.n31 KAPWR.n29 0.221
R57 KAPWR.n33 KAPWR.n31 0.221
R58 KAPWR.n35 KAPWR.n33 0.221
R59 KAPWR.n3 KAPWR.n1 0.203
R60 KAPWR.n7 KAPWR.n6 0.13
R61 KAPWR KAPWR.n36 0.027
R62 VPB VPB.t0 1547.82
R63 VNB VNB.t0 -7851.29
C0 KAPWR VPWR 3.07fF
C1 VGND VPWR 0.11fF
C2 VGND KAPWR 2.43fF
C3 VPB KAPWR 0.13fF
C4 VPB VGND 0.18fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__lpflow_inputiso0n_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__lpflow_inputiso0n_1 VPWR VGND X SLEEP_B A VNB VPB
X0 VPWR.t0 SLEEP_B.t0 a_59_75.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1 X.t0 a_59_75.t3 VPWR.t1 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 VGND.t0 SLEEP_B.t1 a_145_75.t0 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3 a_59_75.t1 A.t0 VPWR.t2 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 X.t1 a_59_75.t4 VGND.t1 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 a_145_75.t1 A.t1 a_59_75.t2 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
R0 SLEEP_B.n0 SLEEP_B.t0 261.886
R1 SLEEP_B.n0 SLEEP_B.t1 155.846
R2 SLEEP_B SLEEP_B.n0 80.864
R3 a_59_75.n2 a_59_75.n1 380.446
R4 a_59_75.n0 a_59_75.t3 236.179
R5 a_59_75.n1 a_59_75.t2 222.061
R6 a_59_75.n0 a_59_75.t4 163.879
R7 a_59_75.n1 a_59_75.n0 76
R8 a_59_75.t0 a_59_75.n2 63.321
R9 a_59_75.n2 a_59_75.t1 63.321
R10 VPWR.n1 VPWR.t2 388.011
R11 VPWR.n1 VPWR.n0 183.665
R12 VPWR.n0 VPWR.t0 116.32
R13 VPWR.n0 VPWR.t1 28.462
R14 VPWR VPWR.n1 0.155
R15 VPB.t0 VPB.t1 319.626
R16 VPB VPB.t2 298.909
R17 VPB.t2 VPB.t0 248.598
R18 X.n0 X.t0 193.162
R19 X X.t1 176.924
R20 X X.n2 11.264
R21 X X.n1 6.656
R22 X.n2 X 6.144
R23 X.n2 X 4.634
R24 X.n1 X.n0 4.077
R25 X.n1 X 3.617
R26 X.n0 X 1.747
R27 a_145_75.t0 a_145_75.t1 77.142
R28 VGND VGND.n0 118.161
R29 VGND.n0 VGND.t0 72.857
R30 VGND.n0 VGND.t1 22.324
R31 VNB VNB.t2 7186.67
R32 VNB.t0 VNB.t1 2650.79
R33 VNB.t2 VNB.t0 2253.66
R34 A.n0 A.t0 256.068
R35 A.n0 A.t1 150.028
R36 A.n1 A.n0 76
R37 A.n2  11.833
R38 A.n1 A 7.68
R39 A.n2 A.n1 4.608
R40 A A.n2 4.588
C0 VPWR X 0.16fF
C1 A SLEEP_B 0.12fF
C2 X VGND 0.15fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__lpflow_inputiso0p_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__lpflow_inputiso0p_1 X SLEEP A VGND VPWR VNB VPB
X0 VPWR.t2 A.t0 a_207_413.t1 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1 X.t0 a_207_413.t3 VPWR.t1 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 a_297_47.t0 a_27_413.t2 a_207_413.t0 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3 X.t1 a_207_413.t4 VGND.t1 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 a_207_413.t2 a_27_413.t3 VPWR.t3 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 VPWR.t0 SLEEP.t0 a_27_413.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 VGND.t2 A.t1 a_297_47.t1 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7 a_27_413.t1 SLEEP.t1 VGND.t0 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
R0 A.n0 A.t1 293.968
R1 A.n0 A.t0 138.336
R2 A.n1 A.n0 76
R3 A A.n1 14.038
R4 A.n1 A 4.954
R5 a_207_413.n2 a_207_413.n1 333.182
R6 a_207_413.n0 a_207_413.t3 240.482
R7 a_207_413.t0 a_207_413.n2 169.75
R8 a_207_413.n0 a_207_413.t4 166.691
R9 a_207_413.n2 a_207_413.n0 98.923
R10 a_207_413.n1 a_207_413.t1 68.011
R11 a_207_413.n1 a_207_413.t2 68.011
R12 VPWR.n9 VPWR.n8 309.954
R13 VPWR.n3 VPWR.n2 292.5
R14 VPWR.n1 VPWR.n0 292.5
R15 VPWR.n8 VPWR.t3 96.154
R16 VPWR.n2 VPWR.t2 86.773
R17 VPWR.n0 VPWR.t1 66.839
R18 VPWR.n8 VPWR.t0 63.321
R19 VPWR.n5 VPWR.n1 5.608
R20 VPWR.n5 VPWR.n4 4.65
R21 VPWR.n7 VPWR.n6 4.65
R22 VPWR.n10 VPWR.n9 3.932
R23 VPWR.n4 VPWR.n3 1
R24 VPWR.n10 VPWR.n7 0.137
R25 VPWR VPWR.n10 0.123
R26 VPWR.n7 VPWR.n5 0.119
R27 VPB.t2 VPB.t1 526.791
R28 VPB.t0 VPB.t3 290.031
R29 VPB.t3 VPB.t2 260.436
R30 VPB VPB.t0 192.367
R31 X.n1 X.t0 212.393
R32 X.n0 X.t1 117.423
R33 X X.n0 79.483
R34 X.n1 X 7.735
R35 X.n0 X 6.666
R36 X X.n1 6.365
R37 a_27_413.t0 a_27_413.n1 433.056
R38 a_27_413.n0 a_27_413.t3 381.656
R39 a_27_413.n0 a_27_413.t2 197.62
R40 a_27_413.n1 a_27_413.t1 151.191
R41 a_27_413.n1 a_27_413.n0 88.993
R42 a_297_47.t0 a_297_47.t1 68.571
R43 VNB VNB.t0 6470.59
R44 VNB.t0 VNB.t2 6082.35
R45 VNB.t2 VNB.t3 2523.53
R46 VNB.t3 VNB.t1 2317.53
R47 VGND.n1 VGND.t0 151.952
R48 VGND.n1 VGND.n0 111.502
R49 VGND.n0 VGND.t2 58.571
R50 VGND.n0 VGND.t1 25.428
R51 VGND VGND.n1 0.045
R52 SLEEP.n0 SLEEP.t0 327.988
R53 SLEEP.n0 SLEEP.t1 199.455
R54 SLEEP.n1 SLEEP.n0 76
R55 SLEEP.n1 SLEEP 12.16
R56 SLEEP SLEEP.n1 2.346
C0 VPWR A 0.15fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__lpflow_inputiso1n_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__lpflow_inputiso1n_1 A SLEEP_B X VGND VPWR VNB VPB
X0 a_219_297.t2 a_27_53.t2 VGND.t3 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1 VGND.t2 SLEEP_B.t0 a_27_53.t0 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 VPWR.t2 A.t0 a_301_297.t1 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3 X.t1 a_219_297.t3 VGND.t0 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 a_301_297.t0 a_27_53.t3 a_219_297.t1 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 X.t0 a_219_297.t4 VPWR.t0 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 a_27_53.t1 SLEEP_B.t1 VPWR.t1 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7 VGND.t1 A.t1 a_219_297.t0 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
R0 a_27_53.n1 a_27_53.t1 379.583
R1 a_27_53.n0 a_27_53.t2 186.028
R2 a_27_53.t0 a_27_53.n1 168.69
R3 a_27_53.n0 a_27_53.t3 137.828
R4 a_27_53.n1 a_27_53.n0 95.393
R5 VGND.n1 VGND.n0 108.687
R6 VGND.n3 VGND.n2 92.5
R7 VGND.n7 VGND.n6 92.5
R8 VGND.n0 VGND.t1 52.857
R9 VGND.n2 VGND.t3 38.571
R10 VGND.n6 VGND.t2 38.571
R11 VGND.n0 VGND.t0 27.568
R12 VGND.n9 VGND.n8 4.65
R13 VGND.n5 VGND.n4 4.65
R14 VGND.n5 VGND.n1 0.864
R15 VGND.n4 VGND.n3 0.196
R16 VGND.n8 VGND.n7 0.196
R17 VGND.n9 VGND.n5 0.119
R18 VGND.n10 VGND.n9 0.119
R19 VGND VGND.n10 0.02
R20 a_219_297.n1 a_219_297.t1 439.31
R21 a_219_297.n0 a_219_297.t4 240.482
R22 a_219_297.n2 a_219_297.n1 171.328
R23 a_219_297.n0 a_219_297.t3 168.182
R24 a_219_297.n1 a_219_297.n0 76
R25 a_219_297.t0 a_219_297.n2 38.571
R26 a_219_297.n2 a_219_297.t2 38.571
R27 VNB VNB.t1 7214.71
R28 VNB.t1 VNB.t2 5823.53
R29 VNB.t2 VNB.t0 2717.65
R30 VNB.t0 VNB.t3 2327.87
R31 SLEEP_B.n0 SLEEP_B.t0 185.375
R32 SLEEP_B.n0 SLEEP_B.t1 137.175
R33 SLEEP_B SLEEP_B.n0 81.632
R34 A A.t0 487.895
R35 A.t0 A.t1 392.026
R36 a_301_297.t0 a_301_297.t1 98.5
R37 VPWR.n1 VPWR.t1 413.04
R38 VPWR.n1 VPWR.n0 173.038
R39 VPWR.n0 VPWR.t2 96.154
R40 VPWR.n0 VPWR.t0 26.595
R41 VPWR VPWR.n1 0.039
R42 VPB.t2 VPB.t0 568.224
R43 VPB.t3 VPB.t1 290.031
R44 VPB.t0 VPB.t3 213.084
R45 VPB VPB.t2 189.408
R46 X X.t0 214.087
R47 X X.t1 194.571
C0 VPWR X 0.13fF
C1 VPWR A 0.25fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__lpflow_inputiso1p_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__lpflow_inputiso1p_1 SLEEP X A VGND VPWR VNB VPB
X0 VGND.t2 SLEEP.t0 a_68_297.t1 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1 a_68_297.t0 A.t0 VGND.t0 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 X.t0 a_68_297.t3 VGND.t1 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 VPWR.t1 SLEEP.t1 a_150_297.t0 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 X.t1 a_68_297.t4 VPWR.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 a_150_297.t1 A.t1 a_68_297.t2 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
R0 SLEEP.n0 SLEEP.t0 206.188
R1 SLEEP.n0 SLEEP.t1 148.348
R2 SLEEP SLEEP.n0 78.656
R3  SLEEP 16.422
R4 a_68_297.n1 a_68_297.t2 370.207
R5 a_68_297.n0 a_68_297.t4 236.179
R6 a_68_297.n2 a_68_297.n1 167.806
R7 a_68_297.n1 a_68_297.n0 165.599
R8 a_68_297.n0 a_68_297.t3 163.879
R9 a_68_297.n2 a_68_297.t1 38.571
R10 a_68_297.t0 a_68_297.n2 38.571
R11 VGND.n1 VGND.t0 158.551
R12 VGND.n1 VGND.n0 123.076
R13 VGND.n0 VGND.t2 55.714
R14 VGND.n0 VGND.t1 26.857
R15 VGND VGND.n1 0.145
R16 VNB VNB.t0 7424.51
R17 VNB.t0 VNB.t2 2717.65
R18 VNB.t2 VNB.t1 2303.7
R19 A.n0 A.t0 192.639
R20 A.n0 A.t1 134.799
R21 A A.n0 77.983
R22  A 12.259
R23 X.n0 X.t1 194.32
R24 X X.t0 128.201
R25 X.n0 X 2.438
R26 X X.n0 1.435
R27 a_150_297.t0 a_150_297.t1 98.5
R28 VPWR VPWR.n0 172.477
R29 VPWR.n0 VPWR.t1 96.154
R30 VPWR.n0 VPWR.t0 25.61
R31 VPB VPB.t2 313.707
R32 VPB.t1 VPB.t0 287.071
R33 VPB.t2 VPB.t1 213.084
C0 X VGND 0.15fF
C1 VPWR X 0.18fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__lpflow_inputisolatch_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__lpflow_inputisolatch_1 SLEEP_B D Q VGND VPWR VNB VPB
X0 a_575_47.t1 a_27_47.t2 a_476_47.t3 VNB.t5 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X1 a_381_369.t0 D.t0 VPWR.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X2 a_476_47.t2 a_27_47.t3 a_381_369.t1 VPB.t5 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3 a_476_47.t0 a_193_47.t2 a_381_47.t0 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X4 VGND.t0 a_629_21.t2 a_575_47.t0 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X5 Q.t0 a_476_47.t4 VGND.t3 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 a_193_47.t1 a_27_47.t4 VPWR.t3 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=550000u l=150000u
X7 a_193_47.t0 a_27_47.t5 VGND.t4 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 VPWR.t5 a_629_21.t3 a_560_413.t1 VPB.t7 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9 VGND.t2 a_476_47.t5 a_629_21.t0 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 Q.t1 a_476_47.t6 VPWR.t2 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 VPWR.t1 a_476_47.t7 a_629_21.t1 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 a_381_47.t1 D.t1 VGND.t1 VNB.t7 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13 VPWR.t4 SLEEP_B.t0 a_27_47.t0 VPB.t6 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=550000u l=150000u
X14 a_560_413.t0 a_193_47.t3 a_476_47.t1 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15 VGND.t5 SLEEP_B.t1 a_27_47.t1 VNB.t6 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
R0 a_27_47.n0 a_27_47.t2 425.944
R1 a_27_47.t0 a_27_47.n3 425.2
R2 a_27_47.n1 a_27_47.n0 280.641
R3 a_27_47.n2 a_27_47.t5 273.133
R4 a_27_47.n1 a_27_47.t4 245.819
R5 a_27_47.n0 a_27_47.t3 219.041
R6 a_27_47.n3 a_27_47.t1 208.264
R7 a_27_47.n3 a_27_47.n2 89.145
R8 a_27_47.n2 a_27_47.n1 38.56
R9 a_476_47.n4 a_476_47.n3 430.17
R10 a_476_47.n0 a_476_47.t6 212.079
R11 a_476_47.n1 a_476_47.t7 212.079
R12 a_476_47.n3 a_476_47.n2 188.122
R13 a_476_47.n3 a_476_47.n1 167.966
R14 a_476_47.n0 a_476_47.t4 139.779
R15 a_476_47.n1 a_476_47.t5 139.779
R16 a_476_47.n2 a_476_47.t0 68.333
R17 a_476_47.t1 a_476_47.n4 63.321
R18 a_476_47.n4 a_476_47.t2 63.321
R19 a_476_47.n1 a_476_47.n0 61.345
R20 a_476_47.n2 a_476_47.t3 46.666
R21 a_575_47.t0 a_575_47.t1 90
R22 VNB.t4 VNB.t7 6082.35
R23 VNB.t0 VNB.t2 5690.29
R24 VNB VNB.t6 4270.59
R25 VNB.t1 VNB.t5 3512.9
R26 VNB.t7 VNB.t1 3011.81
R27 VNB.t5 VNB.t0 2980.65
R28 VNB.t6 VNB.t4 2717.65
R29 VNB.t2 VNB.t3 2030.77
R30 D.n0 D.t0 373.281
R31 D.n0 D.t1 127.283
R32 D D.n0 79.242
R33 VPWR.n9 VPWR.t0 425.096
R34 VPWR.n1 VPWR.t5 385.734
R35 VPWR.n15 VPWR.n14 311.893
R36 VPWR.n2 VPWR.n0 183.831
R37 VPWR.n14 VPWR.t3 48.354
R38 VPWR.n14 VPWR.t4 48.354
R39 VPWR.n0 VPWR.t2 26.595
R40 VPWR.n0 VPWR.t1 26.595
R41 VPWR.n2 VPWR.n1 4.845
R42 VPWR.n4 VPWR.n3 4.65
R43 VPWR.n6 VPWR.n5 4.65
R44 VPWR.n8 VPWR.n7 4.65
R45 VPWR.n11 VPWR.n10 4.65
R46 VPWR.n13 VPWR.n12 4.65
R47 VPWR.n16 VPWR.n15 3.932
R48 VPWR.n10 VPWR.n9 0.232
R49 VPWR.n4 VPWR.n2 0.18
R50 VPWR.n16 VPWR.n13 0.137
R51 VPWR VPWR.n16 0.123
R52 VPWR.n6 VPWR.n4 0.119
R53 VPWR.n8 VPWR.n6 0.119
R54 VPWR.n11 VPWR.n8 0.119
R55 VPWR.n13 VPWR.n11 0.119
R56 a_381_369.t0 a_381_369.t1 132.285
R57 VPB.t7 VPB.t2 562.305
R58 VPB.t4 VPB.t0 556.386
R59 VPB.t1 VPB.t7 292.99
R60 VPB.t0 VPB.t5 281.152
R61 VPB.t2 VPB.t3 248.598
R62 VPB.t5 VPB.t1 248.598
R63 VPB.t6 VPB.t4 248.598
R64 VPB VPB.t6 142.056
R65 a_193_47.t1 a_193_47.n1 354.03
R66 a_193_47.n0 a_193_47.t2 252.105
R67 a_193_47.n1 a_193_47.t0 241.336
R68 a_193_47.n0 a_193_47.t3 224.251
R69 a_193_47.n1 a_193_47.n0 109.176
R70 a_381_47.n0 a_381_47.t0 66.666
R71 a_381_47.n0 a_381_47.t1 26.393
R72 a_381_47.n1 a_381_47.n0 14.4
R73 a_629_21.t1 a_629_21.n2 466.769
R74 a_629_21.n1 a_629_21.t2 375.959
R75 a_629_21.n0 a_629_21.t0 184.62
R76 a_629_21.n1 a_629_21.t3 147.812
R77 a_629_21.n2 a_629_21.n1 93.648
R78 a_629_21.n2 a_629_21.n0 0.775
R79 VGND.n1 VGND.t0 154.76
R80 VGND.n9 VGND.t1 145.81
R81 VGND.n2 VGND.n0 131.996
R82 VGND.n14 VGND.n13 107.239
R83 VGND.n13 VGND.t4 38.571
R84 VGND.n13 VGND.t5 38.571
R85 VGND.n0 VGND.t3 24.923
R86 VGND.n0 VGND.t2 24.923
R87 VGND.n4 VGND.n3 4.65
R88 VGND.n6 VGND.n5 4.65
R89 VGND.n8 VGND.n7 4.65
R90 VGND.n10 VGND.n9 4.65
R91 VGND.n12 VGND.n11 4.65
R92 VGND.n15 VGND.n14 3.932
R93 VGND.n2 VGND.n1 3.907
R94 VGND.n4 VGND.n2 0.2
R95 VGND.n15 VGND.n12 0.137
R96 VGND VGND.n15 0.123
R97 VGND.n6 VGND.n4 0.119
R98 VGND.n8 VGND.n6 0.119
R99 VGND.n10 VGND.n8 0.119
R100 VGND.n12 VGND.n10 0.119
R101 Q.n0 Q.t1 226.977
R102 Q.n1 Q.t0 117.423
R103 Q Q.n1 82.221
R104 Q Q.n0 7.813
R105 Q.n0 Q 7.279
R106 Q.n1 Q 6.961
R107 a_560_413.t0 a_560_413.t1 161.821
R108 SLEEP_B.n0 SLEEP_B.t0 284.913
R109 SLEEP_B.n0 SLEEP_B.t1 235.108
R110 SLEEP_B SLEEP_B.n0 78.1
C0 VPWR Q 0.14fF
C1 VPB VPWR 0.10fF
C2 VPWR VGND 0.12fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__lpflow_isobufsrc_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__lpflow_isobufsrc_1 A X SLEEP VGND VPWR VNB VPB
X0 X.t2 a_74_47.t2 a_265_297.t1 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 VPWR.t1 A.t0 a_74_47.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 a_265_297.t0 SLEEP.t0 VPWR.t0 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 X.t0 SLEEP.t1 VGND.t1 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 VGND.t0 A.t1 a_74_47.t1 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 VGND.t2 a_74_47.t3 X.t1 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
R0 a_74_47.t0 a_74_47.n1 362.467
R1 a_74_47.n0 a_74_47.t2 236.179
R2 a_74_47.n1 a_74_47.t1 210.277
R3 a_74_47.n1 a_74_47.n0 170.4
R4 a_74_47.n0 a_74_47.t3 163.879
R5 a_265_297.t0 a_265_297.t1 41.37
R6 X.n1 X.t2 173.353
R7 X.n1 X.n0 166.613
R8 X.n0 X.t1 24.923
R9 X.n0 X.t0 24.923
R10 X X.n1 1.434
R11 VPB VPB.t0 334.423
R12 VPB.t0 VPB.t1 319.626
R13 VPB.t1 VPB.t2 213.084
R14 A.n0 A.t1 176.733
R15 A A.n0 147.046
R16 A.n0 A.t0 119.623
R17  A 19.342
R18 VPWR VPWR.n0 169.473
R19 VPWR.n0 VPWR.t1 121.952
R20 VPWR.n0 VPWR.t0 25.61
R21 SLEEP.n0 SLEEP.t0 236.179
R22 SLEEP.n0 SLEEP.t1 163.879
R23 SLEEP SLEEP.n0 80.676
R24 VGND.n1 VGND.t2 187.535
R25 VGND.n1 VGND.n0 81.179
R26 VGND.n0 VGND.t0 57.772
R27 VGND.n0 VGND.t1 24.789
R28 VGND VGND.n1 0.295
R29 VNB VNB.t0 8355.68
R30 VNB.t0 VNB.t1 2303.7
R31 VNB.t1 VNB.t2 2030.77
C0 X VGND 0.33fF
C1 VPWR X 0.14fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__lpflow_isobufsrc_2.ext - technology: sky130A

.subckt sky130_fd_sc_hd__lpflow_isobufsrc_2 A SLEEP X VGND VPWR VNB VPB
X0 X.t3 a_251_21.t2 a_27_297.t3 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 X.t5 a_251_21.t3 VGND.t4 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 a_27_297.t0 SLEEP.t0 VPWR.t2 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 VGND.t1 SLEEP.t1 X.t0 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 X.t1 SLEEP.t2 VGND.t2 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 VGND.t3 a_251_21.t4 X.t4 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 VPWR.t1 SLEEP.t3 a_27_297.t1 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 VPWR.t0 A.t0 a_251_21.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 VGND.t0 A.t1 a_251_21.t1 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9 a_27_297.t2 a_251_21.t5 X.t2 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
R0 a_251_21.t0 a_251_21.n2 433.143
R1 a_251_21.n1 a_251_21.t5 212.079
R2 a_251_21.n0 a_251_21.t2 212.079
R3 a_251_21.n2 a_251_21.t1 156.452
R4 a_251_21.n1 a_251_21.t4 139.779
R5 a_251_21.n0 a_251_21.t3 139.779
R6 a_251_21.n2 a_251_21.n1 131.533
R7 a_251_21.n1 a_251_21.n0 61.345
R8 a_27_297.n0 a_27_297.t2 200.245
R9 a_27_297.n0 a_27_297.t1 190.115
R10 a_27_297.n1 a_27_297.n0 90.234
R11 a_27_297.n1 a_27_297.t3 26.595
R12 a_27_297.t0 a_27_297.n1 26.595
R13 X.n2 X.n1 190.893
R14 X X.n4 93.857
R15 X.n2 X.n0 90.831
R16 X.n1 X.t2 26.595
R17 X.n1 X.t3 26.595
R18 X.n4 X.t4 24.923
R19 X.n4 X.t5 24.923
R20 X.n0 X.t0 24.923
R21 X.n0 X.t1 24.923
R22 X X.n3 11.83
R23 X.n3 X.n2 3.103
R24 VPB.t3 VPB.t0 556.386
R25 VPB.t4 VPB.t3 248.598
R26 VPB.t1 VPB.t4 248.598
R27 VPB.t2 VPB.t1 248.598
R28 VPB VPB.t2 201.246
R29 VGND.n1 VGND.t0 169.161
R30 VGND.n5 VGND.n4 115.464
R31 VGND.n0 VGND.t3 114.4
R32 VGND.n10 VGND.t2 104.882
R33 VGND.n4 VGND.t4 24.923
R34 VGND.n4 VGND.t1 24.923
R35 VGND.n1 VGND.n0 12.335
R36 VGND.n11 VGND.n10 4.65
R37 VGND.n3 VGND.n2 4.65
R38 VGND.n7 VGND.n6 4.65
R39 VGND.n9 VGND.n8 4.65
R40 VGND.n6 VGND.n5 2.258
R41 VGND.n3 VGND.n1 0.218
R42 VGND.n7 VGND.n3 0.119
R43 VGND.n9 VGND.n7 0.119
R44 VGND.n11 VGND.n9 0.119
R45 VGND VGND.n11 0.02
R46 VNB VNB.t2 6150.61
R47 VNB.t3 VNB.t0 5321.88
R48 VNB.t4 VNB.t3 2030.77
R49 VNB.t1 VNB.t4 2030.77
R50 VNB.t2 VNB.t1 2030.77
R51 SLEEP.n0 SLEEP.t0 212.079
R52 SLEEP.n1 SLEEP.t3 212.079
R53 SLEEP.n0 SLEEP.t1 139.779
R54 SLEEP.n1 SLEEP.t2 139.779
R55 SLEEP SLEEP.n2 77.6
R56 SLEEP.n2 SLEEP.n0 38.706
R57 SLEEP.n2 SLEEP.n1 22.639
R58 VPWR.n1 VPWR.t0 381.226
R59 VPWR.n1 VPWR.n0 173.445
R60 VPWR.n0 VPWR.t2 26.595
R61 VPWR.n0 VPWR.t1 26.595
R62 VPWR VPWR.n1 0.142
R63 A.n0 A.t0 333.171
R64 A.n0 A.t1 130.731
R65 A.n1 A.n0 84.838
R66  A.n1 16.372
R67 A.n1 A 3.869
C0 X VGND 0.49fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__lpflow_isobufsrc_4.ext - technology: sky130A

.subckt sky130_fd_sc_hd__lpflow_isobufsrc_4 A X SLEEP VGND VPWR VNB VPB
X0 VPWR.t4 SLEEP.t0 a_27_297.t4 VPB.t5 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 X.t4 SLEEP.t1 VGND.t4 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 a_27_297.t3 SLEEP.t2 VPWR.t3 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 VGND.t3 SLEEP.t3 X.t3 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 a_27_297.t5 a_419_21.t2 X.t5 VPB.t6 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 X.t2 SLEEP.t4 VGND.t2 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 VGND.t1 SLEEP.t5 X.t1 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 VGND.t5 a_419_21.t3 X.t6 VNB.t5 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 VGND.t6 a_419_21.t4 X.t7 VNB.t6 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 X.t8 a_419_21.t5 a_27_297.t6 VPB.t7 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 VPWR.t2 SLEEP.t6 a_27_297.t2 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 X.t9 a_419_21.t6 VGND.t7 VNB.t7 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 VGND.t0 A.t0 a_419_21.t0 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 X.t10 a_419_21.t7 VGND.t8 VNB.t8 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14 VPWR.t0 A.t1 a_419_21.t1 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 a_27_297.t7 a_419_21.t8 X.t11 VPB.t8 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16 X.t0 a_419_21.t9 a_27_297.t0 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17 a_27_297.t1 SLEEP.t7 VPWR.t1 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
R0 SLEEP.n0 SLEEP.t7 212.079
R1 SLEEP.n2 SLEEP.t0 212.079
R2 SLEEP.n5 SLEEP.t2 212.079
R3 SLEEP.n8 SLEEP.t6 212.079
R4 SLEEP.n0 SLEEP.t5 139.779
R5 SLEEP.n2 SLEEP.t1 139.779
R6 SLEEP.n5 SLEEP.t3 139.779
R7 SLEEP.n8 SLEEP.t4 139.779
R8 SLEEP.n4 SLEEP.n1 97.76
R9 SLEEP SLEEP.n9 76.64
R10 SLEEP.n4 SLEEP.n3 76
R11 SLEEP.n7 SLEEP.n6 76
R12 SLEEP.n7 SLEEP.n4 21.76
R13 SLEEP SLEEP.n7 21.12
R14 SLEEP.n1 SLEEP.n0 18.987
R15 SLEEP.n9 SLEEP.n8 16.066
R16 SLEEP.n3 SLEEP.n2 7.303
R17 SLEEP.n6 SLEEP.n5 4.381
R18 a_27_297.n3 a_27_297.t2 181.085
R19 a_27_297.n1 a_27_297.t5 169.982
R20 a_27_297.n1 a_27_297.n0 150.25
R21 a_27_297.n3 a_27_297.n2 109.334
R22 a_27_297.n5 a_27_297.n4 91.601
R23 a_27_297.n4 a_27_297.n3 57.04
R24 a_27_297.n4 a_27_297.n1 53.037
R25 a_27_297.n2 a_27_297.t4 26.595
R26 a_27_297.n2 a_27_297.t3 26.595
R27 a_27_297.n0 a_27_297.t6 26.595
R28 a_27_297.n0 a_27_297.t7 26.595
R29 a_27_297.t0 a_27_297.n5 26.595
R30 a_27_297.n5 a_27_297.t1 26.595
R31 VPWR.n1 VPWR.n0 169.933
R32 VPWR.n6 VPWR.n5 164.214
R33 VPWR.n2 VPWR.t0 146.245
R34 VPWR.n0 VPWR.t1 26.595
R35 VPWR.n0 VPWR.t4 26.595
R36 VPWR.n5 VPWR.t3 26.595
R37 VPWR.n5 VPWR.t2 26.595
R38 VPWR.n4 VPWR.n3 4.65
R39 VPWR.n2 VPWR.n1 4.126
R40 VPWR.n7 VPWR.n6 3.966
R41 VPWR.n7 VPWR.n4 0.137
R42 VPWR.n4 VPWR.n2 0.134
R43 VPWR VPWR.n7 0.122
R44 VPB.t6 VPB.t0 574.143
R45 VPB.t7 VPB.t6 248.598
R46 VPB.t8 VPB.t7 248.598
R47 VPB.t1 VPB.t8 248.598
R48 VPB.t2 VPB.t1 248.598
R49 VPB.t5 VPB.t2 248.598
R50 VPB.t4 VPB.t5 248.598
R51 VPB.t3 VPB.t4 248.598
R52 VPB VPB.t3 201.246
R53 VGND.n5 VGND.n4 115.464
R54 VGND.n11 VGND.n10 115.464
R55 VGND.n17 VGND.n16 115.464
R56 VGND.n1 VGND.t0 109.099
R57 VGND.n0 VGND.t6 106.289
R58 VGND.n22 VGND.t2 104.219
R59 VGND.n4 VGND.t8 24.923
R60 VGND.n4 VGND.t5 24.923
R61 VGND.n10 VGND.t7 24.923
R62 VGND.n10 VGND.t1 24.923
R63 VGND.n16 VGND.t4 24.923
R64 VGND.n16 VGND.t3 24.923
R65 VGND.n6 VGND.n5 14.305
R66 VGND.n1 VGND.n0 8.896
R67 VGND.n12 VGND.n11 8.282
R68 VGND.n23 VGND.n22 4.65
R69 VGND.n3 VGND.n2 4.65
R70 VGND.n7 VGND.n6 4.65
R71 VGND.n9 VGND.n8 4.65
R72 VGND.n13 VGND.n12 4.65
R73 VGND.n15 VGND.n14 4.65
R74 VGND.n19 VGND.n18 4.65
R75 VGND.n21 VGND.n20 4.65
R76 VGND.n18 VGND.n17 2.258
R77 VGND.n3 VGND.n1 0.266
R78 VGND.n7 VGND.n3 0.119
R79 VGND.n9 VGND.n7 0.119
R80 VGND.n13 VGND.n9 0.119
R81 VGND.n15 VGND.n13 0.119
R82 VGND.n19 VGND.n15 0.119
R83 VGND.n21 VGND.n19 0.119
R84 VGND.n23 VGND.n21 0.119
R85 VGND VGND.n23 0.02
R86 X X.n0 163.414
R87 X.n9 X.n1 152.296
R88 X.n8 X.n2 94.934
R89 X.n6 X.n4 88.89
R90 X.n6 X.n5 52.624
R91 X.n7 X.n3 49.285
R92 X.n7 X.n6 47.999
R93 X.n9 X.n8 26.763
R94 X.n0 X.t5 26.595
R95 X.n0 X.t8 26.595
R96 X.n1 X.t11 26.595
R97 X.n1 X.t0 26.595
R98 X.n3 X.t6 24.923
R99 X.n3 X.t9 24.923
R100 X.n4 X.t3 24.923
R101 X.n4 X.t2 24.923
R102 X.n5 X.t1 24.923
R103 X.n5 X.t4 24.923
R104 X.n2 X.t7 24.923
R105 X.n2 X.t10 24.923
R106 X X.n9 12.16
R107 X.n8 X.n7 5.688
R108 VNB VNB.t2 6150.61
R109 VNB.t6 VNB.t0 4690.11
R110 VNB.t8 VNB.t6 2030.77
R111 VNB.t5 VNB.t8 2030.77
R112 VNB.t7 VNB.t5 2030.77
R113 VNB.t1 VNB.t7 2030.77
R114 VNB.t4 VNB.t1 2030.77
R115 VNB.t3 VNB.t4 2030.77
R116 VNB.t2 VNB.t3 2030.77
R117 a_419_21.n6 a_419_21.t2 212.079
R118 a_419_21.n0 a_419_21.t5 212.079
R119 a_419_21.n2 a_419_21.t8 212.079
R120 a_419_21.n1 a_419_21.t9 212.079
R121 a_419_21.t1 a_419_21.n8 154.904
R122 a_419_21.n6 a_419_21.t4 139.779
R123 a_419_21.n0 a_419_21.t7 139.779
R124 a_419_21.n2 a_419_21.t3 139.779
R125 a_419_21.n1 a_419_21.t6 139.779
R126 a_419_21.n8 a_419_21.t0 107.578
R127 a_419_21.n4 a_419_21.n3 97.76
R128 a_419_21.n7 a_419_21.n6 73.418
R129 a_419_21.n2 a_419_21.n1 61.345
R130 a_419_21.n3 a_419_21.n2 54.042
R131 a_419_21.n7 a_419_21.n4 29.163
R132 a_419_21.n6 a_419_21.n5 18.987
R133 a_419_21.n8 a_419_21.n7 15.119
R134 a_419_21.n3 a_419_21.n0 7.303
R135 A.n0 A.t1 229.752
R136 A.n0 A.t0 157.452
R137 A A.n0 83.314
C0 X VGND 0.92fF
C1 VPB VPWR 0.11fF
C2 VPWR VGND 0.11fF
C3 A VPWR 0.11fF
C4 SLEEP X 0.25fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__lpflow_isobufsrc_8.ext - technology: sky130A

.subckt sky130_fd_sc_hd__lpflow_isobufsrc_8 A X SLEEP VGND VPWR VNB VPB
X0 X.t7 a_123_297.t4 VGND.t7 VNB sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 X.t6 a_123_297.t5 VGND.t6 VNB sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 a_321_297.t7 a_123_297.t6 VPWR.t7 VPB.t7 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 X.t5 a_123_297.t7 VGND.t5 VNB sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 VPWR.t6 a_123_297.t8 a_321_297.t6 VPB.t6 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 a_321_297.t8 SLEEP.t0 X.t8 VPB.t8 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 a_123_297.t0 A.t0 VGND.t16 VNB sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 a_321_297.t5 a_123_297.t9 VPWR.t5 VPB.t5 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 X.t9 SLEEP.t1 a_321_297.t9 VPB.t9 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 VGND.t4 a_123_297.t10 X.t4 VNB sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 VGND.t8 SLEEP.t2 X.t10 VNB sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 VGND.t9 SLEEP.t3 X.t11 VNB sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 VPWR.t4 a_123_297.t11 a_321_297.t4 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13 a_321_297.t10 SLEEP.t4 X.t12 VPB.t10 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14 VGND.t3 a_123_297.t12 X.t3 VNB sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X15 a_123_297.t1 A.t1 VPWR.t8 VPB.t16 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16 VGND.t2 a_123_297.t13 X.t2 VNB sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X17 a_321_297.t3 a_123_297.t14 VPWR.t3 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X18 VGND.t17 A.t2 a_123_297.t2 VNB sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X19 X.t13 SLEEP.t5 a_321_297.t11 VPB.t11 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X20 X.t14 SLEEP.t6 VGND.t10 VNB sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X21 VPWR.t2 a_123_297.t15 a_321_297.t2 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X22 X.t15 SLEEP.t7 VGND.t11 VNB sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X23 a_321_297.t12 SLEEP.t8 X.t16 VPB.t12 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X24 X.t17 SLEEP.t9 VGND.t12 VNB sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X25 a_321_297.t1 a_123_297.t16 VPWR.t1 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X26 X.t18 SLEEP.t10 a_321_297.t13 VPB.t13 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X27 X.t19 SLEEP.t11 VGND.t13 VNB sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X28 a_321_297.t14 SLEEP.t12 X.t20 VPB.t14 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X29 VGND.t1 a_123_297.t17 X.t1 VNB sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X30 X.t21 SLEEP.t13 a_321_297.t15 VPB.t15 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X31 VGND.t14 SLEEP.t14 X.t22 VNB sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X32 VGND.t15 SLEEP.t15 X.t23 VNB sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X33 VPWR.t9 A.t3 a_123_297.t3 VPB.t17 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X34 VPWR.t0 a_123_297.t18 a_321_297.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X35 X.t0 a_123_297.t19 VGND.t0 VNB sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
R0 a_123_297.n1 a_123_297.t14 212.079
R1 a_123_297.n3 a_123_297.t15 212.079
R2 a_123_297.n6 a_123_297.t16 212.079
R3 a_123_297.n11 a_123_297.t18 212.079
R4 a_123_297.n14 a_123_297.t6 212.079
R5 a_123_297.n17 a_123_297.t8 212.079
R6 a_123_297.n20 a_123_297.t9 212.079
R7 a_123_297.n23 a_123_297.t11 212.079
R8 a_123_297.n1 a_123_297.t13 139.779
R9 a_123_297.n3 a_123_297.t7 139.779
R10 a_123_297.n6 a_123_297.t12 139.779
R11 a_123_297.n11 a_123_297.t5 139.779
R12 a_123_297.n14 a_123_297.t10 139.779
R13 a_123_297.n17 a_123_297.t4 139.779
R14 a_123_297.n20 a_123_297.t17 139.779
R15 a_123_297.n23 a_123_297.t19 139.779
R16 a_123_297.n27 a_123_297.n26 133.042
R17 a_123_297.n5 a_123_297.n2 96.723
R18 a_123_297.n25 a_123_297.n24 76
R19 a_123_297.n5 a_123_297.n4 76
R20 a_123_297.n8 a_123_297.n7 76
R21 a_123_297.n10 a_123_297.n9 76
R22 a_123_297.n13 a_123_297.n12 76
R23 a_123_297.n16 a_123_297.n15 76
R24 a_123_297.n19 a_123_297.n18 76
R25 a_123_297.n22 a_123_297.n21 76
R26 a_123_297.n26 a_123_297.n25 65.371
R27 a_123_297.n26 a_123_297.n0 62.321
R28 a_123_297.n12 a_123_297.n11 30.672
R29 a_123_297.n27 a_123_297.t3 26.595
R30 a_123_297.t1 a_123_297.n27 26.595
R31 a_123_297.n0 a_123_297.t2 24.923
R32 a_123_297.n0 a_123_297.t0 24.923
R33 a_123_297.n8 a_123_297.n5 20.723
R34 a_123_297.n10 a_123_297.n8 20.723
R35 a_123_297.n13 a_123_297.n10 20.723
R36 a_123_297.n16 a_123_297.n13 20.723
R37 a_123_297.n19 a_123_297.n16 20.723
R38 a_123_297.n22 a_123_297.n19 20.723
R39 a_123_297.n25 a_123_297.n22 20.723
R40 a_123_297.n15 a_123_297.n14 18.987
R41 a_123_297.n2 a_123_297.n1 16.066
R42 a_123_297.n24 a_123_297.n23 16.066
R43 a_123_297.n7 a_123_297.n6 7.303
R44 a_123_297.n18 a_123_297.n17 7.303
R45 a_123_297.n4 a_123_297.n3 4.381
R46 a_123_297.n21 a_123_297.n20 4.381
R47 VGND.n0 VGND.t15 192.923
R48 VGND.n2 VGND.n1 115.464
R49 VGND.n8 VGND.n7 115.464
R50 VGND.n14 VGND.n13 115.464
R51 VGND.n18 VGND.n17 115.464
R52 VGND.n24 VGND.n23 115.464
R53 VGND.n30 VGND.n29 115.464
R54 VGND.n36 VGND.n35 115.464
R55 VGND.n46 VGND.t16 112.846
R56 VGND.n41 VGND.t0 56.307
R57 VGND.n41 VGND.t17 56.307
R58 VGND.n1 VGND.t13 24.923
R59 VGND.n1 VGND.t14 24.923
R60 VGND.n7 VGND.t12 24.923
R61 VGND.n7 VGND.t9 24.923
R62 VGND.n13 VGND.t11 24.923
R63 VGND.n13 VGND.t8 24.923
R64 VGND.n17 VGND.t10 24.923
R65 VGND.n17 VGND.t2 24.923
R66 VGND.n23 VGND.t5 24.923
R67 VGND.n23 VGND.t3 24.923
R68 VGND.n29 VGND.t6 24.923
R69 VGND.n29 VGND.t4 24.923
R70 VGND.n35 VGND.t7 24.923
R71 VGND.n35 VGND.t1 24.923
R72 VGND.n15 VGND.n14 15.058
R73 VGND.n42 VGND.n41 14.054
R74 VGND.n19 VGND.n18 13.552
R75 VGND.n9 VGND.n8 9.035
R76 VGND.n25 VGND.n24 7.529
R77 VGND.n4 VGND.n3 4.65
R78 VGND.n6 VGND.n5 4.65
R79 VGND.n10 VGND.n9 4.65
R80 VGND.n12 VGND.n11 4.65
R81 VGND.n16 VGND.n15 4.65
R82 VGND.n20 VGND.n19 4.65
R83 VGND.n22 VGND.n21 4.65
R84 VGND.n26 VGND.n25 4.65
R85 VGND.n28 VGND.n27 4.65
R86 VGND.n32 VGND.n31 4.65
R87 VGND.n34 VGND.n33 4.65
R88 VGND.n38 VGND.n37 4.65
R89 VGND.n40 VGND.n39 4.65
R90 VGND.n43 VGND.n42 4.65
R91 VGND.n45 VGND.n44 4.65
R92 VGND.n48 VGND.n47 4.65
R93 VGND.n37 VGND.n36 4.517
R94 VGND.n3 VGND.n2 3.011
R95 VGND.n47 VGND.n46 2.635
R96 VGND.n31 VGND.n30 1.505
R97 VGND.n4 VGND.n0 0.76
R98 VGND.n6 VGND.n4 0.119
R99 VGND.n10 VGND.n6 0.119
R100 VGND.n12 VGND.n10 0.119
R101 VGND.n16 VGND.n12 0.119
R102 VGND.n20 VGND.n16 0.119
R103 VGND.n22 VGND.n20 0.119
R104 VGND.n26 VGND.n22 0.119
R105 VGND.n28 VGND.n26 0.119
R106 VGND.n32 VGND.n28 0.119
R107 VGND.n34 VGND.n32 0.119
R108 VGND.n38 VGND.n34 0.119
R109 VGND.n40 VGND.n38 0.119
R110 VGND.n43 VGND.n40 0.119
R111 VGND.n45 VGND.n43 0.119
R112 VGND.n48 VGND.n45 0.119
R113 VGND.n49 VGND.n48 0.119
R114 VGND VGND.n49 0.022
R115 X.n2 X.n0 199.508
R116 X.n2 X.n1 155.085
R117 X.n4 X.n3 155.085
R118 X.n6 X.n5 155.085
R119 X.n10 X.n8 88.89
R120 X.n10 X.n9 52.624
R121 X.n12 X.n11 52.624
R122 X.n14 X.n13 52.624
R123 X.n16 X.n15 52.624
R124 X.n18 X.n17 52.624
R125 X.n20 X.n19 52.624
R126 X.n21 X.n7 49.285
R127 X.n21 X.n20 47.999
R128 X.n4 X.n2 44.423
R129 X.n6 X.n4 44.423
R130 X X.n21 40.506
R131 X.n12 X.n10 36.266
R132 X.n14 X.n12 36.266
R133 X.n16 X.n14 36.266
R134 X.n18 X.n16 36.266
R135 X.n20 X.n18 36.266
R136 X.n0 X.t12 26.595
R137 X.n0 X.t13 26.595
R138 X.n1 X.t8 26.595
R139 X.n1 X.t9 26.595
R140 X.n3 X.t20 26.595
R141 X.n3 X.t21 26.595
R142 X.n5 X.t16 26.595
R143 X.n5 X.t18 26.595
R144 X.n7 X.t23 24.923
R145 X.n7 X.t19 24.923
R146 X.n8 X.t1 24.923
R147 X.n8 X.t0 24.923
R148 X.n9 X.t4 24.923
R149 X.n9 X.t7 24.923
R150 X.n11 X.t3 24.923
R151 X.n11 X.t6 24.923
R152 X.n13 X.t2 24.923
R153 X.n13 X.t5 24.923
R154 X.n15 X.t10 24.923
R155 X.n15 X.t14 24.923
R156 X.n17 X.t11 24.923
R157 X.n17 X.t15 24.923
R158 X.n19 X.t22 24.923
R159 X.n19 X.t17 24.923
R160 X X.n6 2.666
R161 VPWR.n3 VPWR.n0 174.105
R162 VPWR.n12 VPWR.n11 169.933
R163 VPWR.n7 VPWR.n6 169.933
R164 VPWR.n2 VPWR.n1 169.933
R165 VPWR.n20 VPWR.t8 156.829
R166 VPWR.n16 VPWR.t9 153.549
R167 VPWR.n11 VPWR.t5 26.595
R168 VPWR.n11 VPWR.t4 26.595
R169 VPWR.n6 VPWR.t7 26.595
R170 VPWR.n6 VPWR.t6 26.595
R171 VPWR.n1 VPWR.t1 26.595
R172 VPWR.n1 VPWR.t0 26.595
R173 VPWR.n0 VPWR.t3 26.595
R174 VPWR.n0 VPWR.t2 26.595
R175 VPWR.n5 VPWR.n4 4.65
R176 VPWR.n8 VPWR.n7 4.65
R177 VPWR.n10 VPWR.n9 4.65
R178 VPWR.n13 VPWR.n12 4.65
R179 VPWR.n15 VPWR.n14 4.65
R180 VPWR.n17 VPWR.n16 4.65
R181 VPWR.n19 VPWR.n18 4.65
R182 VPWR.n21 VPWR.n20 4.65
R183 VPWR.n3 VPWR.n2 3.948
R184 VPWR.n5 VPWR.n3 0.257
R185 VPWR.n8 VPWR.n5 0.119
R186 VPWR.n10 VPWR.n8 0.119
R187 VPWR.n13 VPWR.n10 0.119
R188 VPWR.n15 VPWR.n13 0.119
R189 VPWR.n17 VPWR.n15 0.119
R190 VPWR.n19 VPWR.n17 0.119
R191 VPWR.n21 VPWR.n19 0.119
R192 VPWR VPWR.n21 0.022
R193 a_321_297.n4 a_321_297.t12 225.591
R194 a_321_297.n1 a_321_297.t4 169.699
R195 a_321_297.n4 a_321_297.n3 154.573
R196 a_321_297.n6 a_321_297.n5 154.573
R197 a_321_297.n8 a_321_297.n7 154.573
R198 a_321_297.n13 a_321_297.n12 109.737
R199 a_321_297.n11 a_321_297.n10 109.736
R200 a_321_297.n1 a_321_297.n0 109.736
R201 a_321_297.n9 a_321_297.n2 90.234
R202 a_321_297.n9 a_321_297.n8 64.95
R203 a_321_297.n11 a_321_297.n9 55.464
R204 a_321_297.n6 a_321_297.n4 44.423
R205 a_321_297.n8 a_321_297.n6 44.423
R206 a_321_297.n12 a_321_297.n1 35.961
R207 a_321_297.n12 a_321_297.n11 35.961
R208 a_321_297.n2 a_321_297.t11 26.595
R209 a_321_297.n2 a_321_297.t3 26.595
R210 a_321_297.n3 a_321_297.t13 26.595
R211 a_321_297.n3 a_321_297.t14 26.595
R212 a_321_297.n5 a_321_297.t15 26.595
R213 a_321_297.n5 a_321_297.t8 26.595
R214 a_321_297.n7 a_321_297.t9 26.595
R215 a_321_297.n7 a_321_297.t10 26.595
R216 a_321_297.n10 a_321_297.t2 26.595
R217 a_321_297.n10 a_321_297.t1 26.595
R218 a_321_297.n0 a_321_297.t6 26.595
R219 a_321_297.n0 a_321_297.t5 26.595
R220 a_321_297.n13 a_321_297.t0 26.595
R221 a_321_297.t7 a_321_297.n13 26.595
R222 VPB.t17 VPB.t4 591.9
R223 VPB.t13 VPB.t12 248.598
R224 VPB.t14 VPB.t13 248.598
R225 VPB.t15 VPB.t14 248.598
R226 VPB.t8 VPB.t15 248.598
R227 VPB.t9 VPB.t8 248.598
R228 VPB.t10 VPB.t9 248.598
R229 VPB.t11 VPB.t10 248.598
R230 VPB.t3 VPB.t11 248.598
R231 VPB.t2 VPB.t3 248.598
R232 VPB.t1 VPB.t2 248.598
R233 VPB.t0 VPB.t1 248.598
R234 VPB.t7 VPB.t0 248.598
R235 VPB.t6 VPB.t7 248.598
R236 VPB.t5 VPB.t6 248.598
R237 VPB.t4 VPB.t5 248.598
R238 VPB.t16 VPB.t17 248.598
R239 VPB VPB.t16 233.8
R240 SLEEP.n0 SLEEP.t8 212.079
R241 SLEEP.n1 SLEEP.t10 212.079
R242 SLEEP.n2 SLEEP.t12 212.079
R243 SLEEP.n6 SLEEP.t13 212.079
R244 SLEEP.n9 SLEEP.t0 212.079
R245 SLEEP.n12 SLEEP.t1 212.079
R246 SLEEP.n15 SLEEP.t4 212.079
R247 SLEEP.n18 SLEEP.t5 212.079
R248 SLEEP.n0 SLEEP.t15 139.779
R249 SLEEP.n1 SLEEP.t11 139.779
R250 SLEEP.n2 SLEEP.t14 139.779
R251 SLEEP.n6 SLEEP.t9 139.779
R252 SLEEP.n9 SLEEP.t3 139.779
R253 SLEEP.n12 SLEEP.t7 139.779
R254 SLEEP.n15 SLEEP.t2 139.779
R255 SLEEP.n18 SLEEP.t6 139.779
R256 SLEEP SLEEP.n19 90.08
R257 SLEEP.n5 SLEEP.n4 76
R258 SLEEP.n8 SLEEP.n7 76
R259 SLEEP.n11 SLEEP.n10 76
R260 SLEEP.n14 SLEEP.n13 76
R261 SLEEP.n17 SLEEP.n16 76
R262 SLEEP.n1 SLEEP.n0 61.345
R263 SLEEP.n5 SLEEP.n3 55.015
R264 SLEEP.n7 SLEEP.n6 28.481
R265 SLEEP.n3 SLEEP.n2 26.386
R266 SLEEP.n3 SLEEP.n1 23.92
R267 SLEEP.n8 SLEEP.n5 21.76
R268 SLEEP.n11 SLEEP.n8 21.76
R269 SLEEP.n14 SLEEP.n11 21.76
R270 SLEEP.n17 SLEEP.n14 21.76
R271 SLEEP.n19 SLEEP.n18 18.257
R272 SLEEP.n10 SLEEP.n9 16.796
R273 SLEEP SLEEP.n17 7.68
R274 SLEEP.n16 SLEEP.n15 6.572
R275 SLEEP.n13 SLEEP.n12 5.112
R276 A.n0 A.t3 212.079
R277 A.n2 A.t1 212.079
R278 A.n0 A.t2 174.833
R279 A.n1 A.t0 139.779
R280 A A.n2 112.471
R281 A.n2 A.n1 35.054
R282 A.n1 A.n0 26.29
C0 VPB SLEEP 0.11fF
C1 X VGND 1.79fF
C2 A VGND 0.18fF
C3 SLEEP X 1.01fF
C4 VPB VPWR 0.17fF
C5 VPWR VGND 0.19fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__lpflow_isobufsrc_16.ext - technology: sky130A

.subckt sky130_fd_sc_hd__lpflow_isobufsrc_16 A X SLEEP VGND VPWR VNB VPB
X0 VPWR.t19 a_143_297.t8 a_505_297.t31 VPB.t35 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 X.t47 SLEEP.t0 a_505_297.t13 VPB.t17 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 X.t10 a_143_297.t9 VGND.t18 VNB sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 X.t9 a_143_297.t10 VGND.t17 VNB sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 X.t46 SLEEP.t1 a_505_297.t14 VPB.t18 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 X.t8 a_143_297.t11 VGND.t16 VNB sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 X.t7 a_143_297.t12 VGND.t15 VNB sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 a_505_297.t15 SLEEP.t2 X.t45 VPB.t19 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 a_505_297.t30 a_143_297.t13 VPWR.t18 VPB.t34 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 a_505_297.t29 a_143_297.t14 VPWR.t17 VPB.t33 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 a_143_297.t7 A.t0 VGND.t35 VNB sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 VGND.t34 SLEEP.t3 X.t31 VNB sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 X.t44 SLEEP.t4 a_505_297.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13 a_143_297.t0 A.t1 VGND.t0 VNB sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14 a_505_297.t28 a_143_297.t15 VPWR.t16 VPB.t32 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 VPWR.t15 a_143_297.t16 a_505_297.t27 VPB.t31 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16 X.t43 SLEEP.t5 a_505_297.t1 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17 VGND.t33 SLEEP.t6 X.t30 VNB sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X18 VGND.t32 SLEEP.t7 X.t29 VNB sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X19 VPWR.t0 A.t2 a_143_297.t1 VPB.t13 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X20 VPWR.t14 a_143_297.t17 a_505_297.t26 VPB.t30 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X21 VGND.t14 a_143_297.t18 X.t6 VNB sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X22 VGND.t13 a_143_297.t19 X.t5 VNB sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X23 VGND.t31 SLEEP.t8 X.t28 VNB sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X24 a_143_297.t2 A.t3 VPWR.t1 VPB.t14 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X25 a_505_297.t2 SLEEP.t9 X.t42 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X26 VGND.t30 SLEEP.t10 X.t27 VNB sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X27 VPWR.t13 a_143_297.t20 a_505_297.t25 VPB.t29 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X28 a_505_297.t24 a_143_297.t21 VPWR.t12 VPB.t28 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X29 a_505_297.t3 SLEEP.t11 X.t41 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X30 VGND.t12 a_143_297.t22 X.t4 VNB sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X31 X.t40 SLEEP.t12 a_505_297.t4 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X32 VGND.t11 a_143_297.t23 X.t3 VNB sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X33 X.t39 SLEEP.t13 a_505_297.t5 VPB.t5 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X34 VGND.t10 a_143_297.t24 X.t2 VNB sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X35 VPWR.t2 A.t4 a_143_297.t3 VPB.t15 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X36 VPWR.t11 a_143_297.t25 a_505_297.t23 VPB.t27 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X37 a_505_297.t6 SLEEP.t14 X.t38 VPB.t6 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X38 VGND.t1 A.t5 a_143_297.t4 VNB sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X39 a_505_297.t7 SLEEP.t15 X.t37 VPB.t7 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X40 X.t26 SLEEP.t16 VGND.t29 VNB sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X41 a_505_297.t22 a_143_297.t26 VPWR.t10 VPB.t26 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X42 X.t36 SLEEP.t17 a_505_297.t8 VPB.t8 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X43 X.t1 a_143_297.t27 VGND.t9 VNB sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X44 X.t25 SLEEP.t18 VGND.t28 VNB sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X45 X.t24 SLEEP.t19 VGND.t27 VNB sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X46 X.t35 SLEEP.t20 a_505_297.t9 VPB.t9 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X47 X.t0 a_143_297.t28 VGND.t8 VNB sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X48 X.t23 SLEEP.t21 VGND.t26 VNB sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X49 X.t15 a_143_297.t29 VGND.t7 VNB sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X50 X.t22 SLEEP.t22 VGND.t25 VNB sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X51 a_505_297.t21 a_143_297.t30 VPWR.t9 VPB.t25 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X52 a_505_297.t10 SLEEP.t23 X.t34 VPB.t10 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X53 a_143_297.t5 A.t6 VPWR.t3 VPB.t16 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X54 a_505_297.t11 SLEEP.t24 X.t33 VPB.t11 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X55 VPWR.t8 a_143_297.t31 a_505_297.t20 VPB.t24 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X56 VGND.t6 a_143_297.t32 X.t14 VNB sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X57 VGND.t5 a_143_297.t33 X.t13 VNB sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X58 VGND.t24 SLEEP.t25 X.t21 VNB sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X59 a_505_297.t19 a_143_297.t34 VPWR.t7 VPB.t23 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X60 VPWR.t6 a_143_297.t35 a_505_297.t18 VPB.t22 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X61 a_505_297.t12 SLEEP.t26 X.t32 VPB.t12 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X62 VGND.t4 a_143_297.t36 X.t12 VNB sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X63 VGND.t23 SLEEP.t27 X.t20 VNB sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X64 X.t19 SLEEP.t28 VGND.t22 VNB sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X65 VPWR.t5 a_143_297.t37 a_505_297.t17 VPB.t21 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X66 VGND.t2 A.t7 a_143_297.t6 VNB sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X67 VGND.t21 SLEEP.t29 X.t18 VNB sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X68 a_505_297.t16 a_143_297.t38 VPWR.t4 VPB.t20 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X69 X.t17 SLEEP.t30 VGND.t20 VNB sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X70 X.t11 a_143_297.t39 VGND.t3 VNB sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X71 X.t16 SLEEP.t31 VGND.t19 VNB sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
R0 a_143_297.n1 a_143_297.t14 212.079
R1 a_143_297.n3 a_143_297.t17 212.079
R2 a_143_297.n6 a_143_297.t21 212.079
R3 a_143_297.n11 a_143_297.t25 212.079
R4 a_143_297.n14 a_143_297.t26 212.079
R5 a_143_297.n17 a_143_297.t35 212.079
R6 a_143_297.n20 a_143_297.t38 212.079
R7 a_143_297.n25 a_143_297.t8 212.079
R8 a_143_297.n28 a_143_297.t13 212.079
R9 a_143_297.n31 a_143_297.t16 212.079
R10 a_143_297.n34 a_143_297.t15 212.079
R11 a_143_297.n39 a_143_297.t20 212.079
R12 a_143_297.n42 a_143_297.t30 212.079
R13 a_143_297.n45 a_143_297.t31 212.079
R14 a_143_297.n48 a_143_297.t34 212.079
R15 a_143_297.n51 a_143_297.t37 212.079
R16 a_143_297.n1 a_143_297.t24 139.779
R17 a_143_297.n3 a_143_297.t29 139.779
R18 a_143_297.n6 a_143_297.t23 139.779
R19 a_143_297.n11 a_143_297.t28 139.779
R20 a_143_297.n14 a_143_297.t22 139.779
R21 a_143_297.n17 a_143_297.t11 139.779
R22 a_143_297.n20 a_143_297.t19 139.779
R23 a_143_297.n25 a_143_297.t10 139.779
R24 a_143_297.n28 a_143_297.t18 139.779
R25 a_143_297.n31 a_143_297.t39 139.779
R26 a_143_297.n34 a_143_297.t36 139.779
R27 a_143_297.n39 a_143_297.t12 139.779
R28 a_143_297.n42 a_143_297.t33 139.779
R29 a_143_297.n45 a_143_297.t9 139.779
R30 a_143_297.n48 a_143_297.t32 139.779
R31 a_143_297.n51 a_143_297.t27 139.779
R32 a_143_297.n57 a_143_297.n56 133.913
R33 a_143_297.n59 a_143_297.n58 117.525
R34 a_143_297.n5 a_143_297.n2 96.723
R35 a_143_297.n53 a_143_297.n52 76
R36 a_143_297.n5 a_143_297.n4 76
R37 a_143_297.n8 a_143_297.n7 76
R38 a_143_297.n10 a_143_297.n9 76
R39 a_143_297.n13 a_143_297.n12 76
R40 a_143_297.n16 a_143_297.n15 76
R41 a_143_297.n19 a_143_297.n18 76
R42 a_143_297.n22 a_143_297.n21 76
R43 a_143_297.n24 a_143_297.n23 76
R44 a_143_297.n27 a_143_297.n26 76
R45 a_143_297.n30 a_143_297.n29 76
R46 a_143_297.n33 a_143_297.n32 76
R47 a_143_297.n36 a_143_297.n35 76
R48 a_143_297.n38 a_143_297.n37 76
R49 a_143_297.n41 a_143_297.n40 76
R50 a_143_297.n44 a_143_297.n43 76
R51 a_143_297.n47 a_143_297.n46 76
R52 a_143_297.n50 a_143_297.n49 76
R53 a_143_297.n57 a_143_297.n55 69.5
R54 a_143_297.n54 a_143_297.n0 65.845
R55 a_143_297.n54 a_143_297.n53 64.262
R56 a_143_297.n58 a_143_297.n57 34.909
R57 a_143_297.n40 a_143_297.n39 33.593
R58 a_143_297.n26 a_143_297.n25 30.672
R59 a_143_297.n12 a_143_297.n11 27.751
R60 a_143_297.n56 a_143_297.t3 26.595
R61 a_143_297.n56 a_143_297.t5 26.595
R62 a_143_297.t1 a_143_297.n59 26.595
R63 a_143_297.n59 a_143_297.t2 26.595
R64 a_143_297.n55 a_143_297.t6 24.923
R65 a_143_297.n55 a_143_297.t7 24.923
R66 a_143_297.n0 a_143_297.t4 24.923
R67 a_143_297.n0 a_143_297.t0 24.923
R68 a_143_297.n43 a_143_297.n42 21.909
R69 a_143_297.n8 a_143_297.n5 20.723
R70 a_143_297.n10 a_143_297.n8 20.723
R71 a_143_297.n13 a_143_297.n10 20.723
R72 a_143_297.n16 a_143_297.n13 20.723
R73 a_143_297.n19 a_143_297.n16 20.723
R74 a_143_297.n22 a_143_297.n19 20.723
R75 a_143_297.n24 a_143_297.n22 20.723
R76 a_143_297.n27 a_143_297.n24 20.723
R77 a_143_297.n30 a_143_297.n27 20.723
R78 a_143_297.n33 a_143_297.n30 20.723
R79 a_143_297.n36 a_143_297.n33 20.723
R80 a_143_297.n38 a_143_297.n36 20.723
R81 a_143_297.n41 a_143_297.n38 20.723
R82 a_143_297.n44 a_143_297.n41 20.723
R83 a_143_297.n47 a_143_297.n44 20.723
R84 a_143_297.n50 a_143_297.n47 20.723
R85 a_143_297.n53 a_143_297.n50 20.723
R86 a_143_297.n29 a_143_297.n28 18.987
R87 a_143_297.n15 a_143_297.n14 16.066
R88 a_143_297.n2 a_143_297.n1 13.145
R89 a_143_297.n52 a_143_297.n51 13.145
R90 a_143_297.n58 a_143_297.n54 12.8
R91 a_143_297.n7 a_143_297.n6 10.224
R92 a_143_297.n46 a_143_297.n45 10.224
R93 a_143_297.n21 a_143_297.n20 7.303
R94 a_143_297.n32 a_143_297.n31 7.303
R95 a_143_297.n18 a_143_297.n17 4.381
R96 a_143_297.n35 a_143_297.n34 4.381
R97 a_143_297.n4 a_143_297.n3 1.46
R98 a_143_297.n49 a_143_297.n48 1.46
R99 a_505_297.n19 a_505_297.t6 225.591
R100 a_505_297.n2 a_505_297.t17 169.699
R101 a_505_297.n19 a_505_297.n18 154.573
R102 a_505_297.n21 a_505_297.n20 154.573
R103 a_505_297.n23 a_505_297.n22 154.573
R104 a_505_297.n25 a_505_297.n24 154.573
R105 a_505_297.n27 a_505_297.n26 154.573
R106 a_505_297.n17 a_505_297.n16 154.573
R107 a_505_297.n29 a_505_297.n28 154.572
R108 a_505_297.n2 a_505_297.n1 109.736
R109 a_505_297.n4 a_505_297.n3 109.736
R110 a_505_297.n6 a_505_297.n5 109.736
R111 a_505_297.n8 a_505_297.n7 109.736
R112 a_505_297.n10 a_505_297.n9 109.736
R113 a_505_297.n12 a_505_297.n11 109.736
R114 a_505_297.n14 a_505_297.n13 109.736
R115 a_505_297.n15 a_505_297.n0 90.234
R116 a_505_297.n17 a_505_297.n15 64.95
R117 a_505_297.n15 a_505_297.n14 55.464
R118 a_505_297.n21 a_505_297.n19 44.423
R119 a_505_297.n23 a_505_297.n21 44.423
R120 a_505_297.n25 a_505_297.n23 44.423
R121 a_505_297.n27 a_505_297.n25 44.423
R122 a_505_297.n28 a_505_297.n17 44.423
R123 a_505_297.n28 a_505_297.n27 44.423
R124 a_505_297.n4 a_505_297.n2 35.961
R125 a_505_297.n6 a_505_297.n4 35.961
R126 a_505_297.n8 a_505_297.n6 35.961
R127 a_505_297.n10 a_505_297.n8 35.961
R128 a_505_297.n12 a_505_297.n10 35.961
R129 a_505_297.n14 a_505_297.n12 35.961
R130 a_505_297.n18 a_505_297.t8 26.595
R131 a_505_297.n18 a_505_297.t12 26.595
R132 a_505_297.n20 a_505_297.t1 26.595
R133 a_505_297.n20 a_505_297.t3 26.595
R134 a_505_297.n22 a_505_297.t5 26.595
R135 a_505_297.n22 a_505_297.t7 26.595
R136 a_505_297.n24 a_505_297.t9 26.595
R137 a_505_297.n24 a_505_297.t10 26.595
R138 a_505_297.n26 a_505_297.t13 26.595
R139 a_505_297.n26 a_505_297.t15 26.595
R140 a_505_297.n0 a_505_297.t14 26.595
R141 a_505_297.n0 a_505_297.t29 26.595
R142 a_505_297.n1 a_505_297.t20 26.595
R143 a_505_297.n1 a_505_297.t19 26.595
R144 a_505_297.n3 a_505_297.t25 26.595
R145 a_505_297.n3 a_505_297.t21 26.595
R146 a_505_297.n5 a_505_297.t27 26.595
R147 a_505_297.n5 a_505_297.t28 26.595
R148 a_505_297.n7 a_505_297.t31 26.595
R149 a_505_297.n7 a_505_297.t30 26.595
R150 a_505_297.n9 a_505_297.t18 26.595
R151 a_505_297.n9 a_505_297.t16 26.595
R152 a_505_297.n11 a_505_297.t23 26.595
R153 a_505_297.n11 a_505_297.t22 26.595
R154 a_505_297.n13 a_505_297.t26 26.595
R155 a_505_297.n13 a_505_297.t24 26.595
R156 a_505_297.n16 a_505_297.t4 26.595
R157 a_505_297.n16 a_505_297.t11 26.595
R158 a_505_297.t0 a_505_297.n29 26.595
R159 a_505_297.n29 a_505_297.t2 26.595
R160 VPWR.n3 VPWR.n0 173.557
R161 VPWR.n33 VPWR.n32 169.933
R162 VPWR.n28 VPWR.n27 169.933
R163 VPWR.n23 VPWR.n22 169.933
R164 VPWR.n17 VPWR.n16 169.933
R165 VPWR.n11 VPWR.n10 169.933
R166 VPWR.n7 VPWR.n6 169.933
R167 VPWR.n2 VPWR.n1 169.933
R168 VPWR.n47 VPWR.t3 157.283
R169 VPWR.n37 VPWR.t0 153.549
R170 VPWR.n42 VPWR.n41 133.221
R171 VPWR.n41 VPWR.t1 26.595
R172 VPWR.n41 VPWR.t2 26.595
R173 VPWR.n32 VPWR.t7 26.595
R174 VPWR.n32 VPWR.t5 26.595
R175 VPWR.n27 VPWR.t9 26.595
R176 VPWR.n27 VPWR.t8 26.595
R177 VPWR.n22 VPWR.t16 26.595
R178 VPWR.n22 VPWR.t13 26.595
R179 VPWR.n16 VPWR.t18 26.595
R180 VPWR.n16 VPWR.t15 26.595
R181 VPWR.n10 VPWR.t4 26.595
R182 VPWR.n10 VPWR.t19 26.595
R183 VPWR.n6 VPWR.t10 26.595
R184 VPWR.n6 VPWR.t6 26.595
R185 VPWR.n1 VPWR.t12 26.595
R186 VPWR.n1 VPWR.t11 26.595
R187 VPWR.n0 VPWR.t17 26.595
R188 VPWR.n0 VPWR.t14 26.595
R189 VPWR.n48 VPWR.n47 9.92
R190 VPWR.n43 VPWR.n42 9.035
R191 VPWR.n12 VPWR.n11 7.152
R192 VPWR.n5 VPWR.n4 4.65
R193 VPWR.n9 VPWR.n8 4.65
R194 VPWR.n13 VPWR.n12 4.65
R195 VPWR.n15 VPWR.n14 4.65
R196 VPWR.n19 VPWR.n18 4.65
R197 VPWR.n21 VPWR.n20 4.65
R198 VPWR.n24 VPWR.n23 4.65
R199 VPWR.n26 VPWR.n25 4.65
R200 VPWR.n29 VPWR.n28 4.65
R201 VPWR.n31 VPWR.n30 4.65
R202 VPWR.n34 VPWR.n33 4.65
R203 VPWR.n36 VPWR.n35 4.65
R204 VPWR.n38 VPWR.n37 4.65
R205 VPWR.n40 VPWR.n39 4.65
R206 VPWR.n44 VPWR.n43 4.65
R207 VPWR.n46 VPWR.n45 4.65
R208 VPWR.n3 VPWR.n2 3.764
R209 VPWR.n8 VPWR.n7 2.635
R210 VPWR.n18 VPWR.n17 1.129
R211 VPWR.n5 VPWR.n3 0.233
R212 VPWR.n9 VPWR.n5 0.119
R213 VPWR.n13 VPWR.n9 0.119
R214 VPWR.n15 VPWR.n13 0.119
R215 VPWR.n19 VPWR.n15 0.119
R216 VPWR.n21 VPWR.n19 0.119
R217 VPWR.n24 VPWR.n21 0.119
R218 VPWR.n26 VPWR.n24 0.119
R219 VPWR.n29 VPWR.n26 0.119
R220 VPWR.n31 VPWR.n29 0.119
R221 VPWR.n34 VPWR.n31 0.119
R222 VPWR.n36 VPWR.n34 0.119
R223 VPWR.n38 VPWR.n36 0.119
R224 VPWR.n40 VPWR.n38 0.119
R225 VPWR.n44 VPWR.n40 0.119
R226 VPWR.n46 VPWR.n44 0.119
R227 VPWR.n48 VPWR.n46 0.119
R228 VPWR VPWR.n48 0.022
R229 VPB.t13 VPB.t21 580.062
R230 VPB VPB.t16 292.99
R231 VPB.t8 VPB.t6 248.598
R232 VPB.t12 VPB.t8 248.598
R233 VPB.t1 VPB.t12 248.598
R234 VPB.t3 VPB.t1 248.598
R235 VPB.t5 VPB.t3 248.598
R236 VPB.t7 VPB.t5 248.598
R237 VPB.t9 VPB.t7 248.598
R238 VPB.t10 VPB.t9 248.598
R239 VPB.t17 VPB.t10 248.598
R240 VPB.t19 VPB.t17 248.598
R241 VPB.t0 VPB.t19 248.598
R242 VPB.t2 VPB.t0 248.598
R243 VPB.t4 VPB.t2 248.598
R244 VPB.t11 VPB.t4 248.598
R245 VPB.t18 VPB.t11 248.598
R246 VPB.t33 VPB.t18 248.598
R247 VPB.t30 VPB.t33 248.598
R248 VPB.t28 VPB.t30 248.598
R249 VPB.t27 VPB.t28 248.598
R250 VPB.t26 VPB.t27 248.598
R251 VPB.t22 VPB.t26 248.598
R252 VPB.t20 VPB.t22 248.598
R253 VPB.t35 VPB.t20 248.598
R254 VPB.t34 VPB.t35 248.598
R255 VPB.t31 VPB.t34 248.598
R256 VPB.t32 VPB.t31 248.598
R257 VPB.t29 VPB.t32 248.598
R258 VPB.t25 VPB.t29 248.598
R259 VPB.t24 VPB.t25 248.598
R260 VPB.t23 VPB.t24 248.598
R261 VPB.t21 VPB.t23 248.598
R262 VPB.t14 VPB.t13 248.598
R263 VPB.t15 VPB.t14 248.598
R264 VPB.t16 VPB.t15 248.598
R265 SLEEP.n0 SLEEP.t14 212.079
R266 SLEEP.n1 SLEEP.t17 212.079
R267 SLEEP.n2 SLEEP.t26 212.079
R268 SLEEP.n6 SLEEP.t5 212.079
R269 SLEEP.n9 SLEEP.t11 212.079
R270 SLEEP.n12 SLEEP.t13 212.079
R271 SLEEP.n15 SLEEP.t15 212.079
R272 SLEEP.n20 SLEEP.t20 212.079
R273 SLEEP.n45 SLEEP.t23 212.079
R274 SLEEP.n42 SLEEP.t0 212.079
R275 SLEEP.n39 SLEEP.t2 212.079
R276 SLEEP.n36 SLEEP.t4 212.079
R277 SLEEP.n33 SLEEP.t9 212.079
R278 SLEEP.n28 SLEEP.t12 212.079
R279 SLEEP.n25 SLEEP.t24 212.079
R280 SLEEP.n23 SLEEP.t1 212.079
R281 SLEEP.n0 SLEEP.t3 139.779
R282 SLEEP.n1 SLEEP.t28 139.779
R283 SLEEP.n2 SLEEP.t27 139.779
R284 SLEEP.n6 SLEEP.t21 139.779
R285 SLEEP.n9 SLEEP.t25 139.779
R286 SLEEP.n12 SLEEP.t19 139.779
R287 SLEEP.n15 SLEEP.t10 139.779
R288 SLEEP.n20 SLEEP.t18 139.779
R289 SLEEP.n45 SLEEP.t8 139.779
R290 SLEEP.n42 SLEEP.t16 139.779
R291 SLEEP.n39 SLEEP.t7 139.779
R292 SLEEP.n36 SLEEP.t31 139.779
R293 SLEEP.n33 SLEEP.t6 139.779
R294 SLEEP.n28 SLEEP.t30 139.779
R295 SLEEP.n25 SLEEP.t29 139.779
R296 SLEEP.n23 SLEEP.t22 139.779
R297 SLEEP.n27 SLEEP.n24 96.723
R298 SLEEP.n5 SLEEP.n4 76
R299 SLEEP.n8 SLEEP.n7 76
R300 SLEEP.n11 SLEEP.n10 76
R301 SLEEP.n14 SLEEP.n13 76
R302 SLEEP.n17 SLEEP.n16 76
R303 SLEEP.n19 SLEEP.n18 76
R304 SLEEP.n22 SLEEP.n21 76
R305 SLEEP.n47 SLEEP.n46 76
R306 SLEEP.n44 SLEEP.n43 76
R307 SLEEP.n41 SLEEP.n40 76
R308 SLEEP.n38 SLEEP.n37 76
R309 SLEEP.n35 SLEEP.n34 76
R310 SLEEP.n32 SLEEP.n31 76
R311 SLEEP.n30 SLEEP.n29 76
R312 SLEEP.n27 SLEEP.n26 76
R313 SLEEP.n1 SLEEP.n0 61.345
R314 SLEEP.n5 SLEEP.n3 53.779
R315 SLEEP.n21 SLEEP.n20 30.672
R316 SLEEP.n7 SLEEP.n6 27.751
R317 SLEEP.n34 SLEEP.n33 27.751
R318 SLEEP.n3 SLEEP.n2 27.196
R319 SLEEP.n3 SLEEP.n1 23.06
R320 SLEEP.n8 SLEEP.n5 20.723
R321 SLEEP.n11 SLEEP.n8 20.723
R322 SLEEP.n14 SLEEP.n11 20.723
R323 SLEEP.n17 SLEEP.n14 20.723
R324 SLEEP.n19 SLEEP.n17 20.723
R325 SLEEP.n22 SLEEP.n19 20.723
R326 SLEEP.n47 SLEEP.n44 20.723
R327 SLEEP.n44 SLEEP.n41 20.723
R328 SLEEP.n41 SLEEP.n38 20.723
R329 SLEEP.n38 SLEEP.n35 20.723
R330 SLEEP.n35 SLEEP.n32 20.723
R331 SLEEP.n32 SLEEP.n30 20.723
R332 SLEEP.n30 SLEEP.n27 20.723
R333 SLEEP.n46 SLEEP.n45 18.987
R334 SLEEP.n10 SLEEP.n9 16.066
R335 SLEEP.n37 SLEEP.n36 16.066
R336 SLEEP SLEEP.n22 15.542
R337 SLEEP.n24 SLEEP.n23 13.145
R338 SLEEP.n29 SLEEP.n28 10.224
R339 SLEEP.n16 SLEEP.n15 7.303
R340 SLEEP.n43 SLEEP.n42 7.303
R341 SLEEP SLEEP.n47 5.18
R342 SLEEP.n13 SLEEP.n12 4.381
R343 SLEEP.n40 SLEEP.n39 4.381
R344 SLEEP.n26 SLEEP.n25 1.46
R345 X.n2 X.n0 198.996
R346 X.n2 X.n1 154.573
R347 X.n4 X.n3 154.573
R348 X.n6 X.n5 154.573
R349 X.n8 X.n7 154.573
R350 X.n10 X.n9 154.573
R351 X.n12 X.n11 154.573
R352 X.n14 X.n13 154.573
R353 X.n17 X.n15 88.89
R354 X.n45 X.n44 52.64
R355 X.n17 X.n16 52.624
R356 X.n19 X.n18 52.624
R357 X.n21 X.n20 52.624
R358 X.n23 X.n22 52.624
R359 X.n25 X.n24 52.624
R360 X.n27 X.n26 52.624
R361 X.n29 X.n28 52.624
R362 X.n31 X.n30 52.624
R363 X.n33 X.n32 52.624
R364 X.n35 X.n34 52.624
R365 X.n37 X.n36 52.624
R366 X.n39 X.n38 52.624
R367 X.n41 X.n40 52.624
R368 X.n43 X.n42 52.624
R369 X.n4 X.n2 44.423
R370 X.n6 X.n4 44.423
R371 X.n8 X.n6 44.423
R372 X.n10 X.n8 44.423
R373 X.n12 X.n10 44.423
R374 X.n14 X.n12 44.423
R375 X.n19 X.n17 36.266
R376 X.n21 X.n19 36.266
R377 X.n23 X.n21 36.266
R378 X.n25 X.n23 36.266
R379 X.n27 X.n25 36.266
R380 X.n29 X.n27 36.266
R381 X.n31 X.n29 36.266
R382 X.n33 X.n31 36.266
R383 X.n35 X.n33 36.266
R384 X.n37 X.n35 36.266
R385 X.n39 X.n37 36.266
R386 X.n41 X.n39 36.266
R387 X.n43 X.n41 36.266
R388 X.n45 X.n43 36.266
R389 X.n0 X.t33 26.595
R390 X.n0 X.t46 26.595
R391 X.n1 X.t42 26.595
R392 X.n1 X.t40 26.595
R393 X.n3 X.t45 26.595
R394 X.n3 X.t44 26.595
R395 X.n5 X.t34 26.595
R396 X.n5 X.t47 26.595
R397 X.n7 X.t37 26.595
R398 X.n7 X.t35 26.595
R399 X.n9 X.t41 26.595
R400 X.n9 X.t39 26.595
R401 X.n11 X.t32 26.595
R402 X.n11 X.t43 26.595
R403 X.n13 X.t38 26.595
R404 X.n13 X.t36 26.595
R405 X.n15 X.t14 24.923
R406 X.n15 X.t1 24.923
R407 X.n16 X.t13 24.923
R408 X.n16 X.t10 24.923
R409 X.n18 X.t12 24.923
R410 X.n18 X.t7 24.923
R411 X.n20 X.t6 24.923
R412 X.n20 X.t11 24.923
R413 X.n22 X.t5 24.923
R414 X.n22 X.t9 24.923
R415 X.n24 X.t4 24.923
R416 X.n24 X.t8 24.923
R417 X.n26 X.t3 24.923
R418 X.n26 X.t0 24.923
R419 X.n28 X.t2 24.923
R420 X.n28 X.t15 24.923
R421 X.n30 X.t18 24.923
R422 X.n30 X.t22 24.923
R423 X.n32 X.t30 24.923
R424 X.n32 X.t17 24.923
R425 X.n34 X.t29 24.923
R426 X.n34 X.t16 24.923
R427 X.n36 X.t28 24.923
R428 X.n36 X.t26 24.923
R429 X.n38 X.t27 24.923
R430 X.n38 X.t25 24.923
R431 X.n40 X.t21 24.923
R432 X.n40 X.t24 24.923
R433 X.n42 X.t20 24.923
R434 X.n42 X.t23 24.923
R435 X.n44 X.t31 24.923
R436 X.n44 X.t19 24.923
R437 X X.n45 12.311
R438 X X.n14 2.232
R439 VGND.n2 VGND.t34 194.438
R440 VGND.n1 VGND.n0 115.464
R441 VGND.n6 VGND.n5 115.464
R442 VGND.n12 VGND.n11 115.464
R443 VGND.n18 VGND.n17 115.464
R444 VGND.n24 VGND.n23 115.464
R445 VGND.n28 VGND.n27 115.464
R446 VGND.n34 VGND.n33 115.464
R447 VGND.n40 VGND.n39 115.464
R448 VGND.n46 VGND.n45 115.464
R449 VGND.n52 VGND.n51 115.464
R450 VGND.n58 VGND.n57 115.464
R451 VGND.n62 VGND.n61 115.464
R452 VGND.n68 VGND.n67 115.464
R453 VGND.n74 VGND.n73 115.464
R454 VGND.n80 VGND.n79 115.464
R455 VGND.n95 VGND.t35 103.783
R456 VGND.n91 VGND.n90 70.197
R457 VGND.n85 VGND.t9 56.307
R458 VGND.n85 VGND.t1 56.307
R459 VGND.n0 VGND.t22 24.923
R460 VGND.n0 VGND.t23 24.923
R461 VGND.n5 VGND.t26 24.923
R462 VGND.n5 VGND.t24 24.923
R463 VGND.n11 VGND.t27 24.923
R464 VGND.n11 VGND.t30 24.923
R465 VGND.n17 VGND.t28 24.923
R466 VGND.n17 VGND.t31 24.923
R467 VGND.n23 VGND.t29 24.923
R468 VGND.n23 VGND.t32 24.923
R469 VGND.n27 VGND.t19 24.923
R470 VGND.n27 VGND.t33 24.923
R471 VGND.n33 VGND.t20 24.923
R472 VGND.n33 VGND.t21 24.923
R473 VGND.n39 VGND.t25 24.923
R474 VGND.n39 VGND.t10 24.923
R475 VGND.n45 VGND.t7 24.923
R476 VGND.n45 VGND.t11 24.923
R477 VGND.n51 VGND.t8 24.923
R478 VGND.n51 VGND.t12 24.923
R479 VGND.n57 VGND.t16 24.923
R480 VGND.n57 VGND.t13 24.923
R481 VGND.n61 VGND.t17 24.923
R482 VGND.n61 VGND.t14 24.923
R483 VGND.n67 VGND.t3 24.923
R484 VGND.n67 VGND.t4 24.923
R485 VGND.n73 VGND.t15 24.923
R486 VGND.n73 VGND.t5 24.923
R487 VGND.n79 VGND.t18 24.923
R488 VGND.n79 VGND.t6 24.923
R489 VGND.n90 VGND.t0 24.923
R490 VGND.n90 VGND.t2 24.923
R491 VGND.n29 VGND.n28 15.058
R492 VGND.n59 VGND.n58 15.058
R493 VGND.n2 VGND.n1 14.521
R494 VGND.n25 VGND.n24 13.552
R495 VGND.n63 VGND.n62 13.552
R496 VGND.n86 VGND.n85 13.032
R497 VGND.n35 VGND.n34 9.035
R498 VGND.n53 VGND.n52 9.035
R499 VGND.n19 VGND.n18 7.529
R500 VGND.n69 VGND.n68 7.529
R501 VGND.n4 VGND.n3 4.65
R502 VGND.n8 VGND.n7 4.65
R503 VGND.n10 VGND.n9 4.65
R504 VGND.n14 VGND.n13 4.65
R505 VGND.n16 VGND.n15 4.65
R506 VGND.n20 VGND.n19 4.65
R507 VGND.n22 VGND.n21 4.65
R508 VGND.n26 VGND.n25 4.65
R509 VGND.n30 VGND.n29 4.65
R510 VGND.n32 VGND.n31 4.65
R511 VGND.n36 VGND.n35 4.65
R512 VGND.n38 VGND.n37 4.65
R513 VGND.n42 VGND.n41 4.65
R514 VGND.n44 VGND.n43 4.65
R515 VGND.n48 VGND.n47 4.65
R516 VGND.n50 VGND.n49 4.65
R517 VGND.n54 VGND.n53 4.65
R518 VGND.n56 VGND.n55 4.65
R519 VGND.n60 VGND.n59 4.65
R520 VGND.n64 VGND.n63 4.65
R521 VGND.n66 VGND.n65 4.65
R522 VGND.n70 VGND.n69 4.65
R523 VGND.n72 VGND.n71 4.65
R524 VGND.n76 VGND.n75 4.65
R525 VGND.n78 VGND.n77 4.65
R526 VGND.n82 VGND.n81 4.65
R527 VGND.n84 VGND.n83 4.65
R528 VGND.n87 VGND.n86 4.65
R529 VGND.n89 VGND.n88 4.65
R530 VGND.n92 VGND.n91 4.65
R531 VGND.n94 VGND.n93 4.65
R532 VGND.n7 VGND.n6 4.517
R533 VGND.n81 VGND.n80 4.517
R534 VGND.n96 VGND.n95 3.876
R535 VGND.n41 VGND.n40 3.011
R536 VGND.n47 VGND.n46 3.011
R537 VGND.n13 VGND.n12 1.505
R538 VGND.n75 VGND.n74 1.505
R539 VGND.n4 VGND.n2 0.289
R540 VGND.n96 VGND.n94 0.139
R541 VGND VGND.n96 0.122
R542 VGND.n8 VGND.n4 0.119
R543 VGND.n10 VGND.n8 0.119
R544 VGND.n14 VGND.n10 0.119
R545 VGND.n16 VGND.n14 0.119
R546 VGND.n20 VGND.n16 0.119
R547 VGND.n22 VGND.n20 0.119
R548 VGND.n26 VGND.n22 0.119
R549 VGND.n30 VGND.n26 0.119
R550 VGND.n32 VGND.n30 0.119
R551 VGND.n36 VGND.n32 0.119
R552 VGND.n38 VGND.n36 0.119
R553 VGND.n42 VGND.n38 0.119
R554 VGND.n44 VGND.n42 0.119
R555 VGND.n48 VGND.n44 0.119
R556 VGND.n50 VGND.n48 0.119
R557 VGND.n54 VGND.n50 0.119
R558 VGND.n56 VGND.n54 0.119
R559 VGND.n60 VGND.n56 0.119
R560 VGND.n64 VGND.n60 0.119
R561 VGND.n66 VGND.n64 0.119
R562 VGND.n70 VGND.n66 0.119
R563 VGND.n72 VGND.n70 0.119
R564 VGND.n76 VGND.n72 0.119
R565 VGND.n78 VGND.n76 0.119
R566 VGND.n82 VGND.n78 0.119
R567 VGND.n84 VGND.n82 0.119
R568 VGND.n87 VGND.n84 0.119
R569 VGND.n89 VGND.n87 0.119
R570 VGND.n92 VGND.n89 0.119
R571 VGND.n94 VGND.n92 0.119
R572 A.n0 A.t2 212.079
R573 A.n2 A.t3 212.079
R574 A.n4 A.t4 212.079
R575 A.n6 A.t6 212.079
R576 A.n0 A.t5 171.912
R577 A.n5 A.t0 139.779
R578 A.n3 A.t7 139.779
R579 A.n1 A.t1 139.779
R580 A A.n6 60.544
R581 A.n2 A.n1 32.133
R582 A.n4 A.n3 32.133
R583 A.n6 A.n5 32.133
R584 A.n1 A.n0 29.212
R585 A.n3 A.n2 29.212
R586 A.n5 A.n4 29.212
C0 VPWR VGND 0.36fF
C1 VPB SLEEP 0.22fF
C2 X VGND 3.57fF
C3 A VGND 0.20fF
C4 SLEEP X 2.22fF
C5 VPB VPWR 0.31fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__lpflow_isobufsrckapwr_16.ext - technology: sky130A

.subckt sky130_fd_sc_hd__lpflow_isobufsrckapwr_16 X A SLEEP VGND VPWR KAPWR VNB VPB
X0 VPWR.t3 SLEEP.t0 a_255_297.t5 VPB.t23 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 KAPWR.t19 a_1122_47.t8 X.t7 VPB.t10 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 VGND.t10 SLEEP.t1 a_341_47.t8 VNB.t10 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 VGND.t26 a_1122_47.t9 X.t10 VNB.t26 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 VGND.t25 a_1122_47.t10 X.t9 VNB.t25 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 a_255_297.t4 SLEEP.t2 VPWR.t2 VPB.t22 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 VGND.t24 a_1122_47.t11 X.t8 VNB.t24 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7 X.t6 a_1122_47.t12 KAPWR.t18 VPB.t11 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 a_341_47.t11 a_147_47.t2 VGND.t28 VNB.t28 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 VPWR.t1 SLEEP.t3 a_255_297.t3 VPB.t21 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 KAPWR.t1 a_341_47.t12 a_1122_47.t2 VPB.t19 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 KAPWR.t17 a_1122_47.t13 X.t5 VPB.t12 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 VGND.t23 a_1122_47.t14 X.t23 VNB.t23 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13 X.t4 a_1122_47.t15 KAPWR.t16 VPB.t13 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14 VGND.t5 a_341_47.t13 a_1122_47.t3 VNB.t5 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15 a_255_297.t6 a_147_47.t3 a_341_47.t9 VPB.t27 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16 KAPWR.t15 a_1122_47.t16 X.t3 VPB.t14 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17 X.t22 a_1122_47.t17 VGND.t22 VNB.t22 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18 VGND.t21 a_1122_47.t18 X.t21 VNB.t21 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19 X.t2 a_1122_47.t19 KAPWR.t14 VPB.t15 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X20 a_341_47.t10 a_147_47.t4 a_255_297.t7 VPB.t28 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X21 KAPWR.t13 a_1122_47.t20 X.t1 VPB.t16 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X22 X.t20 a_1122_47.t21 VGND.t20 VNB.t20 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23 a_147_47.t1 A.t0 VGND.t27 VNB.t27 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X24 VGND.t6 a_147_47.t5 a_341_47.t3 VNB.t6 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X25 VGND.t19 a_1122_47.t22 X.t19 VNB.t19 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X26 a_147_47.t0 A.t1 VPWR.t4 VPB.t26 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X27 a_255_297.t1 a_147_47.t6 a_341_47.t4 VPB.t18 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X28 a_1122_47.t4 a_341_47.t14 KAPWR.t2 VPB.t24 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X29 VGND.t0 a_147_47.t7 a_341_47.t1 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X30 X.t0 a_1122_47.t23 KAPWR.t12 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X31 KAPWR.t11 a_1122_47.t24 X.t31 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X32 VGND.t9 SLEEP.t4 a_341_47.t7 VNB.t9 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X33 X.t18 a_1122_47.t25 VGND.t18 VNB.t18 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X34 a_1122_47.t5 a_341_47.t15 VGND.t4 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X35 KAPWR.t10 a_1122_47.t26 X.t30 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X36 X.t29 a_1122_47.t27 KAPWR.t9 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X37 X.t17 a_1122_47.t28 VGND.t17 VNB.t17 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X38 X.t16 a_1122_47.t29 VGND.t16 VNB.t16 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X39 a_1122_47.t6 a_341_47.t16 VGND.t3 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X40 a_255_297.t2 SLEEP.t5 VPWR.t0 VPB.t20 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X41 KAPWR.t3 a_341_47.t17 a_1122_47.t7 VPB.t25 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X42 X.t28 a_1122_47.t30 KAPWR.t8 VPB.t5 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X43 a_341_47.t2 a_147_47.t8 VGND.t1 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X44 X.t27 a_1122_47.t31 KAPWR.t7 VPB.t6 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X45 a_341_47.t6 SLEEP.t6 VGND.t8 VNB.t8 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X46 a_341_47.t5 SLEEP.t7 VGND.t7 VNB.t7 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X47 X.t15 a_1122_47.t32 VGND.t15 VNB.t15 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X48 X.t14 a_1122_47.t33 VGND.t14 VNB.t14 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X49 a_341_47.t0 a_147_47.t9 a_255_297.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X50 VGND.t2 a_341_47.t18 a_1122_47.t0 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X51 X.t13 a_1122_47.t34 VGND.t13 VNB.t13 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X52 KAPWR.t6 a_1122_47.t35 X.t26 VPB.t7 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X53 KAPWR.t5 a_1122_47.t36 X.t25 VPB.t8 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X54 a_1122_47.t1 a_341_47.t19 KAPWR.t0 VPB.t17 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X55 VGND.t12 a_1122_47.t37 X.t12 VNB.t12 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X56 X.t24 a_1122_47.t38 KAPWR.t4 VPB.t9 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X57 VGND.t11 a_1122_47.t39 X.t11 VNB.t11 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
R0 SLEEP.n0 SLEEP.t5 212.079
R1 SLEEP.n7 SLEEP.t0 212.079
R2 SLEEP.n4 SLEEP.t2 212.079
R3 SLEEP.n2 SLEEP.t3 212.079
R4 SLEEP.n0 SLEEP.t1 139.779
R5 SLEEP.n7 SLEEP.t7 139.779
R6 SLEEP.n4 SLEEP.t4 139.779
R7 SLEEP.n2 SLEEP.t6 139.779
R8 SLEEP.n6 SLEEP.n3 97.76
R9 SLEEP SLEEP.n1 87.52
R10 SLEEP.n9 SLEEP.n8 76
R11 SLEEP.n6 SLEEP.n5 76
R12 SLEEP.n9 SLEEP.n6 21.76
R13 SLEEP.n3 SLEEP.n2 18.987
R14 SLEEP.n1 SLEEP.n0 16.066
R15 SLEEP SLEEP.n9 10.24
R16 SLEEP.n5 SLEEP.n4 7.303
R17 SLEEP.n8 SLEEP.n7 4.381
R18 a_255_297.n1 a_255_297.t2 181.085
R19 a_255_297.t0 a_255_297.n5 169.982
R20 a_255_297.n5 a_255_297.n4 150.25
R21 a_255_297.n1 a_255_297.n0 109.334
R22 a_255_297.n3 a_255_297.n2 91.601
R23 a_255_297.n3 a_255_297.n1 57.039
R24 a_255_297.n5 a_255_297.n3 53.035
R25 a_255_297.n2 a_255_297.t3 26.595
R26 a_255_297.n2 a_255_297.t6 26.595
R27 a_255_297.n0 a_255_297.t5 26.595
R28 a_255_297.n0 a_255_297.t4 26.595
R29 a_255_297.n4 a_255_297.t7 26.595
R30 a_255_297.n4 a_255_297.t1 26.595
R31 VPWR.n2 VPWR.n1 169.933
R32 VPWR.n3 VPWR.n0 167.714
R33 VPWR.n16 VPWR.t4 141.877
R34 VPWR.n1 VPWR.t2 26.595
R35 VPWR.n1 VPWR.t1 26.595
R36 VPWR.n0 VPWR.t0 26.595
R37 VPWR.n0 VPWR.t3 26.595
R38 VPWR.n5 VPWR.n4 4.65
R39 VPWR.n7 VPWR.n6 4.65
R40 VPWR.n9 VPWR.n8 4.65
R41 VPWR.n11 VPWR.n10 4.65
R42 VPWR.n13 VPWR.n12 4.65
R43 VPWR.n15 VPWR.n14 4.65
R44 VPWR.n17 VPWR.n16 4.65
R45 VPWR.n3 VPWR.n2 3.671
R46 VPWR.n5 VPWR.n3 0.255
R47 VPWR.n7 VPWR.n5 0.119
R48 VPWR.n9 VPWR.n7 0.119
R49 VPWR.n11 VPWR.n9 0.119
R50 VPWR.n13 VPWR.n11 0.119
R51 VPWR.n15 VPWR.n13 0.119
R52 VPWR.n17 VPWR.n15 0.119
R53 VPWR VPWR.n17 0.02
R54 VPB.t26 VPB.t0 574.143
R55 VPB.t20 VPB 375.856
R56 VPB VPB.t26 301.869
R57 VPB.t5 VPB.t8 254.517
R58 VPB.t16 VPB.t5 254.517
R59 VPB.t11 VPB.t16 254.517
R60 VPB.t7 VPB.t11 254.517
R61 VPB.t4 VPB.t7 254.517
R62 VPB.t3 VPB.t4 254.517
R63 VPB.t15 VPB.t3 254.517
R64 VPB.t13 VPB.t14 254.517
R65 VPB.t10 VPB.t13 254.517
R66 VPB.t6 VPB.t10 254.517
R67 VPB.t2 VPB.t6 254.517
R68 VPB.t1 VPB.t2 254.517
R69 VPB.t12 VPB.t1 254.517
R70 VPB.t9 VPB.t12 254.517
R71 VPB.t25 VPB.t9 254.517
R72 VPB.t24 VPB.t25 254.517
R73 VPB.t19 VPB.t24 254.517
R74 VPB.t17 VPB.t19 254.517
R75 VPB.t14 VPB.t15 251.557
R76 VPB.t23 VPB.t20 248.598
R77 VPB.t22 VPB.t23 248.598
R78 VPB.t21 VPB.t22 248.598
R79 VPB.t27 VPB.t21 248.598
R80 VPB.t28 VPB.t27 248.598
R81 VPB.t18 VPB.t28 248.598
R82 VPB.t0 VPB.t18 248.598
R83 VPB VPB.t17 145.015
R84 a_1122_47.n3 a_1122_47.t36 212.079
R85 a_1122_47.n4 a_1122_47.t30 212.079
R86 a_1122_47.n5 a_1122_47.t20 212.079
R87 a_1122_47.n7 a_1122_47.t12 212.079
R88 a_1122_47.n10 a_1122_47.t35 212.079
R89 a_1122_47.n13 a_1122_47.t27 212.079
R90 a_1122_47.n16 a_1122_47.t26 212.079
R91 a_1122_47.n21 a_1122_47.t19 212.079
R92 a_1122_47.n24 a_1122_47.t16 212.079
R93 a_1122_47.n27 a_1122_47.t15 212.079
R94 a_1122_47.n30 a_1122_47.t8 212.079
R95 a_1122_47.n35 a_1122_47.t31 212.079
R96 a_1122_47.n38 a_1122_47.t24 212.079
R97 a_1122_47.n41 a_1122_47.t23 212.079
R98 a_1122_47.n46 a_1122_47.t13 212.079
R99 a_1122_47.n47 a_1122_47.t38 212.079
R100 a_1122_47.n3 a_1122_47.t14 162.273
R101 a_1122_47.n4 a_1122_47.t25 162.273
R102 a_1122_47.n5 a_1122_47.t18 162.273
R103 a_1122_47.n7 a_1122_47.t29 162.273
R104 a_1122_47.n10 a_1122_47.t22 162.273
R105 a_1122_47.n13 a_1122_47.t33 162.273
R106 a_1122_47.n16 a_1122_47.t39 162.273
R107 a_1122_47.n21 a_1122_47.t34 162.273
R108 a_1122_47.n24 a_1122_47.t10 162.273
R109 a_1122_47.n27 a_1122_47.t28 162.273
R110 a_1122_47.n30 a_1122_47.t37 162.273
R111 a_1122_47.n35 a_1122_47.t32 162.273
R112 a_1122_47.n38 a_1122_47.t9 162.273
R113 a_1122_47.n41 a_1122_47.t17 162.273
R114 a_1122_47.n46 a_1122_47.t11 162.273
R115 a_1122_47.n47 a_1122_47.t21 162.273
R116 a_1122_47.n53 a_1122_47.n52 130.004
R117 a_1122_47.n51 a_1122_47.n1 128.898
R118 a_1122_47.n52 a_1122_47.n0 128.34
R119 a_1122_47.n50 a_1122_47.n2 124.756
R120 a_1122_47.n9 a_1122_47.n6 93.408
R121 a_1122_47.n49 a_1122_47.n48 76
R122 a_1122_47.n9 a_1122_47.n8 76
R123 a_1122_47.n12 a_1122_47.n11 76
R124 a_1122_47.n15 a_1122_47.n14 76
R125 a_1122_47.n18 a_1122_47.n17 76
R126 a_1122_47.n20 a_1122_47.n19 76
R127 a_1122_47.n23 a_1122_47.n22 76
R128 a_1122_47.n26 a_1122_47.n25 76
R129 a_1122_47.n29 a_1122_47.n28 76
R130 a_1122_47.n32 a_1122_47.n31 76
R131 a_1122_47.n34 a_1122_47.n33 76
R132 a_1122_47.n37 a_1122_47.n36 76
R133 a_1122_47.n40 a_1122_47.n39 76
R134 a_1122_47.n43 a_1122_47.n42 76
R135 a_1122_47.n45 a_1122_47.n44 76
R136 a_1122_47.n4 a_1122_47.n3 55.269
R137 a_1122_47.n5 a_1122_47.n4 55.269
R138 a_1122_47.n50 a_1122_47.n49 43.52
R139 a_1122_47.n52 a_1122_47.n51 43.264
R140 a_1122_47.n0 a_1122_47.t0 40
R141 a_1122_47.n0 a_1122_47.t6 40
R142 a_1122_47.n2 a_1122_47.t3 40
R143 a_1122_47.n2 a_1122_47.t5 40
R144 a_1122_47.n6 a_1122_47.n5 35.346
R145 a_1122_47.n48 a_1122_47.n46 28.277
R146 a_1122_47.n1 a_1122_47.t7 27.58
R147 a_1122_47.n1 a_1122_47.t4 27.58
R148 a_1122_47.n53 a_1122_47.t2 27.58
R149 a_1122_47.t1 a_1122_47.n53 27.58
R150 a_1122_47.n48 a_1122_47.n47 26.992
R151 a_1122_47.n8 a_1122_47.n7 23.778
R152 a_1122_47.n22 a_1122_47.n21 21.208
R153 a_1122_47.n36 a_1122_47.n35 19.28
R154 a_1122_47.n12 a_1122_47.n9 17.408
R155 a_1122_47.n15 a_1122_47.n12 17.408
R156 a_1122_47.n18 a_1122_47.n15 17.408
R157 a_1122_47.n20 a_1122_47.n18 17.408
R158 a_1122_47.n23 a_1122_47.n20 17.408
R159 a_1122_47.n26 a_1122_47.n23 17.408
R160 a_1122_47.n29 a_1122_47.n26 17.408
R161 a_1122_47.n32 a_1122_47.n29 17.408
R162 a_1122_47.n34 a_1122_47.n32 17.408
R163 a_1122_47.n37 a_1122_47.n34 17.408
R164 a_1122_47.n40 a_1122_47.n37 17.408
R165 a_1122_47.n43 a_1122_47.n40 17.408
R166 a_1122_47.n45 a_1122_47.n43 17.408
R167 a_1122_47.n49 a_1122_47.n45 17.408
R168 a_1122_47.n31 a_1122_47.n30 12.853
R169 a_1122_47.n11 a_1122_47.n10 12.21
R170 a_1122_47.n17 a_1122_47.n16 10.925
R171 a_1122_47.n25 a_1122_47.n24 10.282
R172 a_1122_47.n39 a_1122_47.n38 7.712
R173 a_1122_47.n42 a_1122_47.n41 3.856
R174 a_1122_47.n28 a_1122_47.n27 1.285
R175 a_1122_47.n14 a_1122_47.n13 0.642
R176 a_1122_47.n51 a_1122_47.n50 0.256
R177 X.n15 X.n13 192.158
R178 X.n15 X.n14 157.028
R179 X.n17 X.n16 157.028
R180 X.n19 X.n18 157.028
R181 X.n21 X.n20 157.028
R182 X.n23 X.n22 157.028
R183 X.n25 X.n24 157.028
R184 X.n2 X.n0 156.137
R185 X.n27 X.n26 153.34
R186 X.n2 X.n1 110.961
R187 X.n4 X.n3 110.961
R188 X.n8 X.n7 110.961
R189 X.n10 X.n9 110.961
R190 X.n12 X.n11 110.961
R191 X.n6 X.n5 109.954
R192 X X.n29 107.105
R193 X.n4 X.n2 45.176
R194 X.n10 X.n8 45.176
R195 X.n12 X.n10 45.176
R196 X.n6 X.n4 44.047
R197 X.n8 X.n6 44.047
R198 X.n0 X.t8 40
R199 X.n0 X.t20 40
R200 X.n1 X.t10 40
R201 X.n1 X.t22 40
R202 X.n3 X.t12 40
R203 X.n3 X.t15 40
R204 X.n5 X.t9 40
R205 X.n5 X.t17 40
R206 X.n7 X.t11 40
R207 X.n7 X.t13 40
R208 X.n9 X.t19 40
R209 X.n9 X.t14 40
R210 X.n11 X.t21 40
R211 X.n11 X.t16 40
R212 X.n29 X.t23 40
R213 X.n29 X.t18 40
R214 X.n17 X.n15 32
R215 X.n19 X.n17 32
R216 X.n23 X.n21 32
R217 X.n25 X.n23 32
R218 X.n21 X.n19 31.2
R219 X.n24 X.t1 27.58
R220 X.n24 X.t6 27.58
R221 X.n13 X.t5 27.58
R222 X.n13 X.t24 27.58
R223 X.n14 X.t31 27.58
R224 X.n14 X.t0 27.58
R225 X.n16 X.t7 27.58
R226 X.n16 X.t27 27.58
R227 X.n18 X.t3 27.58
R228 X.n18 X.t4 27.58
R229 X.n20 X.t30 27.58
R230 X.n20 X.t2 27.58
R231 X.n22 X.t26 27.58
R232 X.n22 X.t29 27.58
R233 X.n26 X.t25 27.58
R234 X.n26 X.t28 27.58
R235 X.n28 X.n12 13.176
R236 X.n27 X.n25 10.447
R237 X.n28 X 3.131
R238 X X.n27 1.757
R239 X X.n28 0.604
R240 KAPWR.n1 KAPWR.t5 182.874
R241 KAPWR.n23 KAPWR.t0 40.036
R242 KAPWR.n12 KAPWR.t12 28.781
R243 KAPWR.n0 KAPWR.t8 27.832
R244 KAPWR.n10 KAPWR.t7 27.827
R245 KAPWR.n8 KAPWR.t16 27.827
R246 KAPWR.n4 KAPWR.t9 27.827
R247 KAPWR.n21 KAPWR.t2 27.58
R248 KAPWR.n21 KAPWR.t1 27.58
R249 KAPWR.n6 KAPWR.t15 27.58
R250 KAPWR.n2 KAPWR.t18 27.58
R251 KAPWR.n2 KAPWR.t6 27.58
R252 KAPWR.n10 KAPWR.t11 26.878
R253 KAPWR.n8 KAPWR.t19 26.878
R254 KAPWR.n4 KAPWR.t10 26.878
R255 KAPWR.n0 KAPWR.t13 26.871
R256 KAPWR.n18 KAPWR.t3 26.595
R257 KAPWR.n6 KAPWR.t14 26.595
R258 KAPWR.n12 KAPWR.t17 25.914
R259 KAPWR.n16 KAPWR.t4 22.111
R260 KAPWR.n3 KAPWR.n2 12.576
R261 KAPWR.n7 KAPWR.n6 12.576
R262 KAPWR.n22 KAPWR.n21 12.457
R263 KAPWR.n11 KAPWR.n10 11.115
R264 KAPWR.n9 KAPWR.n8 11.115
R265 KAPWR.n5 KAPWR.n4 11.115
R266 KAPWR.n1 KAPWR.n0 11.088
R267 KAPWR.n13 KAPWR.n12 11.062
R268 KAPWR.n19 KAPWR.n18 9.3
R269 KAPWR.n17 KAPWR.n16 5.193
R270 KAPWR.n20 KAPWR.n19 4.641
R271 KAPWR.n15 KAPWR.n14 4.465
R272 KAPWR KAPWR.n23 3.222
R273 KAPWR.n18 KAPWR.n17 0.985
R274 KAPWR.n13 KAPWR.n11 0.523
R275 KAPWR.n7 KAPWR.n5 0.503
R276 KAPWR.n11 KAPWR.n9 0.496
R277 KAPWR.n23 KAPWR.n22 0.494
R278 KAPWR.n5 KAPWR.n3 0.484
R279 KAPWR.n9 KAPWR.n7 0.484
R280 KAPWR.n3 KAPWR.n1 0.481
R281 KAPWR.n15 KAPWR.n13 0.481
R282 KAPWR.n22 KAPWR.n20 0.47
R283 KAPWR.n20 KAPWR.n15 0.02
R284 a_341_47.n7 a_341_47.t17 184.766
R285 a_341_47.n8 a_341_47.t14 184.766
R286 a_341_47.n9 a_341_47.t12 184.766
R287 a_341_47.n10 a_341_47.t19 184.766
R288 a_341_47.n21 a_341_47.n20 175.576
R289 a_341_47.n20 a_341_47.n0 152.296
R290 a_341_47.n7 a_341_47.t13 146.206
R291 a_341_47.n8 a_341_47.t15 146.206
R292 a_341_47.n9 a_341_47.t18 146.206
R293 a_341_47.n10 a_341_47.t16 146.206
R294 a_341_47.n15 a_341_47.n10 114.592
R295 a_341_47.n18 a_341_47.n17 89.867
R296 a_341_47.n13 a_341_47.n11 88.89
R297 a_341_47.n13 a_341_47.n12 52.624
R298 a_341_47.n8 a_341_47.n7 40.639
R299 a_341_47.n9 a_341_47.n8 40.639
R300 a_341_47.n10 a_341_47.n9 40.639
R301 a_341_47.n0 a_341_47.t9 26.595
R302 a_341_47.n0 a_341_47.t10 26.595
R303 a_341_47.n21 a_341_47.t4 26.595
R304 a_341_47.t0 a_341_47.n21 26.595
R305 a_341_47.n14 a_341_47.n13 25.154
R306 a_341_47.n17 a_341_47.t3 24.923
R307 a_341_47.n17 a_341_47.t11 24.923
R308 a_341_47.n11 a_341_47.t8 24.923
R309 a_341_47.n11 a_341_47.t5 24.923
R310 a_341_47.n12 a_341_47.t7 24.923
R311 a_341_47.n12 a_341_47.t6 24.923
R312 a_341_47.n20 a_341_47.n19 24.436
R313 a_341_47.n5 a_341_47.t2 18.461
R314 a_341_47.n3 a_341_47.t1 15.692
R315 a_341_47.n6 a_341_47.n5 9.3
R316 a_341_47.n4 a_341_47.n3 9.23
R317 a_341_47.n5 a_341_47.n4 6.461
R318 a_341_47.n15 a_341_47.n14 4.65
R319 a_341_47.n16 a_341_47.n15 4.845
R320 a_341_47.n2 a_341_47.n1 2.666
R321 a_341_47.n19 a_341_47.n18 2.133
R322 a_341_47.n6 a_341_47.n2 1.866
R323 a_341_47.n16 a_341_47.n6 1.866
R324 a_341_47.n19 a_341_47.n16 0.533
R325 VGND.n50 VGND.t10 165.357
R326 VGND.n2 VGND.t23 153.42
R327 VGND.n46 VGND.t3 132.5
R328 VGND.n56 VGND.n55 115.464
R329 VGND.n62 VGND.n61 115.464
R330 VGND.n68 VGND.n67 115.464
R331 VGND.n37 VGND.n36 114.407
R332 VGND.n42 VGND.n41 114.407
R333 VGND.n16 VGND.n15 113.397
R334 VGND.n21 VGND.n20 113.397
R335 VGND.n6 VGND.n5 112.98
R336 VGND.n11 VGND.n10 112.98
R337 VGND.n1 VGND.n0 112.192
R338 VGND.n25 VGND.n24 112.192
R339 VGND.n31 VGND.n30 112.192
R340 VGND.n73 VGND.t28 106.288
R341 VGND.n78 VGND.t27 104.833
R342 VGND.n0 VGND.t18 40
R343 VGND.n0 VGND.t21 40
R344 VGND.n5 VGND.t16 40
R345 VGND.n5 VGND.t19 40
R346 VGND.n10 VGND.t14 40
R347 VGND.n10 VGND.t11 40
R348 VGND.n15 VGND.t25 40
R349 VGND.n20 VGND.t17 40
R350 VGND.n20 VGND.t12 40
R351 VGND.n24 VGND.t15 40
R352 VGND.n24 VGND.t26 40
R353 VGND.n30 VGND.t22 40
R354 VGND.n30 VGND.t24 40
R355 VGND.n36 VGND.t20 40
R356 VGND.n36 VGND.t5 40
R357 VGND.n41 VGND.t4 40
R358 VGND.n41 VGND.t2 40
R359 VGND.n15 VGND.t13 38.571
R360 VGND.n55 VGND.t7 24.923
R361 VGND.n55 VGND.t9 24.923
R362 VGND.n61 VGND.t8 24.923
R363 VGND.n61 VGND.t0 24.923
R364 VGND.n67 VGND.t1 24.923
R365 VGND.n67 VGND.t6 24.923
R366 VGND.n69 VGND.n68 14.305
R367 VGND.n63 VGND.n62 8.282
R368 VGND.n26 VGND.n25 6.023
R369 VGND.n79 VGND.n78 5.779
R370 VGND.n74 VGND.n73 4.894
R371 VGND.n4 VGND.n3 4.65
R372 VGND.n7 VGND.n6 4.65
R373 VGND.n9 VGND.n8 4.65
R374 VGND.n12 VGND.n11 4.65
R375 VGND.n14 VGND.n13 4.65
R376 VGND.n17 VGND.n16 4.65
R377 VGND.n19 VGND.n18 4.65
R378 VGND.n23 VGND.n22 4.65
R379 VGND.n27 VGND.n26 4.65
R380 VGND.n29 VGND.n28 4.65
R381 VGND.n33 VGND.n32 4.65
R382 VGND.n35 VGND.n34 4.65
R383 VGND.n38 VGND.n37 4.65
R384 VGND.n40 VGND.n39 4.65
R385 VGND.n43 VGND.n42 4.65
R386 VGND.n45 VGND.n44 4.65
R387 VGND.n48 VGND.n47 4.65
R388 VGND.n52 VGND.n51 4.65
R389 VGND.n54 VGND.n53 4.65
R390 VGND.n58 VGND.n57 4.65
R391 VGND.n60 VGND.n59 4.65
R392 VGND.n64 VGND.n63 4.65
R393 VGND.n66 VGND.n65 4.65
R394 VGND.n70 VGND.n69 4.65
R395 VGND.n72 VGND.n71 4.65
R396 VGND.n75 VGND.n74 4.65
R397 VGND.n77 VGND.n76 4.65
R398 VGND.n22 VGND.n21 4.517
R399 VGND.n2 VGND.n1 3.953
R400 VGND.n57 VGND.n56 2.258
R401 VGND.n32 VGND.n31 1.505
R402 VGND.n51 VGND.n50 0.984
R403 VGND.n47 VGND.n46 0.59
R404 VGND.n4 VGND.n2 0.242
R405 VGND.n7 VGND.n4 0.119
R406 VGND.n9 VGND.n7 0.119
R407 VGND.n12 VGND.n9 0.119
R408 VGND.n14 VGND.n12 0.119
R409 VGND.n17 VGND.n14 0.119
R410 VGND.n19 VGND.n17 0.119
R411 VGND.n23 VGND.n19 0.119
R412 VGND.n27 VGND.n23 0.119
R413 VGND.n29 VGND.n27 0.119
R414 VGND.n33 VGND.n29 0.119
R415 VGND.n35 VGND.n33 0.119
R416 VGND.n38 VGND.n35 0.119
R417 VGND.n40 VGND.n38 0.119
R418 VGND.n43 VGND.n40 0.119
R419 VGND.n45 VGND.n43 0.119
R420 VGND.n48 VGND.n45 0.119
R421 VGND.n52 VGND.n48 0.119
R422 VGND.n54 VGND.n52 0.119
R423 VGND.n58 VGND.n54 0.119
R424 VGND.n60 VGND.n58 0.119
R425 VGND.n64 VGND.n60 0.119
R426 VGND.n66 VGND.n64 0.119
R427 VGND.n70 VGND.n66 0.119
R428 VGND.n72 VGND.n70 0.119
R429 VGND.n75 VGND.n72 0.119
R430 VGND.n77 VGND.n75 0.119
R431 VGND.n79 VGND.n77 0.119
R432 VGND.n51 VGND.n49 0.098
R433 VGND VGND.n79 0.02
R434 VNB.t27 VNB 7034.27
R435 VNB.t28 VNB.t27 4690.11
R436 VNB.n0 VNB.t10 3865.64
R437 VNB.t18 VNB.t23 2782.35
R438 VNB.t21 VNB.t18 2782.35
R439 VNB.t16 VNB.t21 2782.35
R440 VNB.t19 VNB.t16 2782.35
R441 VNB.t14 VNB.t19 2782.35
R442 VNB.t11 VNB.t14 2782.35
R443 VNB.t13 VNB.t11 2782.35
R444 VNB.t17 VNB.t25 2782.35
R445 VNB.t12 VNB.t17 2782.35
R446 VNB.t15 VNB.t12 2782.35
R447 VNB.t26 VNB.t15 2782.35
R448 VNB.t22 VNB.t26 2782.35
R449 VNB.t24 VNB.t22 2782.35
R450 VNB.t20 VNB.t24 2782.35
R451 VNB.t5 VNB.t20 2782.35
R452 VNB.t4 VNB.t5 2782.35
R453 VNB.t2 VNB.t4 2782.35
R454 VNB.t3 VNB.t2 2782.35
R455 VNB.t25 VNB.t13 2750
R456 VNB VNB.n0 2717.65
R457 VNB.t10 VNB.t7 2030.77
R458 VNB.t7 VNB.t9 2030.77
R459 VNB.t9 VNB.t8 2030.77
R460 VNB.t8 VNB.t0 2030.77
R461 VNB.t0 VNB.t1 2030.77
R462 VNB.t1 VNB.t6 2030.77
R463 VNB.t6 VNB.t28 2030.77
R464 VNB.n0 VNB.t3 1585.29
R465 a_147_47.n2 a_147_47.t3 212.079
R466 a_147_47.n3 a_147_47.t4 212.079
R467 a_147_47.n4 a_147_47.t6 212.079
R468 a_147_47.n1 a_147_47.t9 212.079
R469 a_147_47.t0 a_147_47.n8 154.904
R470 a_147_47.n2 a_147_47.t7 139.779
R471 a_147_47.n3 a_147_47.t8 139.779
R472 a_147_47.n4 a_147_47.t5 139.779
R473 a_147_47.n1 a_147_47.t2 139.779
R474 a_147_47.n8 a_147_47.t1 107.578
R475 a_147_47.n6 a_147_47.n5 97.76
R476 a_147_47.n7 a_147_47.n1 73.418
R477 a_147_47.n3 a_147_47.n2 61.345
R478 a_147_47.n5 a_147_47.n3 54.042
R479 a_147_47.n7 a_147_47.n6 29.163
R480 a_147_47.n1 a_147_47.n0 18.987
R481 a_147_47.n8 a_147_47.n7 15.119
R482 a_147_47.n5 a_147_47.n4 7.303
R483 A.n0 A.t1 229.752
R484 A.n0 A.t0 157.452
R485 A A.n0 86.448
C0 X VGND 1.57fF
C1 VPWR X 0.49fF
C2 KAPWR X 1.87fF
C3 VPB VPWR 0.28fF
C4 KAPWR VGND 0.30fF
C5 VPWR KAPWR 6.14fF
C6 A VPWR 0.11fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__lpflow_lsbuf_lh_hl_isowell_tap_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__lpflow_lsbuf_lh_hl_isowell_tap_1 VPWR A X VPWRIN VPB VGND
X0 a_1028_32.t0 a_620_911.t5 VPWR.t3 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X1 VGND A.t0 a_714_58.t3 VGND sky130_fd_pr__nshort ad=1.4178e+12p pd=1.319e+07u as=0p ps=0u w=650000u l=150000u
X2 VGND.t3 a_505_297.t2 a_620_911.t2 VGND.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 X.t1 a_1028_32.t2 VGND VGND sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 VGND A.t1 a_714_58.t2 VGND sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 a_620_911.t4 a_505_297.t3 VGND.t19 VGND.t18 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 a_714_58.t1 A.t2 VGND VGND sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 a_714_58.t0 A.t3 VGND VGND sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 a_1028_32.t1 a_620_911.t6 VGND.t21 VGND.t20 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 VGND.t17 a_505_297.t4 a_620_911.t3 VGND.t16 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 a_505_297.t0 A.t4 VPWRIN.t1 VPWRIN.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 VPWR.t0 a_714_58.t5 a_620_911.t1 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X12 X.t0 a_1028_32.t3 VPWR.t1 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X13 VPWR.t2 a_620_911.t7 a_714_58.t4 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X14 a_505_297.t1 A.t5 VGND VGND sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15 a_620_911.t0 a_505_297.t5 VGND.t1 VGND.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
R0 a_620_911.t1 a_620_911.n7 395.249
R1 a_620_911.n6 a_620_911.t5 297.232
R2 a_620_911.n0 a_620_911.t6 244.213
R3 a_620_911.n7 a_620_911.n6 192.361
R4 a_620_911.n5 a_620_911.n1 174.104
R5 a_620_911.n6 a_620_911.t7 151.026
R6 a_620_911.n7 a_620_911.n5 122.69
R7 a_620_911.n4 a_620_911.n2 114.361
R8 a_620_911.n1 a_620_911.n0 98.006
R9 a_620_911.n5 a_620_911.n4 93.736
R10 a_620_911.n4 a_620_911.n3 74.456
R11 a_620_911.n3 a_620_911.t2 25.846
R12 a_620_911.n3 a_620_911.t0 25.846
R13 a_620_911.n2 a_620_911.t3 25.846
R14 a_620_911.n2 a_620_911.t4 25.846
R15 VPWR.n2 VPWR.n1 180.465
R16 VPWR.n2 VPWR.n0 179.493
R17 VPWR.n0 VPWR.t3 38.651
R18 VPWR.n1 VPWR.t1 37.405
R19 VPWR.n1 VPWR.t0 37.405
R20 VPWR.n0 VPWR.t2 37.405
R21 VPWR VPWR.n2 18.331
R22 a_1028_32.n1 a_1028_32.n0 704.954
R23 a_1028_32.t0 a_1028_32.n1 230.321
R24 a_1028_32.n0 a_1028_32.t2 195.911
R25 a_1028_32.n1 a_1028_32.t1 98.557
R26 a_1028_32.n0 a_1028_32.t3 59.941
R27 VPB.n2 VPB.t2 255.314
R28 VPB.t1 VPB.t0 151.06
R29 VPB.n5 VPB.n0 105.736
R30 VPB.n3 VPB.n2 7.722
R31 VPB.n5 VPB.n4 6.683
R32 VPB VPB.n5 6.548
R33 VPB.n4 VPB.n3 2.937
R34 VPB.t2 VPB.t1 1.678
R35 VPB.n2 VPB.n1 1.191
R36 A.n0 A.t0 284.379
R37 A.n3 A.t4 268.312
R38 A.n3 A.t5 165.988
R39 A.n4 A.n3 156.261
R40 A.n1 A.t1 146.206
R41 A.n0 A.t2 146.206
R42 A.n2 A.t3 146.206
R43 A.n1 A.n0 138.173
R44 A.n2 A.n1 136.773
R45 A.n4 A.n2 87.848
R46 A A.n4 78.451
R47 a_714_58.n0 a_714_58.t5 407.535
R48 a_714_58.n0 a_714_58.t4 333.495
R49 a_714_58.n2 a_714_58.n0 96.04
R50 a_714_58.n3 a_714_58.n2 73.989
R51 a_714_58.n2 a_714_58.n1 70.404
R52 a_714_58.n1 a_714_58.t2 25.846
R53 a_714_58.n1 a_714_58.t0 25.846
R54 a_714_58.t3 a_714_58.n3 25.846
R55 a_714_58.n3 a_714_58.t1 25.846
R56 VGND.n2 VGND.t20 5441.53
R57 VGND.t20 VGND.t2 3723.08
R58 VGND.t2 VGND.t0 2079.12
R59 VGND.t0 VGND.t16 2079.12
R60 VGND.t16 VGND.t18 2079.12
R61 VGND.n11 VGND.t19 108.15
R62 VGND.n8 VGND.n7 75.935
R63 VGND.n0 VGND.t21 57.23
R64 VGND.n0 VGND.t3 57.23
R65 VGND.n7 VGND.t1 25.846
R66 VGND.n7 VGND.t17 25.846
R67 VGND.n1 VGND.n0 13.427
R68 VGND.n9 VGND.n8 9.411
R69 VGND.n12 VGND.n11 6.4
R70 VGND.n4 VGND.n3 4.65
R71 VGND.n6 VGND.n5 4.65
R72 VGND.n10 VGND.n9 4.65
R73 VGND.n13 VGND.n12 4.65
R74 VGND.n15 VGND.n14 4.65
R75 VGND.n17 VGND.n16 4.65
R76 VGND.n19 VGND.n18 4.65
R77 VGND.n21 VGND.n20 4.65
R78 VGND.n23 VGND.n22 4.65
R79 VGND.n2 VGND.n1 3.972
R80 VGND.n4 VGND.n2 0.165
R81 VGND.n6 VGND.n4 0.119
R82 VGND.n10 VGND.n6 0.119
R83 VGND.n13 VGND.n10 0.119
R84 VGND.n15 VGND.n13 0.119
R85 VGND.n17 VGND.n15 0.119
R86 VGND.n19 VGND.n17 0.119
R87 VGND.n21 VGND.n19 0.119
R88 VGND.n23 VGND.n21 0.119
R89 VGND VGND.n23 0.093
R90 a_505_297.t0 a_505_297.n6 432.19
R91 a_505_297.n0 a_505_297.t2 266.706
R92 a_505_297.n5 a_505_297.n4 235.746
R93 a_505_297.n6 a_505_297.t1 194.9
R94 a_505_297.n3 a_505_297.t3 137.473
R95 a_505_297.n2 a_505_297.n0 133.353
R96 a_505_297.n0 a_505_297.t5 128.533
R97 a_505_297.n1 a_505_297.t4 117.286
R98 a_505_297.n4 a_505_297.n2 19.28
R99 a_505_297.n6 a_505_297.n5 18.133
R100 a_505_297.n2 a_505_297.n1 14.058
R101 a_505_297.n4 a_505_297.n3 4.944
R102 X X.t0 244.564
R103 X X.t1 82.073
R104 X.n0 X 16.756
R105 X X.n0 0.465
R106 X.n0 X 0.426
R107 VPWRIN.n0 VPWRIN.t0 1473.46
R108 VPWRIN.n0 VPWRIN.t1 119.279
R109 VPWRIN VPWRIN.n0 3.752
C0 VPB VPWR 0.62fF
C1 VPWR X 0.12fF
C2 VPWRIN VPWR 1.43fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__lpflow_lsbuf_lh_hl_isowell_tap_2.ext - technology: sky130A

.subckt sky130_fd_sc_hd__lpflow_lsbuf_lh_hl_isowell_tap_2 VPWR A X VPWRIN VPB VGND
X0 a_1032_911.t1 a_620_911.t5 VPWR.t3 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X1 VGND A.t0 a_714_47.t3 VGND sky130_fd_pr__nshort ad=1.62905e+12p pd=1.514e+07u as=0p ps=0u w=650000u l=150000u
X2 VGND.t19 a_505_297.t2 a_620_911.t3 VGND.t18 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 X.t3 a_1032_911.t2 VPWR.t0 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 VGND A.t1 a_714_47.t2 VGND sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 a_620_911.t4 a_505_297.t3 VGND.t21 VGND.t20 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 a_714_47.t1 A.t2 VGND VGND sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 X.t1 a_1032_911.t3 VGND VGND sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 a_714_47.t0 A.t3 VGND VGND sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 VPWR.t1 a_1032_911.t4 X.t2 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 VGND a_1032_911.t5 X.t0 VGND sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 a_1032_911.t0 a_620_911.t6 VGND.t23 VGND.t22 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 VGND.t1 a_505_297.t4 a_620_911.t0 VGND.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 a_505_297.t1 A.t4 VPWRIN.t1 VPWRIN.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14 VPWR.t2 a_714_47.t5 a_620_911.t2 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X15 VPWR.t4 a_620_911.t7 a_714_47.t4 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X16 a_505_297.t0 A.t5 VGND VGND sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17 a_620_911.t1 a_505_297.t5 VGND.t3 VGND.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
R0 a_620_911.t2 a_620_911.n7 395.249
R1 a_620_911.n6 a_620_911.t5 297.232
R2 a_620_911.n0 a_620_911.t6 244.213
R3 a_620_911.n7 a_620_911.n6 192.361
R4 a_620_911.n5 a_620_911.n1 174.104
R5 a_620_911.n6 a_620_911.t7 151.026
R6 a_620_911.n7 a_620_911.n5 122.69
R7 a_620_911.n4 a_620_911.n2 114.361
R8 a_620_911.n1 a_620_911.n0 98.006
R9 a_620_911.n5 a_620_911.n4 93.736
R10 a_620_911.n4 a_620_911.n3 74.456
R11 a_620_911.n3 a_620_911.t3 25.846
R12 a_620_911.n3 a_620_911.t1 25.846
R13 a_620_911.n2 a_620_911.t0 25.846
R14 a_620_911.n2 a_620_911.t4 25.846
R15 VPWR.n3 VPWR.t1 268.841
R16 VPWR.n2 VPWR.n1 180.465
R17 VPWR.n2 VPWR.n0 179.493
R18 VPWR.n0 VPWR.t3 38.651
R19 VPWR.n1 VPWR.t0 38.412
R20 VPWR.n1 VPWR.t2 37.405
R21 VPWR.n0 VPWR.t4 37.405
R22 VPWR.n3 VPWR.n2 16.701
R23 VPWR VPWR.n3 1.63
R24 a_1032_911.n2 a_1032_911.t4 767.979
R25 a_1032_911.t1 a_1032_911.n2 230.321
R26 a_1032_911.n0 a_1032_911.t2 184.766
R27 a_1032_911.t4 a_1032_911.n1 184.766
R28 a_1032_911.n1 a_1032_911.t5 168.699
R29 a_1032_911.n0 a_1032_911.t3 168.699
R30 a_1032_911.n2 a_1032_911.t0 98.557
R31 a_1032_911.n1 a_1032_911.n0 77.12
R32 VPB.n0 VPB.t1 561.077
R33 VPB VPB.n0 48.894
R34 VPB.n0 VPB.t2 18.67
R35 VPB.t1 VPB.t0 11.974
R36 A.n0 A.t0 302.052
R37 A.n3 A.t4 268.312
R38 A.n3 A.t5 165.988
R39 A.n1 A.t1 163.879
R40 A.n0 A.t2 163.879
R41 A.n2 A.t3 163.879
R42 A.n4 A.n3 156.261
R43 A.n1 A.n0 138.173
R44 A.n2 A.n1 136.773
R45 A.n4 A.n2 87.848
R46 A A.n4 78.451
R47 a_714_47.n0 a_714_47.t5 407.535
R48 a_714_47.n0 a_714_47.t4 333.495
R49 a_714_47.n2 a_714_47.n0 96.04
R50 a_714_47.n3 a_714_47.n2 74.751
R51 a_714_47.n2 a_714_47.n1 71.165
R52 a_714_47.n1 a_714_47.t2 25.846
R53 a_714_47.n1 a_714_47.t0 25.846
R54 a_714_47.t3 a_714_47.n3 25.846
R55 a_714_47.n3 a_714_47.t1 25.846
R56 VGND.n2 VGND.t22 6561.39
R57 VGND.t22 VGND.t18 3723.08
R58 VGND.t18 VGND.t2 2079.12
R59 VGND.t2 VGND.t0 2079.12
R60 VGND.t0 VGND.t20 2079.12
R61 VGND.n11 VGND.t21 108.15
R62 VGND.n8 VGND.n7 75.935
R63 VGND.n0 VGND.t23 57.23
R64 VGND.n0 VGND.t19 57.23
R65 VGND.n7 VGND.t3 25.846
R66 VGND.n7 VGND.t1 25.846
R67 VGND.n1 VGND.n0 13.427
R68 VGND.n9 VGND.n8 9.411
R69 VGND.n12 VGND.n11 6.4
R70 VGND.n4 VGND.n3 4.65
R71 VGND.n6 VGND.n5 4.65
R72 VGND.n10 VGND.n9 4.65
R73 VGND.n13 VGND.n12 4.65
R74 VGND.n15 VGND.n14 4.65
R75 VGND.n17 VGND.n16 4.65
R76 VGND.n19 VGND.n18 4.65
R77 VGND.n21 VGND.n20 4.65
R78 VGND.n23 VGND.n22 4.65
R79 VGND.n2 VGND.n1 3.989
R80 VGND.n4 VGND.n2 0.147
R81 VGND.n6 VGND.n4 0.119
R82 VGND.n10 VGND.n6 0.119
R83 VGND.n13 VGND.n10 0.119
R84 VGND.n15 VGND.n13 0.119
R85 VGND.n17 VGND.n15 0.119
R86 VGND.n19 VGND.n17 0.119
R87 VGND.n21 VGND.n19 0.119
R88 VGND.n23 VGND.n21 0.119
R89 VGND VGND.n23 0.093
R90 a_505_297.t1 a_505_297.n6 432.19
R91 a_505_297.n0 a_505_297.t2 266.706
R92 a_505_297.n5 a_505_297.n4 235.746
R93 a_505_297.n6 a_505_297.t0 194.9
R94 a_505_297.n3 a_505_297.t3 137.473
R95 a_505_297.n2 a_505_297.n0 133.353
R96 a_505_297.n0 a_505_297.t5 128.533
R97 a_505_297.n1 a_505_297.t4 117.286
R98 a_505_297.n4 a_505_297.n2 19.28
R99 a_505_297.n6 a_505_297.n5 18.133
R100 a_505_297.n2 a_505_297.n1 14.058
R101 a_505_297.n4 a_505_297.n3 4.944
R102 X X.n1 171.871
R103 X X.n0 58.574
R104 X.n1 X.t2 45.31
R105 X.n0 X.t0 42.461
R106 X.n1 X.t3 27.58
R107 X.n0 X.t1 25.846
R108 X.n2 X 16.756
R109 X X.n2 0.465
R110 X.n2 X 0.426
R111 VPWRIN.n0 VPWRIN.t0 1473.46
R112 VPWRIN.n0 VPWRIN.t1 119.279
R113 VPWRIN VPWRIN.n0 3.752
C0 VPB VPWR 0.63fF
C1 VPWR X 0.20fF
C2 VPWRIN VPWR 1.47fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__lpflow_lsbuf_lh_hl_isowell_tap_4.ext - technology: sky130A

.subckt sky130_fd_sc_hd__lpflow_lsbuf_lh_hl_isowell_tap_4 VPWR A X VPWRIN VPB VGND
X0 a_1032_911.t1 a_620_911.t5 VPWR.t5 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X1 VPWR.t0 a_1032_911.t2 X.t3 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 VGND A.t0 a_714_47.t4 VGND sky130_fd_pr__nshort ad=1.81105e+12p pd=1.7e+07u as=0p ps=0u w=650000u l=150000u
X3 VGND.t1 a_505_297.t2 a_620_911.t1 VGND sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 X.t2 a_1032_911.t3 VPWR.t1 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 VGND A.t1 a_714_47.t3 VGND sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 a_620_911.t2 a_505_297.t3 VGND.t2 VGND sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 a_714_47.t2 A.t2 VGND VGND sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 X.t7 a_1032_911.t4 VGND VGND sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 VGND a_1032_911.t5 X.t6 VGND sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 a_714_47.t1 A.t3 VGND VGND sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 VPWR.t2 a_1032_911.t6 X.t1 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 VGND a_1032_911.t7 X.t5 VGND sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 a_1032_911.t0 a_620_911.t6 VGND.t4 VGND sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14 VGND.t3 a_505_297.t4 a_620_911.t3 VGND sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X15 a_505_297.t0 A.t4 VPWRIN.t1 VPWRIN.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16 VPWR.t6 a_714_47.t5 a_620_911.t4 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X17 X.t4 a_1032_911.t8 VGND VGND sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X18 VPWR.t4 a_620_911.t7 a_714_47.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X19 X.t0 a_1032_911.t9 VPWR.t3 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X20 a_505_297.t1 A.t5 VGND VGND sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21 a_620_911.t0 a_505_297.t5 VGND.t0 VGND sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
R0 a_620_911.t4 a_620_911.n7 395.249
R1 a_620_911.n6 a_620_911.t5 297.232
R2 a_620_911.n0 a_620_911.t6 244.213
R3 a_620_911.n7 a_620_911.n6 192.361
R4 a_620_911.n5 a_620_911.n1 174.104
R5 a_620_911.n6 a_620_911.t7 151.026
R6 a_620_911.n7 a_620_911.n5 122.69
R7 a_620_911.n4 a_620_911.n2 114.361
R8 a_620_911.n1 a_620_911.n0 98.006
R9 a_620_911.n5 a_620_911.n4 93.736
R10 a_620_911.n4 a_620_911.n3 74.456
R11 a_620_911.n3 a_620_911.t1 25.846
R12 a_620_911.n3 a_620_911.t0 25.846
R13 a_620_911.n2 a_620_911.t3 25.846
R14 a_620_911.n2 a_620_911.t2 25.846
R15 VPWR.n2 VPWR.t0 268.542
R16 VPWR.n1 VPWR.n0 186.043
R17 VPWR.n7 VPWR.n6 180.465
R18 VPWR.n7 VPWR.n5 179.493
R19 VPWR.n5 VPWR.t5 38.651
R20 VPWR.n6 VPWR.t1 38.412
R21 VPWR.n6 VPWR.t6 37.405
R22 VPWR.n5 VPWR.t4 37.405
R23 VPWR.n0 VPWR.t3 27.58
R24 VPWR.n0 VPWR.t2 27.58
R25 VPWR.n2 VPWR.n1 20.385
R26 VPWR.n8 VPWR.n7 12.8
R27 VPWR.n4 VPWR.n3 4.65
R28 VPWR.n9 VPWR.n8 4.65
R29 VPWR VPWR.n9 1.377
R30 VPWR.n4 VPWR.n2 0.45
R31 VPWR.n9 VPWR.n4 0.119
R32 a_1032_911.n4 a_1032_911.t2 461.112
R33 a_1032_911.n6 a_1032_911.n5 396.839
R34 a_1032_911.n4 a_1032_911.t9 322.939
R35 a_1032_911.n5 a_1032_911.t6 322.939
R36 a_1032_911.t1 a_1032_911.n6 230.321
R37 a_1032_911.t6 a_1032_911.n3 184.766
R38 a_1032_911.n2 a_1032_911.t3 184.766
R39 a_1032_911.n0 a_1032_911.t5 168.699
R40 a_1032_911.n1 a_1032_911.t8 168.699
R41 a_1032_911.n3 a_1032_911.t7 168.699
R42 a_1032_911.n2 a_1032_911.t4 168.699
R43 a_1032_911.n5 a_1032_911.n4 138.173
R44 a_1032_911.n6 a_1032_911.t0 98.557
R45 a_1032_911.n3 a_1032_911.n2 77.12
R46 a_1032_911.n1 a_1032_911.n0 63.772
R47 a_1032_911.n3 a_1032_911.n1 63.772
R48 VPB.n0 VPB.t2 426.91
R49 VPB VPB.n0 45.669
R50 VPB.n0 VPB.t0 12.642
R51 VPB.t2 VPB.t1 9.033
R52 X.n5 X.n3 168.613
R53 X.n6 X.n0 168.613
R54 X.n5 X.n4 70.809
R55 X X.n1 58.574
R56 X.n0 X.t1 45.31
R57 X.n1 X.t5 42.461
R58 X.n6 X.n5 36.233
R59 X.n3 X.t3 27.58
R60 X.n3 X.t0 27.58
R61 X.n0 X.t2 27.58
R62 X.n1 X.t7 25.846
R63 X.n4 X.t6 25.846
R64 X.n4 X.t4 25.846
R65 X.n6 X.n2 4.887
R66 X X.n6 3.258
R67 X.n6 X 2.363
R68 X.n2 X 0.465
R69 X.n2 X 0.426
R70 A.n0 A.t0 302.052
R71 A.n3 A.t4 268.312
R72 A.n3 A.t5 165.988
R73 A.n1 A.t1 163.879
R74 A.n0 A.t2 163.879
R75 A.n2 A.t3 163.879
R76 A.n4 A.n3 156.261
R77 A.n1 A.n0 138.173
R78 A.n2 A.n1 136.773
R79 A.n4 A.n2 87.848
R80 A A.n4 78.451
R81 a_714_47.n0 a_714_47.t5 407.535
R82 a_714_47.n0 a_714_47.t0 333.495
R83 a_714_47.n2 a_714_47.n0 96.04
R84 a_714_47.n3 a_714_47.n2 74.751
R85 a_714_47.n2 a_714_47.n1 71.165
R86 a_714_47.n1 a_714_47.t3 25.846
R87 a_714_47.n1 a_714_47.t1 25.846
R88 a_714_47.t4 a_714_47.n3 25.846
R89 a_714_47.n3 a_714_47.t2 25.846
R90 VGND.n6 VGND.t2 108.15
R91 VGND.n3 VGND.n2 75.935
R92 VGND.n0 VGND.t4 57.23
R93 VGND.n0 VGND.t1 57.23
R94 VGND.n2 VGND.t0 25.846
R95 VGND.n2 VGND.t3 25.846
R96 VGND.n1 VGND.n0 16.291
R97 VGND.n4 VGND.n3 9.411
R98 VGND.n7 VGND.n6 6.4
R99 VGND.n5 VGND.n4 4.65
R100 VGND.n8 VGND.n7 4.65
R101 VGND.n10 VGND.n9 4.65
R102 VGND.n12 VGND.n11 4.65
R103 VGND.n14 VGND.n13 4.65
R104 VGND.n16 VGND.n15 4.65
R105 VGND.n18 VGND.n17 4.65
R106 VGND.n5 VGND.n1 0.278
R107 VGND.n8 VGND.n5 0.119
R108 VGND.n10 VGND.n8 0.119
R109 VGND.n12 VGND.n10 0.119
R110 VGND.n14 VGND.n12 0.119
R111 VGND.n16 VGND.n14 0.119
R112 VGND.n18 VGND.n16 0.119
R113 VGND VGND.n18 0.093
R114 a_505_297.t0 a_505_297.n6 432.19
R115 a_505_297.n0 a_505_297.t2 266.706
R116 a_505_297.n5 a_505_297.n4 235.746
R117 a_505_297.n6 a_505_297.t1 194.9
R118 a_505_297.n3 a_505_297.t3 137.473
R119 a_505_297.n2 a_505_297.n0 133.353
R120 a_505_297.n0 a_505_297.t5 128.533
R121 a_505_297.n1 a_505_297.t4 117.286
R122 a_505_297.n4 a_505_297.n2 19.28
R123 a_505_297.n6 a_505_297.n5 18.133
R124 a_505_297.n2 a_505_297.n1 14.058
R125 a_505_297.n4 a_505_297.n3 4.944
R126 VPWRIN.n0 VPWRIN.t0 1473.46
R127 VPWRIN.n0 VPWRIN.t1 119.279
R128 VPWRIN VPWRIN.n0 3.752
C0 VPWR VPWRIN 1.65fF
C1 VPWR VPB 0.73fF
C2 VPWR X 0.50fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__lpflow_lsbuf_lh_isowell_4.ext - technology: sky130A

.subckt sky130_fd_sc_hd__lpflow_lsbuf_lh_isowell_4 VGND VPWR A X VNB VPB LOWLVPWR
X0 a_1032_911.t0 a_620_911.t5 VPWR.t5 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X1 VPWR.t0 a_1032_911.t2 X.t7 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 VGND A.t0 a_714_47.t4 VNB sky130_fd_pr__nshort ad=1.81105e+12p pd=1.7e+07u as=0p ps=0u w=650000u l=150000u
X3 VGND.t0 a_505_297.t2 a_620_911.t0 VNB sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 X.t6 a_1032_911.t3 VPWR.t1 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 VGND A.t1 a_714_47.t3 VNB sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 a_620_911.t1 a_505_297.t3 VGND.t1 VNB sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 a_714_47.t2 A.t2 VGND VNB sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 X.t3 a_1032_911.t4 VGND VNB sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 VGND a_1032_911.t5 X.t2 VNB sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 a_714_47.t1 A.t3 VGND VNB sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 VPWR.t2 a_1032_911.t6 X.t5 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 VGND a_1032_911.t7 X.t1 VNB sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 a_1032_911.t1 a_620_911.t6 VGND.t4 VNB sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14 VGND.t2 a_505_297.t4 a_620_911.t2 VNB sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X15 a_505_297.t0 A.t4 LOWLVPWR.t1 LOWLVPWR.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16 VPWR.t3 a_714_47.t5 a_620_911.t4 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X17 X.t0 a_1032_911.t8 VGND VNB sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X18 VPWR.t6 a_620_911.t7 a_714_47.t0 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X19 X.t4 a_1032_911.t9 VPWR.t4 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X20 a_505_297.t1 A.t5 VGND VNB sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21 a_620_911.t3 a_505_297.t5 VGND.t3 VNB sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
R0 a_620_911.t4 a_620_911.n7 395.249
R1 a_620_911.n6 a_620_911.t5 297.232
R2 a_620_911.n0 a_620_911.t6 244.213
R3 a_620_911.n7 a_620_911.n6 192.361
R4 a_620_911.n5 a_620_911.n1 174.104
R5 a_620_911.n6 a_620_911.t7 151.026
R6 a_620_911.n7 a_620_911.n5 122.69
R7 a_620_911.n4 a_620_911.n2 114.361
R8 a_620_911.n1 a_620_911.n0 98.006
R9 a_620_911.n5 a_620_911.n4 93.736
R10 a_620_911.n4 a_620_911.n3 74.456
R11 a_620_911.n3 a_620_911.t0 25.846
R12 a_620_911.n3 a_620_911.t3 25.846
R13 a_620_911.n2 a_620_911.t2 25.846
R14 a_620_911.n2 a_620_911.t1 25.846
R15 VPWR.n2 VPWR.t0 268.542
R16 VPWR.n1 VPWR.n0 186.043
R17 VPWR.n7 VPWR.n6 180.465
R18 VPWR.n7 VPWR.n5 179.493
R19 VPWR.n5 VPWR.t5 38.651
R20 VPWR.n6 VPWR.t1 38.412
R21 VPWR.n6 VPWR.t3 37.405
R22 VPWR.n5 VPWR.t6 37.405
R23 VPWR.n0 VPWR.t4 27.58
R24 VPWR.n0 VPWR.t2 27.58
R25 VPWR.n2 VPWR.n1 20.385
R26 VPWR.n8 VPWR.n7 12.8
R27 VPWR.n4 VPWR.n3 4.65
R28 VPWR.n9 VPWR.n8 4.65
R29 VPWR VPWR.n9 1.377
R30 VPWR.n4 VPWR.n2 0.45
R31 VPWR.n9 VPWR.n4 0.119
R32 a_1032_911.n4 a_1032_911.t2 461.112
R33 a_1032_911.n6 a_1032_911.n5 396.839
R34 a_1032_911.n4 a_1032_911.t9 322.939
R35 a_1032_911.n5 a_1032_911.t6 322.939
R36 a_1032_911.t0 a_1032_911.n6 230.321
R37 a_1032_911.t6 a_1032_911.n3 184.766
R38 a_1032_911.n2 a_1032_911.t3 184.766
R39 a_1032_911.n0 a_1032_911.t5 168.699
R40 a_1032_911.n1 a_1032_911.t8 168.699
R41 a_1032_911.n3 a_1032_911.t7 168.699
R42 a_1032_911.n2 a_1032_911.t4 168.699
R43 a_1032_911.n5 a_1032_911.n4 138.173
R44 a_1032_911.n6 a_1032_911.t1 98.557
R45 a_1032_911.n3 a_1032_911.n2 77.12
R46 a_1032_911.n1 a_1032_911.n0 63.772
R47 a_1032_911.n3 a_1032_911.n1 63.772
R48 VPB VPB.t1 290.57
R49 VPB VPB.t2 161.093
R50 VPB.t2 VPB.t0 9.033
R51 X.n5 X.n3 168.613
R52 X.n6 X.n0 168.613
R53 X.n5 X.n4 70.809
R54 X X.n1 58.574
R55 X.n0 X.t5 45.31
R56 X.n1 X.t1 42.461
R57 X.n6 X.n5 36.233
R58 X.n3 X.t7 27.58
R59 X.n3 X.t4 27.58
R60 X.n0 X.t6 27.58
R61 X.n1 X.t3 25.846
R62 X.n4 X.t2 25.846
R63 X.n4 X.t0 25.846
R64 X.n6 X.n2 4.887
R65 X X.n6 3.258
R66 X.n6 X 2.363
R67 X.n2 X 0.465
R68 X.n2 X 0.426
R69 A.n0 A.t0 302.052
R70 A.n3 A.t4 268.312
R71 A.n3 A.t5 165.988
R72 A.n1 A.t1 163.879
R73 A.n0 A.t2 163.879
R74 A.n2 A.t3 163.879
R75 A.n4 A.n3 156.261
R76 A.n1 A.n0 138.173
R77 A.n2 A.n1 136.773
R78 A.n4 A.n2 87.848
R79 A A.n4 78.451
R80 a_714_47.n0 a_714_47.t5 407.535
R81 a_714_47.n0 a_714_47.t0 333.495
R82 a_714_47.n2 a_714_47.n0 96.04
R83 a_714_47.n3 a_714_47.n2 74.751
R84 a_714_47.n2 a_714_47.n1 71.165
R85 a_714_47.n1 a_714_47.t3 25.846
R86 a_714_47.n1 a_714_47.t1 25.846
R87 a_714_47.t4 a_714_47.n3 25.846
R88 a_714_47.n3 a_714_47.t2 25.846
R89 VGND.n6 VGND.t1 108.15
R90 VGND.n3 VGND.n2 75.935
R91 VGND.n0 VGND.t4 57.23
R92 VGND.n0 VGND.t0 57.23
R93 VGND.n2 VGND.t3 25.846
R94 VGND.n2 VGND.t2 25.846
R95 VGND.n1 VGND.n0 16.292
R96 VGND.n4 VGND.n3 9.411
R97 VGND.n7 VGND.n6 6.4
R98 VGND.n5 VGND.n4 4.65
R99 VGND.n8 VGND.n7 4.65
R100 VGND VGND.n9 0.557
R101 VGND.n5 VGND.n1 0.278
R102 VGND.n9 VGND.n8 0.134
R103 VGND.n8 VGND.n5 0.119
R104 a_505_297.t0 a_505_297.n6 432.19
R105 a_505_297.n0 a_505_297.t2 266.706
R106 a_505_297.n5 a_505_297.n4 235.746
R107 a_505_297.n6 a_505_297.t1 194.9
R108 a_505_297.n3 a_505_297.t3 137.473
R109 a_505_297.n2 a_505_297.n0 133.353
R110 a_505_297.n0 a_505_297.t5 128.533
R111 a_505_297.n1 a_505_297.t4 117.286
R112 a_505_297.n4 a_505_297.n2 19.28
R113 a_505_297.n6 a_505_297.n5 18.133
R114 a_505_297.n2 a_505_297.n1 14.058
R115 a_505_297.n4 a_505_297.n3 4.944
R116 LOWLVPWR.n0 LOWLVPWR.t0 1473.46
R117 LOWLVPWR.n0 LOWLVPWR.t1 119.279
R118 LOWLVPWR LOWLVPWR.n0 3.752
C0 LOWLVPWR VGND 0.26fF
C1 LOWLVPWR VPWR 1.65fF
C2 X VGND 0.56fF
C3 VPWR X 0.50fF
C4 VPWR VGND 0.29fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__lpflow_lsbuf_lh_isowell_tap_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__lpflow_lsbuf_lh_isowell_tap_1 VPWR A X VPB VGND LOWLVPWR
X0 a_1028_32.t1 a_620_911.t5 VPWR.t0 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X1 VGND A.t0 a_714_58.t4 VGND sky130_fd_pr__nshort ad=1.4178e+12p pd=1.319e+07u as=0p ps=0u w=650000u l=150000u
X2 VGND.t5 a_505_297.t2 a_620_911.t0 VGND.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 X.t1 a_1028_32.t2 VGND VGND sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 VGND A.t1 a_714_58.t3 VGND sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 a_620_911.t1 a_505_297.t3 VGND.t7 VGND.t6 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 a_714_58.t2 A.t2 VGND VGND sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 a_714_58.t1 A.t3 VGND VGND sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 a_1028_32.t0 a_620_911.t6 VGND.t3 VGND.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 VGND.t9 a_505_297.t4 a_620_911.t2 VGND.t8 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 a_505_297.t0 A.t4 LOWLVPWR.t1 LOWLVPWR.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 VPWR.t2 a_714_58.t5 a_620_911.t4 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X12 X.t0 a_1028_32.t3 VPWR.t3 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X13 VPWR.t1 a_620_911.t7 a_714_58.t0 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X14 a_505_297.t1 A.t5 VGND VGND sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15 a_620_911.t3 a_505_297.t5 VGND.t11 VGND.t10 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
R0 a_620_911.t4 a_620_911.n7 395.249
R1 a_620_911.n6 a_620_911.t5 297.232
R2 a_620_911.n0 a_620_911.t6 244.213
R3 a_620_911.n7 a_620_911.n6 192.361
R4 a_620_911.n5 a_620_911.n1 174.104
R5 a_620_911.n6 a_620_911.t7 151.026
R6 a_620_911.n7 a_620_911.n5 122.69
R7 a_620_911.n4 a_620_911.n2 114.361
R8 a_620_911.n1 a_620_911.n0 98.006
R9 a_620_911.n5 a_620_911.n4 93.736
R10 a_620_911.n4 a_620_911.n3 74.456
R11 a_620_911.n3 a_620_911.t0 25.846
R12 a_620_911.n3 a_620_911.t3 25.846
R13 a_620_911.n2 a_620_911.t2 25.846
R14 a_620_911.n2 a_620_911.t1 25.846
R15 VPWR.n2 VPWR.n1 180.465
R16 VPWR.n2 VPWR.n0 179.493
R17 VPWR.n0 VPWR.t0 38.651
R18 VPWR.n1 VPWR.t3 37.405
R19 VPWR.n1 VPWR.t2 37.405
R20 VPWR.n0 VPWR.t1 37.405
R21 VPWR VPWR.n2 18.331
R22 a_1028_32.n1 a_1028_32.n0 704.954
R23 a_1028_32.t1 a_1028_32.n1 230.321
R24 a_1028_32.n0 a_1028_32.t2 195.911
R25 a_1028_32.n1 a_1028_32.t0 98.557
R26 a_1028_32.n0 a_1028_32.t3 59.941
R27 VPB.n2 VPB.t2 255.314
R28 VPB.t0 VPB.t1 151.06
R29 VPB.n5 VPB.n0 105.736
R30 VPB.n3 VPB.n2 7.722
R31 VPB.n5 VPB.n4 6.683
R32 VPB VPB.n5 6.548
R33 VPB.n4 VPB.n3 2.937
R34 VPB.t2 VPB.t0 1.678
R35 VPB.n2 VPB.n1 1.191
R36 A.n0 A.t0 284.379
R37 A.n3 A.t4 268.312
R38 A.n3 A.t5 165.988
R39 A.n4 A.n3 156.261
R40 A.n1 A.t1 146.206
R41 A.n0 A.t2 146.206
R42 A.n2 A.t3 146.206
R43 A.n1 A.n0 138.173
R44 A.n2 A.n1 136.773
R45 A.n4 A.n2 87.848
R46 A A.n4 78.451
R47 a_714_58.n0 a_714_58.t5 407.535
R48 a_714_58.n0 a_714_58.t0 333.495
R49 a_714_58.n2 a_714_58.n0 96.04
R50 a_714_58.n3 a_714_58.n2 73.989
R51 a_714_58.n2 a_714_58.n1 70.404
R52 a_714_58.n1 a_714_58.t3 25.846
R53 a_714_58.n1 a_714_58.t1 25.846
R54 a_714_58.t4 a_714_58.n3 25.846
R55 a_714_58.n3 a_714_58.t2 25.846
R56 VGND.n2 VGND.t2 5441.53
R57 VGND.t2 VGND.t4 3723.08
R58 VGND.t4 VGND.t10 2079.12
R59 VGND.t10 VGND.t8 2079.12
R60 VGND.t8 VGND.t6 2079.12
R61 VGND.n11 VGND.t7 108.15
R62 VGND.n8 VGND.n7 75.935
R63 VGND.n0 VGND.t3 57.23
R64 VGND.n0 VGND.t5 57.23
R65 VGND.n7 VGND.t11 25.846
R66 VGND.n7 VGND.t9 25.846
R67 VGND.n1 VGND.n0 13.427
R68 VGND.n9 VGND.n8 9.411
R69 VGND.n12 VGND.n11 6.4
R70 VGND.n4 VGND.n3 4.65
R71 VGND.n6 VGND.n5 4.65
R72 VGND.n10 VGND.n9 4.65
R73 VGND.n13 VGND.n12 4.65
R74 VGND.n15 VGND.n14 4.65
R75 VGND.n17 VGND.n16 4.65
R76 VGND.n19 VGND.n18 4.65
R77 VGND.n21 VGND.n20 4.65
R78 VGND.n23 VGND.n22 4.65
R79 VGND.n2 VGND.n1 3.972
R80 VGND.n4 VGND.n2 0.165
R81 VGND.n6 VGND.n4 0.119
R82 VGND.n10 VGND.n6 0.119
R83 VGND.n13 VGND.n10 0.119
R84 VGND.n15 VGND.n13 0.119
R85 VGND.n17 VGND.n15 0.119
R86 VGND.n19 VGND.n17 0.119
R87 VGND.n21 VGND.n19 0.119
R88 VGND.n23 VGND.n21 0.119
R89 VGND VGND.n23 0.093
R90 a_505_297.t0 a_505_297.n6 432.19
R91 a_505_297.n0 a_505_297.t2 266.706
R92 a_505_297.n5 a_505_297.n4 235.746
R93 a_505_297.n6 a_505_297.t1 194.9
R94 a_505_297.n3 a_505_297.t3 137.473
R95 a_505_297.n2 a_505_297.n0 133.353
R96 a_505_297.n0 a_505_297.t5 128.533
R97 a_505_297.n1 a_505_297.t4 117.286
R98 a_505_297.n4 a_505_297.n2 19.28
R99 a_505_297.n6 a_505_297.n5 18.133
R100 a_505_297.n2 a_505_297.n1 14.058
R101 a_505_297.n4 a_505_297.n3 4.944
R102 X X.t0 244.564
R103 X X.t1 82.073
R104 X.n0 X 16.756
R105 X X.n0 0.465
R106 X.n0 X 0.426
R107 LOWLVPWR.n0 LOWLVPWR.t0 1473.46
R108 LOWLVPWR.n0 LOWLVPWR.t1 119.279
R109 LOWLVPWR LOWLVPWR.n0 3.752
C0 VPB VPWR 0.62fF
C1 VPWR X 0.12fF
C2 LOWLVPWR VPWR 1.43fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__lpflow_lsbuf_lh_isowell_tap_2.ext - technology: sky130A

.subckt sky130_fd_sc_hd__lpflow_lsbuf_lh_isowell_tap_2 VPWR A X VPB VGND LOWLVPWR
X0 a_1032_911.t1 a_620_911.t5 VPWR.t3 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X1 VGND A.t0 a_714_47.t4 VGND sky130_fd_pr__nshort ad=1.62905e+12p pd=1.514e+07u as=0p ps=0u w=650000u l=150000u
X2 VGND.t7 a_505_297.t2 a_620_911.t1 VGND.t6 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 X.t3 a_1032_911.t2 VPWR.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 VGND A.t1 a_714_47.t3 VGND sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 a_620_911.t2 a_505_297.t3 VGND.t9 VGND.t8 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 a_714_47.t2 A.t2 VGND VGND sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 X.t1 a_1032_911.t3 VGND VGND sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 a_714_47.t1 A.t3 VGND VGND sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 VPWR.t1 a_1032_911.t4 X.t2 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 VGND a_1032_911.t5 X.t0 VGND sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 a_1032_911.t0 a_620_911.t6 VGND.t5 VGND.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 VGND.t11 a_505_297.t4 a_620_911.t3 VGND.t10 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 a_505_297.t0 A.t4 LOWLVPWR.t1 LOWLVPWR.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14 VPWR.t2 a_714_47.t5 a_620_911.t0 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X15 VPWR.t4 a_620_911.t7 a_714_47.t0 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X16 a_505_297.t1 A.t5 VGND VGND sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17 a_620_911.t4 a_505_297.t5 VGND.t13 VGND.t12 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
R0 a_620_911.t0 a_620_911.n7 395.249
R1 a_620_911.n6 a_620_911.t5 297.232
R2 a_620_911.n0 a_620_911.t6 244.213
R3 a_620_911.n7 a_620_911.n6 192.361
R4 a_620_911.n5 a_620_911.n1 174.104
R5 a_620_911.n6 a_620_911.t7 151.026
R6 a_620_911.n7 a_620_911.n5 122.69
R7 a_620_911.n4 a_620_911.n2 114.361
R8 a_620_911.n1 a_620_911.n0 98.006
R9 a_620_911.n5 a_620_911.n4 93.736
R10 a_620_911.n4 a_620_911.n3 74.456
R11 a_620_911.n3 a_620_911.t1 25.846
R12 a_620_911.n3 a_620_911.t4 25.846
R13 a_620_911.n2 a_620_911.t3 25.846
R14 a_620_911.n2 a_620_911.t2 25.846
R15 VPWR.n3 VPWR.t1 268.841
R16 VPWR.n2 VPWR.n1 180.465
R17 VPWR.n2 VPWR.n0 179.493
R18 VPWR.n0 VPWR.t3 38.651
R19 VPWR.n1 VPWR.t0 38.412
R20 VPWR.n1 VPWR.t2 37.405
R21 VPWR.n0 VPWR.t4 37.405
R22 VPWR.n3 VPWR.n2 16.701
R23 VPWR VPWR.n3 1.63
R24 a_1032_911.n2 a_1032_911.t4 767.979
R25 a_1032_911.t1 a_1032_911.n2 230.321
R26 a_1032_911.n0 a_1032_911.t2 184.766
R27 a_1032_911.t4 a_1032_911.n1 184.766
R28 a_1032_911.n1 a_1032_911.t5 168.699
R29 a_1032_911.n0 a_1032_911.t3 168.699
R30 a_1032_911.n2 a_1032_911.t0 98.557
R31 a_1032_911.n1 a_1032_911.n0 77.12
R32 VPB.n0 VPB.t0 561.077
R33 VPB VPB.n0 48.894
R34 VPB.n0 VPB.t2 18.67
R35 VPB.t0 VPB.t1 11.974
R36 A.n0 A.t0 302.052
R37 A.n3 A.t4 268.312
R38 A.n3 A.t5 165.988
R39 A.n1 A.t1 163.879
R40 A.n0 A.t2 163.879
R41 A.n2 A.t3 163.879
R42 A.n4 A.n3 156.261
R43 A.n1 A.n0 138.173
R44 A.n2 A.n1 136.773
R45 A.n4 A.n2 87.848
R46 A A.n4 78.451
R47 a_714_47.n0 a_714_47.t5 407.535
R48 a_714_47.n0 a_714_47.t0 333.495
R49 a_714_47.n2 a_714_47.n0 96.04
R50 a_714_47.n3 a_714_47.n2 74.751
R51 a_714_47.n2 a_714_47.n1 71.165
R52 a_714_47.n1 a_714_47.t3 25.846
R53 a_714_47.n1 a_714_47.t1 25.846
R54 a_714_47.t4 a_714_47.n3 25.846
R55 a_714_47.n3 a_714_47.t2 25.846
R56 VGND.n2 VGND.t4 6561.39
R57 VGND.t4 VGND.t6 3723.08
R58 VGND.t6 VGND.t12 2079.12
R59 VGND.t12 VGND.t10 2079.12
R60 VGND.t10 VGND.t8 2079.12
R61 VGND.n11 VGND.t9 108.15
R62 VGND.n8 VGND.n7 75.935
R63 VGND.n0 VGND.t5 57.23
R64 VGND.n0 VGND.t7 57.23
R65 VGND.n7 VGND.t13 25.846
R66 VGND.n7 VGND.t11 25.846
R67 VGND.n1 VGND.n0 13.427
R68 VGND.n9 VGND.n8 9.411
R69 VGND.n12 VGND.n11 6.4
R70 VGND.n4 VGND.n3 4.65
R71 VGND.n6 VGND.n5 4.65
R72 VGND.n10 VGND.n9 4.65
R73 VGND.n13 VGND.n12 4.65
R74 VGND.n15 VGND.n14 4.65
R75 VGND.n17 VGND.n16 4.65
R76 VGND.n19 VGND.n18 4.65
R77 VGND.n21 VGND.n20 4.65
R78 VGND.n23 VGND.n22 4.65
R79 VGND.n2 VGND.n1 3.989
R80 VGND.n4 VGND.n2 0.147
R81 VGND.n6 VGND.n4 0.119
R82 VGND.n10 VGND.n6 0.119
R83 VGND.n13 VGND.n10 0.119
R84 VGND.n15 VGND.n13 0.119
R85 VGND.n17 VGND.n15 0.119
R86 VGND.n19 VGND.n17 0.119
R87 VGND.n21 VGND.n19 0.119
R88 VGND.n23 VGND.n21 0.119
R89 VGND VGND.n23 0.093
R90 a_505_297.t0 a_505_297.n6 432.19
R91 a_505_297.n0 a_505_297.t2 266.706
R92 a_505_297.n5 a_505_297.n4 235.746
R93 a_505_297.n6 a_505_297.t1 194.9
R94 a_505_297.n3 a_505_297.t3 137.473
R95 a_505_297.n2 a_505_297.n0 133.353
R96 a_505_297.n0 a_505_297.t5 128.533
R97 a_505_297.n1 a_505_297.t4 117.286
R98 a_505_297.n4 a_505_297.n2 19.28
R99 a_505_297.n6 a_505_297.n5 18.133
R100 a_505_297.n2 a_505_297.n1 14.058
R101 a_505_297.n4 a_505_297.n3 4.944
R102 X X.n1 171.871
R103 X X.n0 58.574
R104 X.n1 X.t2 45.31
R105 X.n0 X.t0 42.461
R106 X.n1 X.t3 27.58
R107 X.n0 X.t1 25.846
R108 X.n2 X 16.756
R109 X X.n2 0.465
R110 X.n2 X 0.426
R111 LOWLVPWR.n0 LOWLVPWR.t0 1473.46
R112 LOWLVPWR.n0 LOWLVPWR.t1 119.279
R113 LOWLVPWR LOWLVPWR.n0 3.752
C0 VPB VPWR 0.63fF
C1 VPWR X 0.20fF
C2 LOWLVPWR VPWR 1.47fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__lpflow_lsbuf_lh_isowell_tap_4.ext - technology: sky130A

.subckt sky130_fd_sc_hd__lpflow_lsbuf_lh_isowell_tap_4 VPWR A X VPB VGND LOWLVPWR
X0 a_1032_911.t1 a_620_911.t5 VPWR.t5 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X1 VPWR.t0 a_1032_911.t2 X.t3 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 VGND A.t0 a_714_47.t4 VGND sky130_fd_pr__nshort ad=1.81105e+12p pd=1.7e+07u as=0p ps=0u w=650000u l=150000u
X3 VGND.t2 a_505_297.t2 a_620_911.t2 VGND sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 X.t2 a_1032_911.t3 VPWR.t1 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 VGND A.t1 a_714_47.t3 VGND sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 a_620_911.t3 a_505_297.t3 VGND.t3 VGND sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 a_714_47.t2 A.t2 VGND VGND sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 X.t7 a_1032_911.t4 VGND VGND sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 VGND a_1032_911.t5 X.t6 VGND sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 a_714_47.t1 A.t3 VGND VGND sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 VPWR.t3 a_1032_911.t6 X.t1 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 VGND a_1032_911.t7 X.t5 VGND sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 a_1032_911.t0 a_620_911.t6 VGND.t4 VGND sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14 VGND.t0 a_505_297.t4 a_620_911.t0 VGND sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X15 a_505_297.t0 A.t4 LOWLVPWR.t1 LOWLVPWR.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16 VPWR.t2 a_714_47.t5 a_620_911.t4 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X17 X.t4 a_1032_911.t8 VGND VGND sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X18 VPWR.t6 a_620_911.t7 a_714_47.t0 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X19 X.t0 a_1032_911.t9 VPWR.t4 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X20 a_505_297.t1 A.t5 VGND VGND sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21 a_620_911.t1 a_505_297.t5 VGND.t1 VGND sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
R0 a_620_911.t4 a_620_911.n7 395.249
R1 a_620_911.n6 a_620_911.t5 297.232
R2 a_620_911.n0 a_620_911.t6 244.213
R3 a_620_911.n7 a_620_911.n6 192.361
R4 a_620_911.n5 a_620_911.n1 174.104
R5 a_620_911.n6 a_620_911.t7 151.026
R6 a_620_911.n7 a_620_911.n5 122.69
R7 a_620_911.n4 a_620_911.n2 114.361
R8 a_620_911.n1 a_620_911.n0 98.006
R9 a_620_911.n5 a_620_911.n4 93.736
R10 a_620_911.n4 a_620_911.n3 74.456
R11 a_620_911.n3 a_620_911.t2 25.846
R12 a_620_911.n3 a_620_911.t1 25.846
R13 a_620_911.n2 a_620_911.t0 25.846
R14 a_620_911.n2 a_620_911.t3 25.846
R15 VPWR.n2 VPWR.t0 268.542
R16 VPWR.n1 VPWR.n0 186.043
R17 VPWR.n7 VPWR.n6 180.465
R18 VPWR.n7 VPWR.n5 179.493
R19 VPWR.n5 VPWR.t5 38.651
R20 VPWR.n6 VPWR.t1 38.412
R21 VPWR.n6 VPWR.t2 37.405
R22 VPWR.n5 VPWR.t6 37.405
R23 VPWR.n0 VPWR.t4 27.58
R24 VPWR.n0 VPWR.t3 27.58
R25 VPWR.n2 VPWR.n1 20.385
R26 VPWR.n8 VPWR.n7 12.8
R27 VPWR.n4 VPWR.n3 4.65
R28 VPWR.n9 VPWR.n8 4.65
R29 VPWR VPWR.n9 1.377
R30 VPWR.n4 VPWR.n2 0.45
R31 VPWR.n9 VPWR.n4 0.119
R32 a_1032_911.n4 a_1032_911.t2 461.112
R33 a_1032_911.n6 a_1032_911.n5 396.839
R34 a_1032_911.n4 a_1032_911.t9 322.939
R35 a_1032_911.n5 a_1032_911.t6 322.939
R36 a_1032_911.t1 a_1032_911.n6 230.321
R37 a_1032_911.t6 a_1032_911.n3 184.766
R38 a_1032_911.n2 a_1032_911.t3 184.766
R39 a_1032_911.n0 a_1032_911.t5 168.699
R40 a_1032_911.n1 a_1032_911.t8 168.699
R41 a_1032_911.n3 a_1032_911.t7 168.699
R42 a_1032_911.n2 a_1032_911.t4 168.699
R43 a_1032_911.n5 a_1032_911.n4 138.173
R44 a_1032_911.n6 a_1032_911.t0 98.557
R45 a_1032_911.n3 a_1032_911.n2 77.12
R46 a_1032_911.n1 a_1032_911.n0 63.772
R47 a_1032_911.n3 a_1032_911.n1 63.772
R48 VPB.n0 VPB.t2 426.91
R49 VPB VPB.n0 45.669
R50 VPB.n0 VPB.t1 12.642
R51 VPB.t2 VPB.t0 9.033
R52 X.n5 X.n3 168.613
R53 X.n6 X.n0 168.613
R54 X.n5 X.n4 70.809
R55 X X.n1 58.574
R56 X.n0 X.t1 45.31
R57 X.n1 X.t5 42.461
R58 X.n6 X.n5 36.233
R59 X.n3 X.t3 27.58
R60 X.n3 X.t0 27.58
R61 X.n0 X.t2 27.58
R62 X.n1 X.t7 25.846
R63 X.n4 X.t6 25.846
R64 X.n4 X.t4 25.846
R65 X.n6 X.n2 4.887
R66 X X.n6 3.258
R67 X.n6 X 2.363
R68 X.n2 X 0.465
R69 X.n2 X 0.426
R70 A.n0 A.t0 302.052
R71 A.n3 A.t4 268.312
R72 A.n3 A.t5 165.988
R73 A.n1 A.t1 163.879
R74 A.n0 A.t2 163.879
R75 A.n2 A.t3 163.879
R76 A.n4 A.n3 156.261
R77 A.n1 A.n0 138.173
R78 A.n2 A.n1 136.773
R79 A.n4 A.n2 87.848
R80 A A.n4 78.451
R81 a_714_47.n0 a_714_47.t5 407.535
R82 a_714_47.n0 a_714_47.t0 333.495
R83 a_714_47.n2 a_714_47.n0 96.04
R84 a_714_47.n3 a_714_47.n2 74.751
R85 a_714_47.n2 a_714_47.n1 71.165
R86 a_714_47.n1 a_714_47.t3 25.846
R87 a_714_47.n1 a_714_47.t1 25.846
R88 a_714_47.t4 a_714_47.n3 25.846
R89 a_714_47.n3 a_714_47.t2 25.846
R90 VGND.n6 VGND.t3 108.15
R91 VGND.n3 VGND.n2 75.935
R92 VGND.n0 VGND.t4 57.23
R93 VGND.n0 VGND.t2 57.23
R94 VGND.n2 VGND.t1 25.846
R95 VGND.n2 VGND.t0 25.846
R96 VGND.n1 VGND.n0 16.291
R97 VGND.n4 VGND.n3 9.411
R98 VGND.n7 VGND.n6 6.4
R99 VGND.n5 VGND.n4 4.65
R100 VGND.n8 VGND.n7 4.65
R101 VGND.n10 VGND.n9 4.65
R102 VGND.n12 VGND.n11 4.65
R103 VGND.n14 VGND.n13 4.65
R104 VGND.n16 VGND.n15 4.65
R105 VGND.n18 VGND.n17 4.65
R106 VGND.n5 VGND.n1 0.278
R107 VGND.n8 VGND.n5 0.119
R108 VGND.n10 VGND.n8 0.119
R109 VGND.n12 VGND.n10 0.119
R110 VGND.n14 VGND.n12 0.119
R111 VGND.n16 VGND.n14 0.119
R112 VGND.n18 VGND.n16 0.119
R113 VGND VGND.n18 0.093
R114 a_505_297.t0 a_505_297.n6 432.19
R115 a_505_297.n0 a_505_297.t2 266.706
R116 a_505_297.n5 a_505_297.n4 235.746
R117 a_505_297.n6 a_505_297.t1 194.9
R118 a_505_297.n3 a_505_297.t3 137.473
R119 a_505_297.n2 a_505_297.n0 133.353
R120 a_505_297.n0 a_505_297.t5 128.533
R121 a_505_297.n1 a_505_297.t4 117.286
R122 a_505_297.n4 a_505_297.n2 19.28
R123 a_505_297.n6 a_505_297.n5 18.133
R124 a_505_297.n2 a_505_297.n1 14.058
R125 a_505_297.n4 a_505_297.n3 4.944
R126 LOWLVPWR.n0 LOWLVPWR.t0 1473.46
R127 LOWLVPWR.n0 LOWLVPWR.t1 119.279
R128 LOWLVPWR LOWLVPWR.n0 3.752
C0 VPB VPWR 0.73fF
C1 VPWR X 0.50fF
C2 LOWLVPWR VPWR 1.65fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__macro_sparecell.ext - technology: sky130A

.subckt sky130_fd_sc_hd__nand2_2 Y A B VGND VPWR VNB VPB
X0 VPWR A Y VPB sky130_fd_pr__phighvt ad=7.9e+11p pd=7.58e+06u as=5.4e+11p ps=5.08e+06u w=1e+06u l=150000u
X1 Y A VPWR VPB sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 VPWR B Y VPB sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 a_27_47# B VGND VNB sky130_fd_pr__nshort ad=5.135e+11p pd=5.48e+06u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X4 a_27_47# A Y VNB sky130_fd_pr__nshort ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X5 Y A a_27_47# VNB sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 Y B VPWR VPB sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 VGND B a_27_47# VNB sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
C0 Y A 0.32fF
C1 Y VPWR 0.72fF
C2 Y a_27_47# 0.20fF
C3 a_27_47# B 0.13fF
C4 VGND a_27_47# 0.41fF
.ends

.subckt sky130_fd_sc_hd__inv_2 A Y VPWR VGND VNB VPB
X0 Y.t2 A.t0 VPWR.t1 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 VGND.t1 A.t1 Y.t0 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 Y.t3 A.t2 VGND.t0 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 VPWR.t0 A.t3 Y.t1 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
R0 A.n0 A.t3 212.079
R1 A.n1 A.t0 212.079
R2 A.n0 A.t1 139.779
R3 A.n1 A.t2 139.779
R4 A A.n1 113.072
R5 A.n1 A.n0 61.345
R6 VPWR.n0 VPWR.t0 162.171
R7 VPWR.n0 VPWR.t1 159.068
R8 VPWR VPWR.n0 0.126
R9 Y.n2 Y.n1 111.319
R10 Y Y.n0 50.466
R11 Y.n1 Y.t1 26.595
R12 Y.n1 Y.t2 26.595
R13 Y.n0 Y.t0 24.923
R14 Y.n0 Y.t3 24.923
R15 Y.n3 Y 11.264
R16 Y Y.n3 6.144
R17 Y.n3 Y 4.654
R18 Y Y.n2 2.048
R19 Y.n2 Y 1.551
R20 VPB.t1 VPB.t0 248.598
R21 VPB VPB.t1 198.286
R22 VGND.n0 VGND.t1 120.227
R23 VGND.n0 VGND.t0 117.585
R24 VGND VGND.n0 0.126
R25 VNB VNB.t0 6126.44
R26 VNB.t0 VNB.t1 2030.77
C0 VPWR Y 0.38fF
C1 Y VGND 0.27fF
.ends

.subckt sky130_fd_sc_hd__nor2_2 B Y A VGND VPWR VNB VPB a_27_297#
X0 Y B a_27_297# VPB sky130_fd_pr__phighvt ad=2.7e+11p pd=2.54e+06u as=8.1e+11p ps=7.62e+06u w=1e+06u l=150000u
X1 Y B VGND VNB sky130_fd_pr__nshort ad=3.51e+11p pd=3.68e+06u as=5.265e+11p ps=5.52e+06u w=650000u l=150000u
X2 a_27_297# A VPWR VPB sky130_fd_pr__phighvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X3 VGND A Y VNB sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 Y A VGND VNB sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 VGND B Y VNB sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 VPWR A a_27_297# VPB sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 a_27_297# B Y VPB sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
C0 Y B 0.25fF
C1 a_27_297# VPWR 0.50fF
C2 Y a_27_297# 0.30fF
C3 a_27_297# A 0.12fF
C4 Y VGND 0.48fF
.ends

.subckt sky130_fd_sc_hd__conb_1 LO HI VPB VNB VGND VPWR
R0 HI VPWR sky130_fd_pr__res_generic_po w=480000u l=45000u
R1 VGND LO sky130_fd_pr__res_generic_po w=480000u l=45000u
C0 HI LO 0.14fF
C1 HI VGND 0.20fF
C2 VPWR LO 0.30fF
.ends

.subckt sky130_fd_sc_hd__macro_sparecell VGND VPWR LO VNB VPB
Xsky130_fd_sc_hd__nand2_2_1 sky130_fd_sc_hd__nor2_2_1/B LO LO VGND VPWR VNB VPB sky130_fd_sc_hd__nand2_2
Xsky130_fd_sc_hd__nand2_2_0 sky130_fd_sc_hd__nor2_2_0/B LO LO VGND VPWR VNB VPB sky130_fd_sc_hd__nand2_2
Xsky130_fd_sc_hd__inv_2_0 sky130_fd_sc_hd__inv_2_0/A sky130_fd_sc_hd__inv_2_0/Y VPWR
+ VGND VNB VPB sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__inv_2_1 sky130_fd_sc_hd__inv_2_1/A sky130_fd_sc_hd__inv_2_1/Y VPWR
+ VGND VNB VPB sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__nor2_2_0 sky130_fd_sc_hd__nor2_2_0/B sky130_fd_sc_hd__inv_2_0/A
+ sky130_fd_sc_hd__nor2_2_0/B VGND VPWR VNB VPB sky130_fd_sc_hd__nor2_2_0/a_27_297#
+ sky130_fd_sc_hd__nor2_2
Xsky130_fd_sc_hd__nor2_2_1 sky130_fd_sc_hd__nor2_2_1/B sky130_fd_sc_hd__inv_2_1/A
+ sky130_fd_sc_hd__nor2_2_1/B VGND VPWR VNB VPB sky130_fd_sc_hd__nor2_2_1/a_27_297#
+ sky130_fd_sc_hd__nor2_2
Xsky130_fd_sc_hd__conb_1_0 LO sky130_fd_sc_hd__conb_1_0/HI VPB VNB VGND VPWR sky130_fd_sc_hd__conb_1
X0 VPWR LO.t8 sky130_fd_sc_hd__nor2_2_0/B VPB sky130_fd_pr__phighvt ad=3.16e+12p pd=3.032e+07u as=5.4e+11p ps=5.08e+06u w=0u l=0u
X1 sky130_fd_sc_hd__nor2_2_1/B LO.t6 VPWR VPB sky130_fd_pr__phighvt ad=5.4e+11p pd=5.08e+06u as=0p ps=0u w=0u l=0u
X2 sky130_fd_sc_hd__nand2_2_1/a_27_47# LO.t4 sky130_fd_sc_hd__nor2_2_1/B VNB sky130_fd_pr__nshort ad=5.135e+11p pd=5.48e+06u as=1.755e+11p ps=1.84e+06u w=0u l=0u
X3 sky130_fd_sc_hd__nor2_2_0/B LO.t9 VPWR VPB sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=0u l=0u
X4 sky130_fd_sc_hd__nor2_2_0/B LO.t13 sky130_fd_sc_hd__nand2_2_0/a_27_47# VNB sky130_fd_pr__nshort ad=1.755e+11p pd=1.84e+06u as=5.135e+11p ps=5.48e+06u w=0u l=0u
X5 VPWR LO.t10 sky130_fd_sc_hd__nor2_2_0/B VPB sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=0u l=0u
X6 VGND LO.t7 sky130_fd_sc_hd__nand2_2_1/a_27_47# VNB sky130_fd_pr__nshort ad=2.08e+12p pd=2.2e+07u as=0p ps=0u w=0u l=0u
X7 sky130_fd_sc_hd__nor2_2_0/B LO.t14 VPWR VPB sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=0u l=0u
X8 VPWR.t0 sky130_fd_sc_hd__inv_2_1/A sky130_fd_sc_hd__inv_2_1/Y.t2 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=0u l=0u
X9 sky130_fd_sc_hd__nor2_2_1/B LO.t5 sky130_fd_sc_hd__nand2_2_1/a_27_47# VNB sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=0u l=0u
X10 VPWR LO.t2 sky130_fd_sc_hd__nor2_2_1/B VPB sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=0u l=0u
X11 sky130_fd_sc_hd__inv_2_1/Y.t0 sky130_fd_sc_hd__inv_2_1/A VGND.t0 VNB sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=0u l=0u
X12 sky130_fd_sc_hd__nor2_2_1/B LO.t1 VPWR VPB sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=0u l=0u
X13 VGND.t1 sky130_fd_sc_hd__inv_2_1/A sky130_fd_sc_hd__inv_2_1/Y.t1 VNB sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=0u l=0u
X14 VPWR LO.t0 sky130_fd_sc_hd__nor2_2_1/B VPB sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=0u l=0u
X15 VGND LO.t15 sky130_fd_sc_hd__nand2_2_0/a_27_47# VNB sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=0u l=0u
X16 sky130_fd_sc_hd__inv_2_1/Y.t3 sky130_fd_sc_hd__inv_2_1/A VPWR.t1 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=0u l=0u
X17 sky130_fd_sc_hd__nand2_2_0/a_27_47# LO.t11 VGND VNB sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=0u l=0u
X18 sky130_fd_sc_hd__nand2_2_0/a_27_47# LO.t12 sky130_fd_sc_hd__nor2_2_0/B VNB sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=0u l=0u
X19 sky130_fd_sc_hd__nand2_2_1/a_27_47# LO.t3 VGND VNB sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=0u l=0u
R0 LO.n8 LO.t6 212.079
R1 LO.n9 LO.t2 212.079
R2 LO.n12 LO.t1 212.079
R3 LO.n13 LO.t0 212.079
R4 LO.n4 LO.t10 212.079
R5 LO.n5 LO.t14 212.079
R6 LO.n0 LO.t8 212.079
R7 LO.n1 LO.t9 212.079
R8 LO.n8 LO.t7 139.779
R9 LO.n9 LO.t3 139.779
R10 LO.n12 LO.t5 139.779
R11 LO.n13 LO.t4 139.779
R12 LO.n4 LO.t11 139.779
R13 LO.n5 LO.t15 139.779
R14 LO.n0 LO.t12 139.779
R15 LO.n1 LO.t13 139.779
R16 LO LO.n6 79.584
R17 LO.n11 LO.n10 76
R18 LO.n15 LO.n14 76
R19 LO.n3 LO.n2 76
R20 LO.n10 LO.n8 30.672
R21 LO.n10 LO.n9 30.672
R22 LO.n14 LO.n12 30.672
R23 LO.n14 LO.n13 30.672
R24 LO.n6 LO.n4 30.672
R25 LO.n6 LO.n5 30.672
R26 LO.n2 LO.n0 30.672
R27 LO.n2 LO.n1 30.672
R28 sky130_fd_sc_hd__nand2_2_1/ LO.n11 18.432
R29 LO.n19 LO.n3 15.872
R30 sky130_fd_sc_hd__nand2_2_1/ LO.n15 14.336
R31 LO.n7 LO 13.312
R32 LO.n16 sky130_fd_sc_hd__nand2_2_1/ 11.521
R33 LO.n16 sky130_fd_sc_hd__nand2_2_1/ 11.306
R34 LO.n17 LO 10.926
R35 LO.n7 sky130_fd_sc_hd__nand2_2_0/ 10.24
R36 LO.n15 LO 9.216
R37 sky130_fd_sc_hd__nand2_2_0/ LO.n19 7.168
R38 LO.n19 LO.n18 5.314
R39 LO.n11 LO 5.12
R40 LO.n18 LO.n7 4.65
R41 LO LO.n16 0.797
R42 LO.n18 LO.n17 0.664
R43 LO.n3 LO 0.512
R44 LO.n17 LO 0.046
R45 VPWR.n43 VPWR.t0 156.087
R46 VPWR.n41 VPWR.n3 128.563
R47 VPWR.n13 VPWR.n12 35.57
R48 VPWR.n36 VPWR.n4 34.635
R49 VPWR.n40 VPWR.n4 34.635
R50 VPWR.n30 VPWR.n29 34.635
R51 VPWR.n23 VPWR.n22 34.635
R52 VPWR.n17 VPWR.n16 34.635
R53 VPWR.n29 VPWR.n28 34.634
R54 VPWR.n18 VPWR.n17 34.634
R55 VPWR.n34 VPWR.n6 31.623
R56 VPWR.n41 VPWR.n40 26.729
R57 VPWR.n28 VPWR.n8 25.976
R58 VPWR.n18 VPWR.n10 25.976
R59 VPWR.n42 VPWR.n41 25.223
R60 VPWR.n43 VPWR.n42 25.223
R61 VPWR.n3 VPWR.n2 24.625
R62 VPWR.n3 VPWR.t1 24.625
R63 VPWR.n24 VPWR.n8 23.717
R64 VPWR.n22 VPWR.n10 23.717
R65 VPWR.n35 VPWR.n34 22.964
R66 VPWR.n36 VPWR.n35 21.458
R67 VPWR.n30 VPWR.n6 18.447
R68 VPWR.n16 VPWR.n12 18.447
R69 VPWR.n24 VPWR.n23 9.788
R70 VPWR.n14 VPWR.n12 4.65
R71 VPWR.n16 VPWR.n15 4.65
R72 VPWR.n17 VPWR.n11 4.65
R73 VPWR.n19 VPWR.n18 4.65
R74 VPWR.n20 VPWR.n10 4.65
R75 VPWR.n22 VPWR.n21 4.65
R76 VPWR.n23 VPWR.n9 4.65
R77 VPWR.n25 VPWR.n24 4.65
R78 VPWR.n26 VPWR.n8 4.65
R79 VPWR.n28 VPWR.n27 4.65
R80 VPWR.n29 VPWR.n7 4.65
R81 VPWR.n31 VPWR.n30 4.65
R82 VPWR.n32 VPWR.n6 4.65
R83 VPWR.n34 VPWR.n33 4.65
R84 VPWR.n35 VPWR.n5 4.65
R85 VPWR.n37 VPWR.n36 4.65
R86 VPWR.n38 VPWR.n4 4.65
R87 VPWR.n40 VPWR.n39 4.65
R88 VPWR.n41 VPWR.n1 4.65
R89 VPWR.n42 VPWR.n0 4.65
R90 VPWR VPWR.n43 4.65
R91 VPWR.n13 VPWR 0.555
R92 VPWR.n15 VPWR.n14 0.119
R93 VPWR.n15 VPWR.n11 0.119
R94 VPWR.n19 VPWR.n11 0.119
R95 VPWR.n20 VPWR.n19 0.119
R96 VPWR.n21 VPWR.n9 0.119
R97 VPWR.n25 VPWR.n9 0.119
R98 VPWR.n27 VPWR.n7 0.119
R99 VPWR.n31 VPWR.n7 0.119
R100 VPWR.n32 VPWR.n31 0.119
R101 VPWR.n33 VPWR.n32 0.119
R102 VPWR.n37 VPWR.n5 0.119
R103 VPWR.n38 VPWR.n37 0.119
R104 VPWR.n39 VPWR.n38 0.119
R105 VPWR.n39 VPWR.n1 0.119
R106 VPWR VPWR.n0 0.119
R107 VPWR.n14 VPWR 0.098
R108 VPWR.n21 VPWR 0.098
R109 VPWR.n26 VPWR 0.097
R110 VPWR VPWR.n0 0.097
R111 VPWR.n27 VPWR 0.096
R112 VPWR VPWR.n5 0.096
R113 VPWR VPWR.n13 0.041
R114 VPWR VPWR.n26 0.023
R115 VPWR.n33 VPWR 0.023
R116 VPWR VPWR.n25 0.022
R117 VPWR.n1 VPWR 0.022
R118 VPWR VPWR.n20 0.02
R119 VPB VPB 1361.37
R120 VPB VPB 1361.37
R121 VPB VPB 1358.41
R122 VPB.n0 VPB 958.878
R123 VPB VPB 819.781
R124 VPB VPB 275.233
R125 VPB.n1 VPB.n0 248.598
R126 VPB.t1 VPB.t0 248.598
R127 VPB.t0 VPB 198.286
R128 VPB VPB.n1 150.934
R129 VPB VPB.t1 97.663
R130 VGND.n2 VGND.n1 457.213
R131 VGND.n42 VGND.t1 117.781
R132 VGND.n40 VGND.t0 115.342
R133 VGND.n13 VGND.n12 34.635
R134 VGND.n14 VGND.n13 34.635
R135 VGND.n14 VGND.n8 34.635
R136 VGND.n19 VGND.n18 34.635
R137 VGND.n23 VGND.n7 34.635
R138 VGND.n24 VGND.n23 34.635
R139 VGND.n28 VGND.n6 34.635
R140 VGND.n29 VGND.n28 34.635
R141 VGND.n30 VGND.n29 34.635
R142 VGND.n36 VGND.n35 34.635
R143 VGND.n18 VGND.n8 34.634
R144 VGND.n24 VGND.n6 34.634
R145 VGND.n35 VGND.n34 34.634
R146 VGND.n12 VGND.n10 28.078
R147 VGND.n41 VGND.n40 25.223
R148 VGND.n42 VGND.n41 25.223
R149 VGND.n34 VGND.n4 24.47
R150 VGND.n30 VGND.n4 24.094
R151 VGND.n36 VGND.n2 19.952
R152 VGND.n40 VGND.n2 19.576
R153 VGND.n19 VGND.n7 9.035
R154 VGND VGND.n42 4.65
R155 VGND.n12 VGND.n11 4.65
R156 VGND.n13 VGND.n9 4.65
R157 VGND.n15 VGND.n14 4.65
R158 VGND.n16 VGND.n8 4.65
R159 VGND.n18 VGND.n17 4.65
R160 VGND.n20 VGND.n19 4.65
R161 VGND.n21 VGND.n7 4.65
R162 VGND.n23 VGND.n22 4.65
R163 VGND.n25 VGND.n24 4.65
R164 VGND.n26 VGND.n6 4.65
R165 VGND.n28 VGND.n27 4.65
R166 VGND.n29 VGND.n5 4.65
R167 VGND.n31 VGND.n30 4.65
R168 VGND.n32 VGND.n4 4.65
R169 VGND.n34 VGND.n33 4.65
R170 VGND.n35 VGND.n3 4.65
R171 VGND.n37 VGND.n36 4.65
R172 VGND.n38 VGND.n2 4.65
R173 VGND.n40 VGND.n39 4.65
R174 VGND.n41 VGND.n0 4.65
R175 VGND.n10 VGND 0.557
R176 VGND.n11 VGND.n9 0.119
R177 VGND.n15 VGND.n9 0.119
R178 VGND.n16 VGND.n15 0.119
R179 VGND.n17 VGND.n16 0.119
R180 VGND.n21 VGND.n20 0.119
R181 VGND.n22 VGND.n21 0.119
R182 VGND.n27 VGND.n26 0.119
R183 VGND.n27 VGND.n5 0.119
R184 VGND.n31 VGND.n5 0.119
R185 VGND.n32 VGND.n31 0.119
R186 VGND.n33 VGND.n3 0.119
R187 VGND.n37 VGND.n3 0.119
R188 VGND.n38 VGND.n37 0.119
R189 VGND.n39 VGND.n38 0.119
R190 VGND VGND.n0 0.119
R191 VGND.n11 VGND 0.098
R192 VGND.n20 VGND 0.098
R193 VGND.n25 VGND 0.097
R194 VGND VGND.n0 0.097
R195 VGND.n26 VGND 0.096
R196 VGND.n33 VGND 0.096
R197 VGND VGND.n10 0.039
R198 VGND VGND.n25 0.023
R199 VGND VGND.n32 0.023
R200 VGND.n22 VGND 0.022
R201 VGND.n39 VGND 0.022
R202 VGND.n17 VGND 0.02
R203 sky130_fd_sc_hd__inv_2_1/Y.n3 sky130_fd_sc_hd__inv_2_1/Y.n2 111.32
R204 sky130_fd_sc_hd__inv_2_1/Y sky130_fd_sc_hd__inv_2_1/Y.n0 50.466
R205 sky130_fd_sc_hd__inv_2_1/Y.n2 sky130_fd_sc_hd__inv_2_1/Y.t3 26.595
R206 sky130_fd_sc_hd__inv_2_1/Y.n2 sky130_fd_sc_hd__inv_2_1/Y.t2 26.595
R207 sky130_fd_sc_hd__inv_2_1/Y.n0 sky130_fd_sc_hd__inv_2_1/Y.t0 24.923
R208 sky130_fd_sc_hd__inv_2_1/Y.n0 sky130_fd_sc_hd__inv_2_1/Y.t1 24.923
R209 sky130_fd_sc_hd__inv_2_1/Y sky130_fd_sc_hd__inv_2_1/Y.n1 11.264
R210 sky130_fd_sc_hd__inv_2_1/Y.n1 sky130_fd_sc_hd__inv_2_1/Y 6.144
R211 sky130_fd_sc_hd__inv_2_1/Y.n1 sky130_fd_sc_hd__inv_2_1/Y 4.654
R212 sky130_fd_sc_hd__inv_2_1/Y.n3 sky130_fd_sc_hd__inv_2_1/Y 2.048
R213 sky130_fd_sc_hd__inv_2_1/Y sky130_fd_sc_hd__inv_2_1/Y.n3 1.551
C0 LO VGND 0.21fF
C1 VGND sky130_fd_sc_hd__nor2_2_1/B 0.14fF
C2 VGND sky130_fd_sc_hd__nor2_2_0/B 0.14fF
C3 VPWR VGND -0.19fF
C4 LO VPWR 0.33fF
C5 VPWR sky130_fd_sc_hd__nor2_2_1/a_27_297# 0.13fF
C6 VPWR sky130_fd_sc_hd__nor2_2_0/a_27_297# 0.12fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__maj3_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__maj3_1 C X B A VGND VPWR VNB VPB
X0 X.t0 a_27_47.t6 VGND.t0 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 X.t1 a_27_47.t7 VPWR.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 a_109_341.t1 C.t0 a_27_47.t5 VPB.t6 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3 a_27_47.t0 B.t0 a_265_341.t1 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 VGND.t2 A.t0 a_109_47.t0 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 a_265_341.t0 A.t1 VPWR.t1 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 VPWR.t2 A.t2 a_109_341.t0 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7 a_421_47.t0 B.t1 a_27_47.t1 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 a_265_47.t1 A.t3 VGND.t1 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9 VGND.t3 C.t1 a_421_47.t1 VNB.t6 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10 a_27_47.t2 B.t2 a_265_47.t0 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11 VPWR.t3 C.t2 a_421_341.t1 VPB.t5 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12 a_421_341.t0 B.t3 a_27_47.t3 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13 a_109_47.t1 C.t3 a_27_47.t4 VNB.t5 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
R0 a_27_47.n1 a_27_47.t5 413.667
R1 a_27_47.n5 a_27_47.n4 320.216
R2 a_27_47.n3 a_27_47.t7 236.179
R3 a_27_47.n3 a_27_47.t6 163.879
R4 a_27_47.n4 a_27_47.n3 160.48
R5 a_27_47.n1 a_27_47.t4 145.594
R6 a_27_47.n2 a_27_47.n1 98.575
R7 a_27_47.n2 a_27_47.n0 92.5
R8 a_27_47.n4 a_27_47.n2 66.26
R9 a_27_47.n5 a_27_47.t3 63.321
R10 a_27_47.t0 a_27_47.n5 63.321
R11 a_27_47.n0 a_27_47.t1 38.571
R12 a_27_47.n0 a_27_47.t2 38.571
R13 VGND.n2 VGND.n0 111.323
R14 VGND.n2 VGND.n1 111.279
R15 VGND.n1 VGND.t0 78.791
R16 VGND.n1 VGND.t3 70
R17 VGND.n0 VGND.t1 38.571
R18 VGND.n0 VGND.t2 38.571
R19 VGND VGND.n2 0.251
R20 X.n3 X.n2 292.5
R21 X.n2 X 157.814
R22 X X.n0 94.194
R23 X.n1 X.n0 92.5
R24 X.n2 X.t1 47.28
R25 X.n0 X.t0 44.307
R26 X.n5 X 15.928
R27 X.n1 X 11.105
R28 X.n4 X.n3 6.4
R29 X.n3 X 4.848
R30 X X.n5 3.413
R31 X X.n4 2.844
R32 X.n5 X 2.258
R33 X.n4 X 1.939
R34 X X.n1 1.694
R35 VNB VNB.t5 6438.23
R36 VNB.t6 VNB.t0 3882.35
R37 VNB.t3 VNB.t2 2717.65
R38 VNB.t4 VNB.t1 2717.65
R39 VNB.t2 VNB.t6 2329.41
R40 VNB.t1 VNB.t3 2329.41
R41 VNB.t5 VNB.t4 2329.41
R42 VPWR.n2 VPWR.n0 337.189
R43 VPWR.n2 VPWR.n1 174.604
R44 VPWR.n1 VPWR.t3 105.607
R45 VPWR.n0 VPWR.t1 63.321
R46 VPWR.n0 VPWR.t2 63.321
R47 VPWR.n1 VPWR.t0 57.307
R48 VPWR VPWR.n2 0.257
R49 VPB.t5 VPB.t0 423.208
R50 VPB.t3 VPB.t4 248.598
R51 VPB.t2 VPB.t1 248.598
R52 VPB.t4 VPB.t5 213.084
R53 VPB.t1 VPB.t3 213.084
R54 VPB.t6 VPB.t2 213.084
R55 VPB VPB.t6 189.408
R56 C.t2 C.t0 970.426
R57 C.t0 C.t3 472.36
R58 C.n0 C.t2 208.298
R59 C.n0 C.t1 195.445
R60 C C.n0 78.07
R61  C 12.8
R62 a_109_341.t0 a_109_341.t1 98.5
R63 B.n0 B.t3 189.586
R64 B.n1 B.t0 189.586
R65 B.n0 B.t1 176.733
R66 B.n1 B.t2 176.733
R67 B.n3 B.n2 76
R68 B.n2 B.n0 30.672
R69 B.n2 B.n1 30.672
R70  B.n3 9.007
R71 B.n3 B 1.738
R72 a_265_341.t0 a_265_341.t1 98.5
R73 A.n0 A.t1 189.586
R74 A.n1 A.t2 189.586
R75 A.n0 A.t3 176.733
R76 A.n1 A.t0 176.733
R77 A.n3 A.n2 89.381
R78 A.n2 A.n0 30.672
R79 A.n2 A.n1 30.672
R80  A.n3 9.035
R81 A.n3 A 3.296
R82 a_109_47.t0 a_109_47.t1 60
R83 a_421_47.t0 a_421_47.t1 60
R84 a_265_47.t0 a_265_47.t1 60
R85 a_421_341.t0 a_421_341.t1 98.5
C0 VPWR X 0.11fF
C1 A VPWR 0.17fF
C2 C A 0.15fF
C3 C B 0.15fF
C4 A B 0.14fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__maj3_2.ext - technology: sky130A

.subckt sky130_fd_sc_hd__maj3_2 VGND VPWR B A C X VNB VPB
X0 VGND.t2 C.t0 a_441_47.t0 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1 a_285_369.t1 A.t0 VPWR.t4 VPB.t7 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X2 a_47_47.t2 B.t0 a_285_47.t0 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3 VPWR.t3 A.t1 a_129_369.t1 VPB.t6 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X4 a_129_47.t0 C.t1 a_47_47.t1 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 VPWR.t2 C.t2 a_441_369.t0 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X6 VPWR.t0 a_47_47.t6 X.t3 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 X.t1 a_47_47.t7 VGND.t0 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 a_129_369.t0 C.t3 a_47_47.t0 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X9 X.t2 a_47_47.t8 VPWR.t1 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 VGND.t3 A.t2 a_129_47.t1 VNB.t6 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11 a_441_369.t1 B.t1 a_47_47.t5 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X12 a_47_47.t3 B.t2 a_285_369.t0 VPB.t5 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X13 a_441_47.t1 B.t3 a_47_47.t4 VNB.t5 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14 VGND.t1 a_47_47.t9 X.t0 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X15 a_285_47.t1 A.t3 VGND.t4 VNB.t7 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
R0 C.n0 C.t0 321.771
R1 C.n1 C.t3 299.374
R2 C.n1 C.t1 206.188
R3 C.n0 C.t2 183.597
R4 C C.n2 140.378
R5 C.n2 C.n1 76
R6 C.n3 C.n0 76
R7 C C.n3 16.384
R8 C.n3 C 6.912
R9 C.n2  2.011
R10 a_441_47.t0 a_441_47.t1 60
R11 VGND.n4 VGND.t1 110.716
R12 VGND.n3 VGND.n2 107.239
R13 VGND.n1 VGND.n0 106.463
R14 VGND.n2 VGND.t0 88.109
R15 VGND.n2 VGND.t2 67.142
R16 VGND.n0 VGND.t4 38.571
R17 VGND.n0 VGND.t3 38.571
R18 VGND.n4 VGND.n3 5.953
R19 VGND.n6 VGND.n5 4.65
R20 VGND.n8 VGND.n7 4.65
R21 VGND.n10 VGND.n9 4.65
R22 VGND.n11 VGND.n1 3.919
R23 VGND VGND.n11 0.24
R24 VGND.n6 VGND.n4 0.201
R25 VGND.n11 VGND.n10 0.14
R26 VGND.n8 VGND.n6 0.119
R27 VGND.n10 VGND.n8 0.119
R28 VNB VNB.t2 7117.65
R29 VNB.t3 VNB.t0 4002.52
R30 VNB.t4 VNB.t5 2717.65
R31 VNB.t6 VNB.t7 2717.65
R32 VNB.t5 VNB.t3 2329.41
R33 VNB.t7 VNB.t4 2329.41
R34 VNB.t2 VNB.t6 2329.41
R35 VNB.t0 VNB.t1 2030.77
R36 A.n0 A.t0 269.919
R37 A.n1 A.t1 269.919
R38 A.n0 A.t3 176.733
R39 A.n1 A.t2 176.733
R40 A.n3 A.n2 76
R41 A.n2 A.n0 30.672
R42 A.n2 A.n1 30.672
R43 A.n3 A 14.933
R44 A A.n3 2.909
R45 VPWR.n10 VPWR.n9 307.239
R46 VPWR.n2 VPWR.n1 164.49
R47 VPWR.n0 VPWR.t0 154.768
R48 VPWR.n1 VPWR.t1 133.183
R49 VPWR.n1 VPWR.t2 41.554
R50 VPWR.n9 VPWR.t4 41.554
R51 VPWR.n9 VPWR.t3 41.554
R52 VPWR.n4 VPWR.n3 4.65
R53 VPWR.n6 VPWR.n5 4.65
R54 VPWR.n8 VPWR.n7 4.65
R55 VPWR.n11 VPWR.n10 3.919
R56 VPWR.n3 VPWR.n2 0.376
R57 VPWR VPWR.n11 0.24
R58 VPWR.n4 VPWR.n0 0.201
R59 VPWR.n11 VPWR.n8 0.14
R60 VPWR.n6 VPWR.n4 0.119
R61 VPWR.n8 VPWR.n6 0.119
R62 a_285_369.t0 a_285_369.t1 64.64
R63 VPB.t3 VPB.t1 443.925
R64 VPB VPB.t2 251.557
R65 VPB.t1 VPB.t0 248.598
R66 VPB.t5 VPB.t4 248.598
R67 VPB.t6 VPB.t7 248.598
R68 VPB.t4 VPB.t3 213.084
R69 VPB.t7 VPB.t5 213.084
R70 VPB.t2 VPB.t6 213.084
R71 B.n0 B.t1 269.919
R72 B.n1 B.t2 269.919
R73 B.n0 B.t3 176.733
R74 B.n1 B.t0 176.733
R75 B B.n2 78.427
R76 B.n2 B.n1 35.054
R77 B.n2 B.n0 26.29
R78 a_285_47.t0 a_285_47.t1 60
R79 a_47_47.n6 a_47_47.n0 238.413
R80 a_47_47.n1 a_47_47.t6 221.719
R81 a_47_47.n2 a_47_47.t8 221.719
R82 a_47_47.t0 a_47_47.n6 214.566
R83 a_47_47.n4 a_47_47.n2 192.696
R84 a_47_47.n1 a_47_47.t9 149.419
R85 a_47_47.n2 a_47_47.t7 149.419
R86 a_47_47.n5 a_47_47.t1 139.652
R87 a_47_47.n4 a_47_47.n3 107.239
R88 a_47_47.n5 a_47_47.n4 92.611
R89 a_47_47.n6 a_47_47.n5 80.571
R90 a_47_47.n2 a_47_47.n1 74.977
R91 a_47_47.n0 a_47_47.t5 41.554
R92 a_47_47.n0 a_47_47.t3 41.554
R93 a_47_47.n3 a_47_47.t4 38.571
R94 a_47_47.n3 a_47_47.t2 38.571
R95 a_129_369.t0 a_129_369.t1 64.64
R96 a_129_47.t0 a_129_47.t1 60
R97 a_441_369.t0 a_441_369.t1 64.64
R98 X.n1 X.n0 161.755
R99 X X.n2 93.469
R100 X.n0 X.t3 26.595
R101 X.n0 X.t2 26.595
R102 X.n2 X.t0 24.923
R103 X.n2 X.t1 24.923
R104 X X.n1 12.218
C0 X VGND 0.19fF
C1 A B 0.17fF
C2 C VPWR 0.12fF
C3 VPWR X 0.26fF
C4 C A 0.34fF
C5 VPWR VGND 0.11fF
C6 C B 0.18fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__maj3_4.ext - technology: sky130A

.subckt sky130_fd_sc_hd__maj3_4 X B C A VGND VPWR VNB VPB
X0 X.t7 a_47_297.t6 VGND.t6 VNB.t9 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 a_151_297.t1 C.t0 a_47_297.t4 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 VPWR.t1 A.t0 a_151_297.t0 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 VGND.t0 A.t1 a_151_47.t0 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 VGND.t5 a_47_297.t7 X.t6 VNB.t8 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 VGND.t4 a_47_297.t8 X.t5 VNB.t7 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 VPWR.t2 C.t1 a_482_297.t1 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 a_314_47.t0 A.t2 VGND.t1 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 a_482_47.t1 B.t0 a_47_297.t0 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 X.t4 a_47_297.t9 VGND.t3 VNB.t6 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 VPWR.t6 a_47_297.t10 X.t3 VPB.t9 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 a_482_297.t0 B.t1 a_47_297.t1 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 VGND.t2 C.t2 a_482_47.t0 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 X.t2 a_47_297.t11 VPWR.t5 VPB.t8 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14 a_47_297.t2 B.t2 a_314_297.t1 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 VPWR.t4 a_47_297.t12 X.t1 VPB.t7 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16 a_47_297.t3 B.t3 a_314_47.t1 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X17 a_314_297.t0 A.t3 VPWR.t0 VPB.t5 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X18 a_151_47.t1 C.t3 a_47_297.t5 VNB.t5 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X19 X.t0 a_47_297.t13 VPWR.t3 VPB.t6 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
R0 a_47_297.n13 a_47_297.n12 215.501
R1 a_47_297.n0 a_47_297.t10 212.079
R2 a_47_297.n2 a_47_297.t11 212.079
R3 a_47_297.n5 a_47_297.t12 212.079
R4 a_47_297.n6 a_47_297.t13 212.079
R5 a_47_297.n11 a_47_297.t4 199.115
R6 a_47_297.n0 a_47_297.t8 139.779
R7 a_47_297.n2 a_47_297.t9 139.779
R8 a_47_297.n5 a_47_297.t7 139.779
R9 a_47_297.n6 a_47_297.t6 139.779
R10 a_47_297.n10 a_47_297.n8 104.708
R11 a_47_297.n4 a_47_297.n1 101.6
R12 a_47_297.n11 a_47_297.t5 85.62
R13 a_47_297.n4 a_47_297.n3 76
R14 a_47_297.n8 a_47_297.n7 76
R15 a_47_297.n12 a_47_297.n11 60.871
R16 a_47_297.n10 a_47_297.n9 51.267
R17 a_47_297.n1 a_47_297.n0 30.672
R18 a_47_297.n3 a_47_297.n2 30.672
R19 a_47_297.n7 a_47_297.n5 30.672
R20 a_47_297.n7 a_47_297.n6 30.672
R21 a_47_297.t1 a_47_297.n13 26.595
R22 a_47_297.n13 a_47_297.t2 26.595
R23 a_47_297.n8 a_47_297.n4 25.6
R24 a_47_297.n9 a_47_297.t0 24.923
R25 a_47_297.n9 a_47_297.t3 24.923
R26 a_47_297.n12 a_47_297.n10 14.506
R27 VGND.n2 VGND.t4 202.953
R28 VGND.n4 VGND.n3 114.711
R29 VGND.n1 VGND.n0 107.239
R30 VGND.n10 VGND.n9 106.598
R31 VGND.n9 VGND.t2 47.076
R32 VGND.n9 VGND.t6 42.461
R33 VGND.n3 VGND.t3 24.923
R34 VGND.n3 VGND.t5 24.923
R35 VGND.n0 VGND.t1 24.923
R36 VGND.n0 VGND.t0 24.923
R37 VGND.n6 VGND.n5 4.65
R38 VGND.n8 VGND.n7 4.65
R39 VGND.n11 VGND.n10 4.65
R40 VGND.n13 VGND.n12 4.65
R41 VGND.n15 VGND.n14 4.65
R42 VGND.n17 VGND.n16 4.65
R43 VGND.n18 VGND.n1 4.112
R44 VGND.n5 VGND.n4 3.764
R45 VGND.n6 VGND.n2 0.861
R46 VGND VGND.n18 0.247
R47 VGND.n18 VGND.n17 0.134
R48 VGND.n8 VGND.n6 0.119
R49 VGND.n11 VGND.n8 0.119
R50 VGND.n13 VGND.n11 0.119
R51 VGND.n15 VGND.n13 0.119
R52 VGND.n17 VGND.n15 0.119
R53 X.n5 X.n3 146.188
R54 X.n5 X.n4 107.787
R55 X.n2 X.n0 88.17
R56 X.n2 X.n1 52.043
R57 X.n3 X.t1 26.595
R58 X.n3 X.t0 26.595
R59 X.n4 X.t3 26.595
R60 X.n4 X.t2 26.595
R61 X.n0 X.t6 24.923
R62 X.n0 X.t7 24.923
R63 X.n1 X.t5 24.923
R64 X.n1 X.t4 24.923
R65 X X.n5 17.476
R66 X.n6 X 14.523
R67 X.n6 X.n2 11.452
R68 X X.n6 2.215
R69 VNB VNB.t5 7244.34
R70 VNB.t4 VNB.t9 3070.33
R71 VNB.t6 VNB.t7 2030.77
R72 VNB.t8 VNB.t6 2030.77
R73 VNB.t9 VNB.t8 2030.77
R74 VNB.t1 VNB.t0 2030.77
R75 VNB.t3 VNB.t1 2030.77
R76 VNB.t2 VNB.t3 2030.77
R77 VNB.t5 VNB.t2 1909.89
R78 VNB.t0 VNB.t4 1740.66
R79 C C.n0 368.659
R80 C.n0 C.t1 236.549
R81 C.n1 C.t0 236.179
R82 C.n0 C.t2 164.249
R83 C.n1 C.t3 163.879
R84 C C.n1 76.914
R85 a_151_297.t0 a_151_297.t1 48.265
R86 VPB.t3 VPB.t6 375.856
R87 VPB VPB.t4 319.626
R88 VPB.t8 VPB.t9 248.598
R89 VPB.t7 VPB.t8 248.598
R90 VPB.t6 VPB.t7 248.598
R91 VPB.t1 VPB.t0 248.598
R92 VPB.t5 VPB.t1 248.598
R93 VPB.t2 VPB.t5 248.598
R94 VPB.t4 VPB.t2 233.8
R95 VPB.t0 VPB.t3 213.084
R96 A.n0 A.t3 212.079
R97 A.n1 A.t0 212.079
R98 A.n0 A.t2 139.779
R99 A.n1 A.t1 139.779
R100 A.n3 A.n2 76
R101 A.n2 A.n0 30.672
R102 A.n2 A.n1 30.672
R103 A.n3 A 9.353
R104 A A.n3 1.805
R105 VPWR.n1 VPWR.n0 307.239
R106 VPWR.n2 VPWR.t6 205.078
R107 VPWR.n4 VPWR.n3 175.281
R108 VPWR.n10 VPWR.n9 119.91
R109 VPWR.n9 VPWR.t3 48.265
R110 VPWR.n9 VPWR.t2 47.28
R111 VPWR.n3 VPWR.t5 26.595
R112 VPWR.n3 VPWR.t4 26.595
R113 VPWR.n0 VPWR.t0 26.595
R114 VPWR.n0 VPWR.t1 26.595
R115 VPWR.n6 VPWR.n5 4.65
R116 VPWR.n8 VPWR.n7 4.65
R117 VPWR.n11 VPWR.n10 4.65
R118 VPWR.n13 VPWR.n12 4.65
R119 VPWR.n15 VPWR.n14 4.65
R120 VPWR.n17 VPWR.n16 4.65
R121 VPWR.n18 VPWR.n1 4.112
R122 VPWR.n5 VPWR.n4 3.764
R123 VPWR.n6 VPWR.n2 0.746
R124 VPWR VPWR.n18 0.247
R125 VPWR.n18 VPWR.n17 0.134
R126 VPWR.n8 VPWR.n6 0.119
R127 VPWR.n11 VPWR.n8 0.119
R128 VPWR.n13 VPWR.n11 0.119
R129 VPWR.n15 VPWR.n13 0.119
R130 VPWR.n17 VPWR.n15 0.119
R131 a_151_47.t0 a_151_47.t1 45.23
R132 a_482_297.t0 a_482_297.t1 41.37
R133 a_314_47.t0 a_314_47.t1 49.846
R134 B.n0 B.t1 212.079
R135 B.n1 B.t2 212.079
R136 B.n0 B.t0 139.779
R137 B.n1 B.t3 139.779
R138 B B.n2 83.424
R139 B.n2 B.n0 30.672
R140 B.n2 B.n1 30.672
R141 a_482_47.t0 a_482_47.t1 38.769
R142 a_314_297.t0 a_314_297.t1 53.19
C0 C B 0.12fF
C1 X VGND 0.39fF
C2 C VPWR 0.40fF
C3 VPB VPWR 0.10fF
C4 VPWR X 0.71fF
C5 C A 0.19fF
C6 VPWR VGND 0.11fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__mux2_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__mux2_1 VGND VPWR S A1 A0 X VNB VPB
X0 VPWR.t0 a_505_21.t2 a_535_374.t1 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1 a_505_21.t0 S.t0 VPWR.t2 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 a_218_374.t1 S.t1 VPWR.t3 VPB.t5 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3 VGND.t0 a_505_21.t3 a_439_47.t0 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 a_76_199.t2 A0.t0 a_218_374.t0 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 a_505_21.t1 S.t2 VGND.t2 VNB.t5 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 a_439_47.t1 A0.t1 a_76_199.t3 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7 a_535_374.t0 A1.t0 a_76_199.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 a_76_199.t1 A1.t1 a_218_47.t0 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9 a_218_47.t1 S.t3 VGND.t3 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10 VPWR.t1 a_76_199.t4 X.t0 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 VGND.t1 a_76_199.t5 X.t1 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
R0 a_505_21.t0 a_505_21.n1 410.968
R1 a_505_21.n0 a_505_21.t2 329.804
R2 a_505_21.n0 a_505_21.t3 209.596
R3 a_505_21.n1 a_505_21.t1 154.058
R4 a_505_21.n1 a_505_21.n0 126.07
R5 a_535_374.t0 a_535_374.t1 98.5
R6 VPWR.n2 VPWR.n0 348.653
R7 VPWR.n2 VPWR.n1 141.932
R8 VPWR.n1 VPWR.t3 123.494
R9 VPWR.n0 VPWR.t0 86.773
R10 VPWR.n0 VPWR.t2 68.011
R11 VPWR.n1 VPWR.t1 28.757
R12 VPWR VPWR.n2 0.139
R13 VPB.t3 VPB.t0 633.333
R14 VPB.t2 VPB.t5 322.585
R15 VPB.t5 VPB.t3 304.828
R16 VPB.t1 VPB.t4 284.112
R17 VPB.t0 VPB.t1 213.084
R18 VPB VPB.t2 59.19
R19 S S.n1 352.003
R20 S.n0 S.t2 329.901
R21 S.n1 S.t1 272.061
R22 S.n1 S.t3 206.188
R23 S.n0 S.t0 148.348
R24 S S.n0 76.673
R25 a_218_374.t0 a_218_374.t1 171.202
R26 a_439_47.t0 a_439_47.t1 94.285
R27 VGND.n13 VGND.n12 107.239
R28 VGND.n3 VGND.n2 95.288
R29 VGND.n1 VGND.n0 92.5
R30 VGND.n12 VGND.t3 74.285
R31 VGND.n0 VGND.t0 61.428
R32 VGND.n2 VGND.t2 38.571
R33 VGND.n12 VGND.t1 25.428
R34 VGND.n5 VGND.n4 4.65
R35 VGND.n7 VGND.n6 4.65
R36 VGND.n9 VGND.n8 4.65
R37 VGND.n11 VGND.n10 4.65
R38 VGND.n14 VGND.n13 3.932
R39 VGND.n5 VGND.n3 3.094
R40 VGND.n3 VGND.n1 2.626
R41 VGND.n14 VGND.n11 0.137
R42 VGND VGND.n14 0.121
R43 VGND.n7 VGND.n5 0.119
R44 VGND.n9 VGND.n7 0.119
R45 VGND.n11 VGND.n9 0.119
R46 VNB VNB.n0 6526.25
R47 VNB.t1 VNB.t5 5435.29
R48 VNB.t0 VNB.t2 4044.12
R49 VNB.t2 VNB.t1 3105.88
R50 VNB.t4 VNB.t0 3105.88
R51 VNB.n0 VNB.t3 544.086
R52 VNB.n0 VNB.t4 517.647
R53 A0.n0 A0.t0 471.287
R54 A0.n0 A0.t1 148.348
R55 A0 A0.n0 78.096
R56 a_76_199.n3 a_76_199.n2 247.831
R57 a_76_199.n0 a_76_199.t4 241.534
R58 a_76_199.t0 a_76_199.n3 207.514
R59 a_76_199.n3 a_76_199.t2 184.804
R60 a_76_199.n0 a_76_199.t5 169.234
R61 a_76_199.n2 a_76_199.n0 147.529
R62 a_76_199.n2 a_76_199.n1 113.901
R63 a_76_199.n1 a_76_199.t3 94.285
R64 a_76_199.n1 a_76_199.t1 41.428
R65 A1.n0 A1.t1 338.429
R66 A1.n0 A1.t0 224.348
R67 A1 A1.n0 29.642
R68 a_218_47.t0 a_218_47.t1 94.285
R69 X.n2 X.n1 292.5
R70 X.n3 X.n2 147.091
R71 X.n0 X.t1 117.423
R72 X.n1 X.n0 74.319
R73 X.n2 X.t0 26.595
R74 X.n3 X 10.551
R75 X.n1 X 4.776
R76 X.n0 X 2.509
R77 X X.n3 2.402
C0 A1 VGND 0.10fF
C1 S A1 0.11fF
C2 VPWR S 0.56fF
C3 A0 A1 0.38fF
C4 X VPWR 0.22fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__mux2_2.ext - technology: sky130A

.subckt sky130_fd_sc_hd__mux2_2 VGND VPWR A1 A0 S X VNB VPB
X0 VPWR.t4 S.t0 a_591_369.t1 VPB.t6 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1 a_591_369.t0 A0.t0 a_79_21.t2 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X2 VPWR.t1 a_79_21.t4 X.t1 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 a_79_21.t0 A1.t0 a_306_369.t1 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X4 VGND.t1 a_79_21.t5 X.t3 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 VGND.t4 S.t1 a_578_47.t1 VNB.t5 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 a_306_369.t0 a_257_199.t2 VPWR.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X7 a_79_21.t3 A0.t1 a_288_47.t1 VNB.t6 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 a_288_47.t0 a_257_199.t3 VGND.t2 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9 a_257_199.t1 S.t2 VGND.t3 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10 a_578_47.t0 A1.t1 a_79_21.t1 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11 X.t0 a_79_21.t6 VPWR.t2 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 a_257_199.t0 S.t3 VPWR.t3 VPB.t5 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X13 X.t2 a_79_21.t7 VGND.t0 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
R0 S.n0 S.t3 269.919
R1 S.n1 S.t0 269.919
R2 S.n0 S.t2 176.733
R3 S.n1 S.t1 176.733
R4 S.n3 S.n2 76
R5 S.n2 S.n1 31.403
R6 S.n2 S.n0 29.942
R7 S.n3 S 19.2
R8 S S.n3 3.705
R9 a_591_369.t0 a_591_369.t1 64.64
R10 VPWR.n3 VPWR.n0 318.728
R11 VPWR.n2 VPWR.n1 309.272
R12 VPWR.n6 VPWR.t2 152.162
R13 VPWR.n1 VPWR.t0 70.796
R14 VPWR.n1 VPWR.t1 46.995
R15 VPWR.n0 VPWR.t3 41.554
R16 VPWR.n0 VPWR.t4 41.554
R17 VPWR.n5 VPWR.n4 4.65
R18 VPWR.n7 VPWR.n6 4.65
R19 VPWR.n3 VPWR.n2 3.936
R20 VPWR.n5 VPWR.n3 0.14
R21 VPWR.n7 VPWR.n5 0.119
R22 VPWR VPWR.n7 0.02
R23 VPB.t0 VPB.t1 511.993
R24 VPB.t2 VPB.t0 334.423
R25 VPB.t1 VPB.t4 331.464
R26 VPB.t6 VPB.t5 248.598
R27 VPB.t3 VPB.t2 248.598
R28 VPB.t4 VPB.t6 213.084
R29 VPB VPB.t3 189.408
R30 A0.n1 A0.t0 291.73
R31 A0.n0 A0.t1 208.281
R32 A0.n1 A0 14.038
R33 A0 A0.n1 4.954
R34 A0 A0.n0 3.555
R35 A0.n0 A0 3.352
R36 a_79_21.n4 a_79_21.n3 473.24
R37 a_79_21.n1 a_79_21.t4 212.079
R38 a_79_21.n0 a_79_21.t6 212.079
R39 a_79_21.n1 a_79_21.t5 139.779
R40 a_79_21.n0 a_79_21.t7 139.779
R41 a_79_21.n3 a_79_21.n2 139.689
R42 a_79_21.n2 a_79_21.t1 102.078
R43 a_79_21.n3 a_79_21.n1 83.303
R44 a_79_21.n2 a_79_21.t3 75.266
R45 a_79_21.t0 a_79_21.n4 72.335
R46 a_79_21.n1 a_79_21.n0 61.345
R47 a_79_21.n4 a_79_21.t2 53.867
R48 X X.n2 180.864
R49 X.n1 X.n0 146.351
R50 X.n0 X.t1 26.595
R51 X.n0 X.t0 26.595
R52 X.n2 X.t3 24.923
R53 X.n2 X.t2 24.923
R54 X X.n1 10.552
R55 X.n1 X 3.409
R56 A1.n0 A1.t0 457.021
R57 A1.n0 A1.t1 135.398
R58 A1 A1.n0 81.296
R59 a_306_369.t0 a_306_369.t1 220.085
R60 VGND.n3 VGND.n0 123.523
R61 VGND.n6 VGND.t0 108.779
R62 VGND.n2 VGND.n1 107.239
R63 VGND.n1 VGND.t2 54.285
R64 VGND.n0 VGND.t3 38.571
R65 VGND.n0 VGND.t4 38.571
R66 VGND.n1 VGND.t1 25.934
R67 VGND.n7 VGND.n6 4.65
R68 VGND.n5 VGND.n4 4.65
R69 VGND.n3 VGND.n2 4.013
R70 VGND.n5 VGND.n3 0.137
R71 VGND.n7 VGND.n5 0.119
R72 VGND VGND.n7 0.02
R73 VNB.t6 VNB.t3 6308.82
R74 VNB VNB.t0 6053.91
R75 VNB.t2 VNB.t6 3073.53
R76 VNB.t3 VNB.t5 2750
R77 VNB.t5 VNB.t4 2717.65
R78 VNB.t1 VNB.t2 2255.35
R79 VNB.t0 VNB.t1 2030.77
R80 a_578_47.t0 a_578_47.t1 78.571
R81 a_257_199.n0 a_257_199.t2 299.374
R82 a_257_199.n1 a_257_199.n0 286.822
R83 a_257_199.t0 a_257_199.n1 214.451
R84 a_257_199.n0 a_257_199.t3 206.188
R85 a_257_199.n1 a_257_199.t1 192.059
R86 a_288_47.t0 a_288_47.t1 92.857
C0 VPWR VGND 0.10fF
C1 X VGND 0.15fF
C2 VPWR X 0.20fF
C3 A1 A0 0.19fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__mux2_4.ext - technology: sky130A

.subckt sky130_fd_sc_hd__mux2_4 X S A0 A1 VPWR VGND VNB VPB
X0 a_204_297.t0 A1.t0 a_396_47.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 VPWR.t3 a_396_47.t4 X.t7 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 X.t6 a_396_47.t5 VPWR.t2 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 VPWR.t5 S.t0 a_314_297.t1 VPB.t7 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 a_204_297.t1 a_27_47.t2 VPWR.t4 VPB.t6 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 a_396_47.t3 A0.t0 a_314_297.t0 VPB.t5 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 a_206_47.t0 a_27_47.t3 VGND.t0 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 X.t1 a_396_47.t6 VGND.t4 VNB.t6 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 X.t0 a_396_47.t7 VGND.t3 VNB.t5 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 VPWR.t1 a_396_47.t8 X.t5 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 a_490_47.t0 A1.t1 a_396_47.t1 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 VGND.t6 S.t1 a_490_47.t1 VNB.t8 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 VGND.t2 a_396_47.t9 X.t3 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 a_396_47.t2 A0.t1 a_206_47.t1 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14 VGND.t1 a_396_47.t10 X.t2 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X15 VPWR.t6 S.t2 a_27_47.t0 VPB.t8 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16 X.t4 a_396_47.t11 VPWR.t0 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17 VGND.t5 S.t3 a_27_47.t1 VNB.t7 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
R0 A1.n0 A1.t0 241.534
R1 A1.n0 A1.t1 169.234
R2 A1 A1.n0 90.351
R3 a_396_47.n13 a_396_47.n12 432.169
R4 a_396_47.n12 a_396_47.n0 239.321
R5 a_396_47.n1 a_396_47.t8 212.079
R6 a_396_47.n3 a_396_47.t11 212.079
R7 a_396_47.n6 a_396_47.t4 212.079
R8 a_396_47.n9 a_396_47.t5 212.079
R9 a_396_47.n1 a_396_47.t10 139.779
R10 a_396_47.n3 a_396_47.t7 139.779
R11 a_396_47.n6 a_396_47.t9 139.779
R12 a_396_47.n9 a_396_47.t6 139.779
R13 a_396_47.n5 a_396_47.n2 101.6
R14 a_396_47.n5 a_396_47.n4 76
R15 a_396_47.n8 a_396_47.n7 76
R16 a_396_47.n11 a_396_47.n10 76
R17 a_396_47.n13 a_396_47.t3 32.505
R18 a_396_47.t0 a_396_47.n13 30.535
R19 a_396_47.n0 a_396_47.t1 29.538
R20 a_396_47.n0 a_396_47.t2 29.538
R21 a_396_47.n2 a_396_47.n1 27.021
R22 a_396_47.n8 a_396_47.n5 25.6
R23 a_396_47.n11 a_396_47.n8 25.6
R24 a_396_47.n4 a_396_47.n3 15.336
R25 a_396_47.n12 a_396_47.n11 14.682
R26 a_396_47.n10 a_396_47.n9 8.033
R27 a_396_47.n7 a_396_47.n6 3.651
R28 a_204_297.t0 a_204_297.t1 810.824
R29 VPB.t0 VPB.t7 588.94
R30 VPB.t6 VPB.t5 568.224
R31 VPB.t8 VPB.t6 281.152
R32 VPB.t5 VPB.t0 278.193
R33 VPB.t1 VPB.t2 248.598
R34 VPB.t4 VPB.t1 248.598
R35 VPB.t3 VPB.t4 248.598
R36 VPB.t7 VPB.t3 248.598
R37 VPB VPB.t8 189.408
R38 X.n2 X.n1 231.818
R39 X.n5 X.n4 171.935
R40 X.n2 X.n0 168.571
R41 X.n5 X.n3 108.688
R42 X X.n2 39.07
R43 X X.n5 29.609
R44 X.n0 X.t5 26.595
R45 X.n0 X.t4 26.595
R46 X.n1 X.t7 26.595
R47 X.n1 X.t6 26.595
R48 X.n4 X.t3 24.923
R49 X.n4 X.t1 24.923
R50 X.n3 X.t2 24.923
R51 X.n3 X.t0 24.923
R52 VPWR.n6 VPWR.n5 307.239
R53 VPWR.n2 VPWR.t1 194.747
R54 VPWR.n19 VPWR.n18 165.68
R55 VPWR.n1 VPWR.n0 164.214
R56 VPWR.n18 VPWR.t4 37.43
R57 VPWR.n0 VPWR.t0 26.595
R58 VPWR.n0 VPWR.t3 26.595
R59 VPWR.n5 VPWR.t2 26.595
R60 VPWR.n5 VPWR.t5 26.595
R61 VPWR.n18 VPWR.t6 26.595
R62 VPWR.n4 VPWR.n3 4.65
R63 VPWR.n7 VPWR.n6 4.65
R64 VPWR.n9 VPWR.n8 4.65
R65 VPWR.n11 VPWR.n10 4.65
R66 VPWR.n13 VPWR.n12 4.65
R67 VPWR.n15 VPWR.n14 4.65
R68 VPWR.n17 VPWR.n16 4.65
R69 VPWR.n20 VPWR.n19 3.932
R70 VPWR.n2 VPWR.n1 3.704
R71 VPWR.n4 VPWR.n2 0.269
R72 VPWR.n20 VPWR.n17 0.137
R73 VPWR VPWR.n20 0.121
R74 VPWR.n7 VPWR.n4 0.119
R75 VPWR.n9 VPWR.n7 0.119
R76 VPWR.n11 VPWR.n9 0.119
R77 VPWR.n13 VPWR.n11 0.119
R78 VPWR.n15 VPWR.n13 0.119
R79 VPWR.n17 VPWR.n15 0.119
R80 S S.n1 275.528
R81 S.n1 S.t2 241.534
R82 S.n0 S.t0 212.079
R83 S.n1 S.t3 169.234
R84 S.n0 S.t1 139.779
R85 S S.n0 63.644
R86 a_314_297.t0 a_314_297.t1 975.255
R87 a_27_47.n0 a_27_47.t2 241.534
R88 a_27_47.t0 a_27_47.n1 196.066
R89 a_27_47.n1 a_27_47.t1 195.476
R90 a_27_47.n0 a_27_47.t3 169.234
R91 a_27_47.n1 a_27_47.n0 150.164
R92 A0.n0 A0.t0 229.752
R93 A0.n0 A0.t1 157.452
R94 A0.n1 A0.n0 76
R95 A0.n1 A0 13.511
R96 A0 A0.n1 2.607
R97 VGND.n2 VGND.t1 194.253
R98 VGND.n1 VGND.n0 107.239
R99 VGND.n6 VGND.n5 107.239
R100 VGND.n19 VGND.n18 107.239
R101 VGND.n18 VGND.t0 36.923
R102 VGND.n0 VGND.t3 24.923
R103 VGND.n0 VGND.t2 24.923
R104 VGND.n5 VGND.t4 24.923
R105 VGND.n5 VGND.t6 24.923
R106 VGND.n18 VGND.t5 24.923
R107 VGND.n4 VGND.n3 4.65
R108 VGND.n7 VGND.n6 4.65
R109 VGND.n9 VGND.n8 4.65
R110 VGND.n11 VGND.n10 4.65
R111 VGND.n13 VGND.n12 4.65
R112 VGND.n15 VGND.n14 4.65
R113 VGND.n17 VGND.n16 4.65
R114 VGND.n20 VGND.n19 3.932
R115 VGND.n2 VGND.n1 3.704
R116 VGND.n4 VGND.n2 0.269
R117 VGND.n20 VGND.n17 0.137
R118 VGND VGND.n20 0.121
R119 VGND.n7 VGND.n4 0.119
R120 VGND.n9 VGND.n7 0.119
R121 VGND.n11 VGND.n9 0.119
R122 VGND.n13 VGND.n11 0.119
R123 VGND.n15 VGND.n13 0.119
R124 VGND.n17 VGND.n15 0.119
R125 a_206_47.t0 a_206_47.t1 147.692
R126 VNB VNB.t7 6053.91
R127 VNB.t2 VNB.t8 4810.99
R128 VNB.t0 VNB.t1 4593.41
R129 VNB.t7 VNB.t0 2345.05
R130 VNB.t1 VNB.t2 2272.53
R131 VNB.t5 VNB.t3 2030.77
R132 VNB.t4 VNB.t5 2030.77
R133 VNB.t6 VNB.t4 2030.77
R134 VNB.t8 VNB.t6 2030.77
R135 a_490_47.t0 a_490_47.t1 156
C0 VPWR VGND 0.12fF
C1 S VGND 0.13fF
C2 VPB VPWR 0.11fF
C3 S A1 0.17fF
C4 X VGND 0.33fF
C5 VPWR X 0.47fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__mux2_8.ext - technology: sky130A

.subckt sky130_fd_sc_hd__mux2_8 S A1 VPWR VGND A0 X VNB VPB
X0 VGND.t7 a_79_21.t8 X.t15 VNB.t7 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 VGND.t6 a_79_21.t9 X.t14 VNB.t6 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 a_79_21.t0 A0.t0 a_792_297.t3 VPB.t16 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 X.t7 a_79_21.t10 VPWR.t7 VPB.t7 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 VPWR.t6 a_79_21.t11 X.t6 VPB.t6 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 a_1259_199.t0 S.t0 VGND.t12 VNB.t12 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 X.t5 a_79_21.t12 VPWR.t5 VPB.t5 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 a_1302_47.t3 A0.t1 a_79_21.t2 VNB.t13 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X8 VPWR.t4 a_79_21.t13 X.t4 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 a_792_297.t0 S.t1 VPWR.t8 VPB.t8 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 a_1259_199.t1 S.t2 VPWR.t9 VPB.t9 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 VGND.t5 a_79_21.t14 X.t13 VNB.t5 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 VGND.t4 a_79_21.t15 X.t12 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 VGND.t10 a_1259_199.t2 a_1302_47.t1 VNB.t10 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X14 a_79_21.t4 A1.t0 a_792_47.t3 VNB.t15 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X15 a_79_21.t3 A0.t2 a_1302_47.t2 VNB.t14 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X16 VPWR.t3 a_79_21.t16 X.t3 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17 VPWR.t10 S.t3 a_792_297.t1 VPB.t10 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X18 X.t11 a_79_21.t17 VGND.t3 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X19 a_792_297.t2 A0.t3 a_79_21.t1 VPB.t15 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X20 X.t10 a_79_21.t18 VGND.t2 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X21 X.t2 a_79_21.t19 VPWR.t2 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X22 a_1302_47.t0 a_1259_199.t3 VGND.t11 VNB.t11 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X23 VPWR.t11 a_1259_199.t4 a_1302_297.t1 VPB.t11 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X24 X.t9 a_79_21.t20 VGND.t1 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X25 a_1302_297.t0 a_1259_199.t5 VPWR.t12 VPB.t12 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X26 a_792_47.t2 A1.t1 a_79_21.t5 VNB.t16 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X27 VPWR.t1 a_79_21.t21 X.t1 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X28 a_1302_297.t3 A1.t2 a_79_21.t6 VPB.t13 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X29 VGND.t8 S.t4 a_792_47.t1 VNB.t8 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X30 X.t0 a_79_21.t22 VPWR.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X31 a_79_21.t7 A1.t3 a_1302_297.t2 VPB.t14 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X32 X.t8 a_79_21.t23 VGND.t0 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X33 a_792_47.t0 S.t5 VGND.t9 VNB.t9 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
R0 a_79_21.n26 a_79_21.n0 498.805
R1 a_79_21.n27 a_79_21.n26 292.5
R2 a_79_21.n21 a_79_21.t16 205.652
R3 a_79_21.n22 a_79_21.t19 205.652
R4 a_79_21.n17 a_79_21.t21 205.652
R5 a_79_21.n14 a_79_21.t10 205.652
R6 a_79_21.n11 a_79_21.t11 205.652
R7 a_79_21.n8 a_79_21.t12 205.652
R8 a_79_21.n6 a_79_21.t13 205.652
R9 a_79_21.n5 a_79_21.t22 205.652
R10 a_79_21.n26 a_79_21.n25 178.446
R11 a_79_21.n3 a_79_21.n1 156.103
R12 a_79_21.n21 a_79_21.t9 139.779
R13 a_79_21.n22 a_79_21.t20 139.779
R14 a_79_21.n17 a_79_21.t8 139.779
R15 a_79_21.n14 a_79_21.t18 139.779
R16 a_79_21.n11 a_79_21.t15 139.779
R17 a_79_21.n8 a_79_21.t17 139.779
R18 a_79_21.n6 a_79_21.t14 139.779
R19 a_79_21.n5 a_79_21.t23 139.779
R20 a_79_21.n10 a_79_21.n7 101.6
R21 a_79_21.n25 a_79_21.n3 95.623
R22 a_79_21.n3 a_79_21.n2 92.5
R23 a_79_21.n20 a_79_21.n4 76
R24 a_79_21.n19 a_79_21.n18 76
R25 a_79_21.n16 a_79_21.n15 76
R26 a_79_21.n13 a_79_21.n12 76
R27 a_79_21.n10 a_79_21.n9 76
R28 a_79_21.n24 a_79_21.n23 76
R29 a_79_21.n6 a_79_21.n5 57.84
R30 a_79_21.n7 a_79_21.n6 35.805
R31 a_79_21.n23 a_79_21.n21 30.297
R32 a_79_21.n23 a_79_21.n22 27.542
R33 a_79_21.n0 a_79_21.t6 26.595
R34 a_79_21.n0 a_79_21.t7 26.595
R35 a_79_21.n27 a_79_21.t1 26.595
R36 a_79_21.t0 a_79_21.n27 26.595
R37 a_79_21.n25 a_79_21.n24 26.352
R38 a_79_21.n24 a_79_21.n20 25.6
R39 a_79_21.n20 a_79_21.n19 25.6
R40 a_79_21.n19 a_79_21.n16 25.6
R41 a_79_21.n16 a_79_21.n13 25.6
R42 a_79_21.n13 a_79_21.n10 25.6
R43 a_79_21.n2 a_79_21.t5 25.312
R44 a_79_21.n2 a_79_21.t4 25.312
R45 a_79_21.n1 a_79_21.t2 25.312
R46 a_79_21.n1 a_79_21.t3 25.312
R47 a_79_21.n9 a_79_21.n8 24.788
R48 a_79_21.n12 a_79_21.n11 13.771
R49 a_79_21.n18 a_79_21.n17 8.262
R50 a_79_21.n15 a_79_21.n14 2.754
R51 X.n3 X.n2 231.818
R52 X.n6 X.n5 173.516
R53 X.n10 X.n9 168.923
R54 X.n3 X.n1 168.571
R55 X.n4 X.n0 168.571
R56 X.n13 X.n12 113.633
R57 X.n10 X.n8 108.688
R58 X.n11 X.n7 105.676
R59 X.n4 X.n3 63.247
R60 X.n11 X.n10 63.247
R61 X.n6 X.n4 53.082
R62 X.n13 X.n11 53.082
R63 X X.n6 32.29
R64 X.n2 X.t3 26.595
R65 X.n2 X.t2 26.595
R66 X.n1 X.t1 26.595
R67 X.n1 X.t7 26.595
R68 X.n0 X.t6 26.595
R69 X.n0 X.t5 26.595
R70 X.n5 X.t4 26.595
R71 X.n5 X.t0 26.595
R72 X.n7 X.t12 24.923
R73 X.n7 X.t11 24.923
R74 X.n8 X.t15 24.923
R75 X.n8 X.t10 24.923
R76 X.n9 X.t14 24.923
R77 X.n9 X.t9 24.923
R78 X.n12 X.t13 24.923
R79 X.n12 X.t8 24.923
R80 X X.n13 22.4
R81 VGND.n34 VGND.t0 190.095
R82 VGND.n3 VGND.n0 111.352
R83 VGND.n2 VGND.n1 107.239
R84 VGND.n15 VGND.n14 107.239
R85 VGND.n19 VGND.n18 107.239
R86 VGND.n25 VGND.n24 107.239
R87 VGND.n30 VGND.n29 107.239
R88 VGND.n0 VGND.t10 40.312
R89 VGND.n1 VGND.t8 37.5
R90 VGND.n14 VGND.t9 35.625
R91 VGND.n1 VGND.t11 25.312
R92 VGND.n18 VGND.t1 24.923
R93 VGND.n18 VGND.t7 24.923
R94 VGND.n24 VGND.t2 24.923
R95 VGND.n24 VGND.t4 24.923
R96 VGND.n29 VGND.t3 24.923
R97 VGND.n29 VGND.t5 24.923
R98 VGND.n0 VGND.t12 22.167
R99 VGND.n14 VGND.t6 22.167
R100 VGND.n35 VGND.n34 4.65
R101 VGND.n5 VGND.n4 4.65
R102 VGND.n7 VGND.n6 4.65
R103 VGND.n9 VGND.n8 4.65
R104 VGND.n11 VGND.n10 4.65
R105 VGND.n13 VGND.n12 4.65
R106 VGND.n17 VGND.n16 4.65
R107 VGND.n21 VGND.n20 4.65
R108 VGND.n23 VGND.n22 4.65
R109 VGND.n26 VGND.n25 4.65
R110 VGND.n28 VGND.n27 4.65
R111 VGND.n31 VGND.n30 4.65
R112 VGND.n33 VGND.n32 4.65
R113 VGND.n3 VGND.n2 3.909
R114 VGND.n20 VGND.n19 3.388
R115 VGND.n16 VGND.n15 0.376
R116 VGND.n5 VGND.n3 0.14
R117 VGND.n7 VGND.n5 0.119
R118 VGND.n9 VGND.n7 0.119
R119 VGND.n11 VGND.n9 0.119
R120 VGND.n13 VGND.n11 0.119
R121 VGND.n17 VGND.n13 0.119
R122 VGND.n21 VGND.n17 0.119
R123 VGND.n23 VGND.n21 0.119
R124 VGND.n26 VGND.n23 0.119
R125 VGND.n28 VGND.n26 0.119
R126 VGND.n31 VGND.n28 0.119
R127 VGND.n33 VGND.n31 0.119
R128 VGND.n35 VGND.n33 0.119
R129 VGND VGND.n35 0.02
R130 VNB VNB.t0 6053.91
R131 VNB.t13 VNB.t10 5866.67
R132 VNB.t16 VNB.t8 5866.67
R133 VNB.t11 VNB.t14 3104.44
R134 VNB.t8 VNB.t11 2371.11
R135 VNB.t10 VNB.t12 2309.39
R136 VNB.t6 VNB.t9 2248.62
R137 VNB.t9 VNB.t15 2175.55
R138 VNB.t14 VNB.t13 2053.33
R139 VNB.t15 VNB.t16 2053.33
R140 VNB.t1 VNB.t6 2030.77
R141 VNB.t7 VNB.t1 2030.77
R142 VNB.t2 VNB.t7 2030.77
R143 VNB.t4 VNB.t2 2030.77
R144 VNB.t3 VNB.t4 2030.77
R145 VNB.t5 VNB.t3 2030.77
R146 VNB.t0 VNB.t5 2030.77
R147 A0.n1 A0.t3 215.544
R148 A0.n2 A0.n0 203.621
R149 A0.n1 A0.t0 202.768
R150 A0.n0 A0.t1 180.319
R151 A0.n0 A0.t2 135.421
R152 A0.n2 A0.n1 126.823
R153 A0 A0.n2 4.813
R154 a_792_297.n1 a_792_297.n0 706.976
R155 a_792_297.n0 a_792_297.t3 180.255
R156 a_792_297.n0 a_792_297.t0 31.52
R157 a_792_297.n1 a_792_297.t1 26.595
R158 a_792_297.t2 a_792_297.n1 26.595
R159 VPB.t12 VPB.t14 837.538
R160 VPB.t8 VPB.t16 725.077
R161 VPB.t11 VPB.t9 295.95
R162 VPB.t10 VPB.t12 287.071
R163 VPB.t3 VPB.t8 281.152
R164 VPB.t13 VPB.t11 248.598
R165 VPB.t14 VPB.t13 248.598
R166 VPB.t15 VPB.t10 248.598
R167 VPB.t16 VPB.t15 248.598
R168 VPB.t2 VPB.t3 248.598
R169 VPB.t1 VPB.t2 248.598
R170 VPB.t7 VPB.t1 248.598
R171 VPB.t6 VPB.t7 248.598
R172 VPB.t5 VPB.t6 248.598
R173 VPB.t4 VPB.t5 248.598
R174 VPB.t0 VPB.t4 248.598
R175 VPB VPB.t0 189.408
R176 VPWR.n2 VPWR.n1 314.711
R177 VPWR.n3 VPWR.n0 311.359
R178 VPWR.n15 VPWR.n14 307.239
R179 VPWR.n34 VPWR.t0 190.542
R180 VPWR.n30 VPWR.n29 164.214
R181 VPWR.n25 VPWR.n24 164.214
R182 VPWR.n19 VPWR.n18 164.214
R183 VPWR.n0 VPWR.t11 42.355
R184 VPWR.n1 VPWR.t12 39.4
R185 VPWR.n14 VPWR.t8 37.43
R186 VPWR.n29 VPWR.t5 26.595
R187 VPWR.n29 VPWR.t4 26.595
R188 VPWR.n24 VPWR.t7 26.595
R189 VPWR.n24 VPWR.t6 26.595
R190 VPWR.n18 VPWR.t2 26.595
R191 VPWR.n18 VPWR.t1 26.595
R192 VPWR.n14 VPWR.t3 26.595
R193 VPWR.n1 VPWR.t10 26.595
R194 VPWR.n0 VPWR.t9 26.595
R195 VPWR.n3 VPWR.n2 7.904
R196 VPWR.n5 VPWR.n4 4.65
R197 VPWR.n7 VPWR.n6 4.65
R198 VPWR.n9 VPWR.n8 4.65
R199 VPWR.n11 VPWR.n10 4.65
R200 VPWR.n13 VPWR.n12 4.65
R201 VPWR.n17 VPWR.n16 4.65
R202 VPWR.n21 VPWR.n20 4.65
R203 VPWR.n23 VPWR.n22 4.65
R204 VPWR.n26 VPWR.n25 4.65
R205 VPWR.n28 VPWR.n27 4.65
R206 VPWR.n31 VPWR.n30 4.65
R207 VPWR.n33 VPWR.n32 4.65
R208 VPWR.n35 VPWR.n34 4.65
R209 VPWR.n20 VPWR.n19 3.388
R210 VPWR.n16 VPWR.n15 0.376
R211 VPWR.n5 VPWR.n3 0.134
R212 VPWR.n7 VPWR.n5 0.119
R213 VPWR.n9 VPWR.n7 0.119
R214 VPWR.n11 VPWR.n9 0.119
R215 VPWR.n13 VPWR.n11 0.119
R216 VPWR.n17 VPWR.n13 0.119
R217 VPWR.n21 VPWR.n17 0.119
R218 VPWR.n23 VPWR.n21 0.119
R219 VPWR.n26 VPWR.n23 0.119
R220 VPWR.n28 VPWR.n26 0.119
R221 VPWR.n31 VPWR.n28 0.119
R222 VPWR.n33 VPWR.n31 0.119
R223 VPWR.n35 VPWR.n33 0.119
R224 VPWR VPWR.n35 0.02
R225 S.n2 S.t3 241.534
R226 S.n1 S.t1 240.999
R227 S.n3 S.n1 237.752
R228 S.n0 S.t2 236.932
R229 S.n2 S.t4 170.841
R230 S.n1 S.t5 170.306
R231 S.n0 S.t0 164.632
R232 S S.n0 96.75
R233 S.n3 S.n2 88.975
R234 S S.n3 7.777
R235 a_1259_199.n3 a_1259_199.n2 277.411
R236 a_1259_199.t1 a_1259_199.n3 243.043
R237 a_1259_199.n0 a_1259_199.t4 239.503
R238 a_1259_199.n2 a_1259_199.t5 235.819
R239 a_1259_199.n1 a_1259_199.t0 204.763
R240 a_1259_199.n0 a_1259_199.t2 168.81
R241 a_1259_199.n2 a_1259_199.t3 165.126
R242 a_1259_199.n1 a_1259_199.n0 76
R243 a_1259_199.n3 a_1259_199.n1 25.223
R244 a_1302_47.n1 a_1302_47.n0 257.282
R245 a_1302_47.t1 a_1302_47.n1 171.562
R246 a_1302_47.n0 a_1302_47.t2 47.812
R247 a_1302_47.n0 a_1302_47.t0 43.125
R248 a_1302_47.n1 a_1302_47.t3 25.312
R249 A1.n0 A1.t3 214.859
R250 A1.n0 A1.t2 202.517
R251 A1.n1 A1.t1 177.648
R252 A1.n1 A1.t0 137.386
R253 A1 A1.n1 13.197
R254 A1 A1.n0 10.445
R255 a_792_47.n1 a_792_47.n0 248.247
R256 a_792_47.t1 a_792_47.n1 171.562
R257 a_792_47.n0 a_792_47.t0 30
R258 a_792_47.n0 a_792_47.t3 25.312
R259 a_792_47.n1 a_792_47.t2 25.312
R260 a_1302_297.n1 a_1302_297.n0 723.164
R261 a_1302_297.n0 a_1302_297.t2 222.61
R262 a_1302_297.n0 a_1302_297.t0 26.595
R263 a_1302_297.t1 a_1302_297.n1 26.595
R264 a_1302_297.n1 a_1302_297.t3 26.595
C0 X VGND 0.59fF
C1 A0 VGND 0.16fF
C2 S VPWR 0.21fF
C3 VPWR X 0.91fF
C4 S A0 0.23fF
C5 VPWR VGND 0.13fF
C6 S A1 0.71fF
C7 VPB VPWR 0.19fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__mux2i_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__mux2i_1 A1 S A0 Y VGND VPWR VNB VPB
X0 a_27_297.t0 S.t0 VPWR.t1 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 VGND.t1 S.t1 a_283_205.t0 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 a_204_297.t0 A1.t0 Y.t0 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 a_193_47.t0 A1.t1 Y.t1 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 Y.t3 A0.t0 a_27_297.t1 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 VPWR.t0 a_283_205.t2 a_204_297.t1 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 VPWR.t2 S.t2 a_283_205.t1 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 VGND.t2 a_283_205.t3 a_27_47.t1 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 a_193_47.t1 S.t3 VGND.t0 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 Y.t2 A0.t1 a_27_47.t0 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
R0 S.n1 S.t2 234.572
R1 S.n1 S.n0 225.367
R2 S.n0 S.t0 211.862
R3 S.n0 S.t3 194.406
R4 S.n2 S.t1 191.193
R5 S.n3 S.n2 97.582
R6 S.n2 S.n1 32.133
R7 S.n3 S 10.889
R8 S S.n3 2.101
R9 VPWR.n1 VPWR.t2 197.272
R10 VPWR.n1 VPWR.n0 178.25
R11 VPWR.n0 VPWR.t1 65.995
R12 VPWR.n0 VPWR.t0 52.205
R13 VPWR VPWR.n1 0.454
R14 a_27_297.t0 a_27_297.t1 458.235
R15 VPB.t2 VPB.t1 574.143
R16 VPB.t0 VPB.t2 443.925
R17 VPB.t3 VPB.t0 322.585
R18 VPB.t4 VPB.t3 269.314
R19 VPB VPB.t4 204.205
R20 a_283_205.n0 a_283_205.t2 237.785
R21 a_283_205.n0 a_283_205.t3 197.619
R22 a_283_205.t1 a_283_205.n1 157.243
R23 a_283_205.n1 a_283_205.n0 142.451
R24 a_283_205.n1 a_283_205.t0 109.483
R25 VGND.n1 VGND.t1 202.036
R26 VGND.n1 VGND.n0 119.025
R27 VGND.n0 VGND.t0 24.923
R28 VGND.n0 VGND.t2 24.923
R29 VGND VGND.n1 0.504
R30 VNB VNB.t1 6078.09
R31 VNB.t0 VNB.t4 4641.76
R32 VNB.t2 VNB.t3 4545.05
R33 VNB.t4 VNB.t2 2030.77
R34 VNB.t1 VNB.t0 2030.77
R35 A1.n0 A1.t0 234.17
R36 A1.n0 A1.t1 161.87
R37 A1 A1.n0 93.483
R38 Y.n2 Y.n1 146.375
R39  Y.n0 138.647
R40 Y.n1 Y.t0 33.49
R41 Y.n1 Y.t3 26.595
R42 Y.n0 Y.t1 24.923
R43 Y.n0 Y.t2 24.923
R44 Y.n3 Y.n2 12.55
R45 Y.n2 Y 4.228
R46 Y.n3  0.673
R47  Y.n3 0.512
R48 a_204_297.t0 a_204_297.t1 77.815
R49 a_193_47.t0 a_193_47.t1 391.508
R50 A0.n0 A0.t1 1554.34
R51 A0.n0 A0.t0 229.368
R52 A0 A0.n0 82.257
R53 a_27_47.t0 a_27_47.t1 352.648
C0 A1 Y 0.12fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__mux2i_2.ext - technology: sky130A

.subckt sky130_fd_sc_hd__mux2i_2 Y A1 A0 S VPWR VGND VNB VPB
X0 a_361_47.t1 A0.t0 Y.t3 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 Y.t1 A0.t1 a_193_297.t1 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 VPWR.t4 a_27_47.t2 a_361_297.t3 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 a_361_297.t2 a_27_47.t3 VPWR.t3 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 VPWR.t0 S.t0 a_193_297.t2 VPB.t6 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 Y.t2 A0.t2 a_361_47.t0 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 a_193_297.t3 S.t1 VPWR.t1 VPB.t7 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 a_361_297.t0 A1.t0 Y.t4 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 a_193_47.t1 S.t2 VGND.t0 VNB.t6 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 a_361_47.t2 a_27_47.t4 VGND.t4 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 a_193_297.t0 A0.t3 Y.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 Y.t5 A1.t1 a_361_297.t1 VPB.t5 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 Y.t6 A1.t2 a_193_47.t3 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 VGND.t1 S.t3 a_193_47.t0 VNB.t7 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14 VGND.t3 a_27_47.t5 a_361_47.t3 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X15 a_193_47.t2 A1.t3 Y.t7 VNB.t5 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X16 VPWR.t2 S.t4 a_27_47.t0 VPB.t8 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17 VGND.t2 S.t5 a_27_47.t1 VNB.t8 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
R0 A0.n0 A0.t1 212.079
R1 A0.n1 A0.t3 212.079
R2 A0.n0 A0.t2 139.779
R3 A0.n1 A0.t0 139.779
R4 A0.n4 A0.n3 130.626
R5 A0.n6 A0.n2 76
R6 A0.n5 A0.n4 76
R7 A0.n2 A0.n1 32.863
R8 A0.n2 A0.n0 28.481
R9 A0.n6 A0.n5 21.76
R10 A0.n3 A0 18.88
R11 A0.n3 A0 10.56
R12 A0 A0.n6 4.8
R13 A0.n5 A0 2.88
R14 Y.n1 Y.t0 626.232
R15 Y.n2 Y.t5 446.203
R16 Y.n1 Y.n0 292.5
R17 Y.n4 Y.t3 238.823
R18 Y.n5 Y.t6 153.423
R19 Y Y.n5 106.164
R20 Y.n4 Y.n3 92.5
R21 Y.n5 Y.n4 81.317
R22 Y.n2 Y.n1 65.505
R23 Y.n3 Y.t7 32.307
R24 Y.n0 Y.t4 30.535
R25 Y.n0 Y.t1 30.535
R26 Y.n3 Y.t2 24.923
R27 Y Y.n2 22.772
R28 a_361_47.n1 a_361_47.n0 304.129
R29 a_361_47.n0 a_361_47.t3 24.923
R30 a_361_47.n0 a_361_47.t2 24.923
R31 a_361_47.n1 a_361_47.t0 24.923
R32 a_361_47.t1 a_361_47.n1 24.923
R33 VNB VNB.t8 6053.91
R34 VNB.t3 VNB.t1 4545.05
R35 VNB.t0 VNB.t5 2224.18
R36 VNB.t5 VNB.t4 2054.95
R37 VNB.t1 VNB.t0 2030.77
R38 VNB.t2 VNB.t3 2030.77
R39 VNB.t7 VNB.t2 2030.77
R40 VNB.t6 VNB.t7 2030.77
R41 VNB.t8 VNB.t6 2030.77
R42 a_193_297.n1 a_193_297.n0 760.622
R43 a_193_297.n0 a_193_297.t2 26.595
R44 a_193_297.n0 a_193_297.t3 26.595
R45 a_193_297.t1 a_193_297.n1 26.595
R46 a_193_297.n1 a_193_297.t0 26.595
R47 VPB.t2 VPB.t0 556.386
R48 VPB.t1 VPB.t4 272.274
R49 VPB.t4 VPB.t5 251.557
R50 VPB.t0 VPB.t1 248.598
R51 VPB.t3 VPB.t2 248.598
R52 VPB.t6 VPB.t3 248.598
R53 VPB.t7 VPB.t6 248.598
R54 VPB.t8 VPB.t7 248.598
R55 VPB VPB.t8 189.408
R56 a_27_47.t0 a_27_47.n3 579.89
R57 a_27_47.n0 a_27_47.t2 212.079
R58 a_27_47.n1 a_27_47.t3 212.079
R59 a_27_47.n3 a_27_47.n2 202.282
R60 a_27_47.n3 a_27_47.t1 195.685
R61 a_27_47.n0 a_27_47.t5 149.419
R62 a_27_47.n1 a_27_47.t4 149.419
R63 a_27_47.n2 a_27_47.n0 53.02
R64 a_27_47.n2 a_27_47.n1 14.46
R65 a_361_297.n1 a_361_297.n0 764.971
R66 a_361_297.t0 a_361_297.n1 27.58
R67 a_361_297.n0 a_361_297.t3 26.595
R68 a_361_297.n0 a_361_297.t2 26.595
R69 a_361_297.n1 a_361_297.t1 26.595
R70 VPWR.n2 VPWR.t4 584.683
R71 VPWR.n1 VPWR.n0 307.239
R72 VPWR.n6 VPWR.n5 307.239
R73 VPWR.n0 VPWR.t3 26.595
R74 VPWR.n0 VPWR.t0 26.595
R75 VPWR.n5 VPWR.t1 26.595
R76 VPWR.n5 VPWR.t2 26.595
R77 VPWR.n4 VPWR.n3 4.65
R78 VPWR.n2 VPWR.n1 3.951
R79 VPWR.n7 VPWR.n6 3.932
R80 VPWR.n4 VPWR.n2 0.243
R81 VPWR.n7 VPWR.n4 0.137
R82 VPWR VPWR.n7 0.121
R83 S.n0 S.t0 212.079
R84 S.n1 S.t1 212.079
R85 S.n2 S.t4 212.079
R86 S.n0 S.t3 139.779
R87 S.n1 S.t2 139.779
R88 S.n2 S.t5 139.779
R89 S S.n3 79.684
R90 S.n1 S.n0 61.345
R91 S.n3 S.n1 54.772
R92  S 17.435
R93 S.n3 S.n2 6.572
R94 A1.n1 A1.t1 212.079
R95 A1.n0 A1.t0 212.079
R96 A1.n1 A1.t2 139.779
R97 A1.n0 A1.t3 139.779
R98 A1.n2 A1.n1 98.639
R99 A1.n1 A1.n0 62.075
R100 A1.n2 A1 11.224
R101 A1 A1.n2 2.166
R102 VGND.n2 VGND.t3 207.952
R103 VGND.n6 VGND.n5 107.7
R104 VGND.n1 VGND.n0 69.685
R105 VGND.n0 VGND.t4 24.923
R106 VGND.n0 VGND.t1 24.923
R107 VGND.n5 VGND.t0 24.923
R108 VGND.n5 VGND.t2 24.923
R109 VGND.n4 VGND.n3 4.65
R110 VGND.n7 VGND.n6 3.932
R111 VGND.n2 VGND.n1 3.842
R112 VGND.n4 VGND.n2 0.358
R113 VGND.n7 VGND.n4 0.137
R114 VGND VGND.n7 0.121
R115 a_193_47.n1 a_193_47.n0 123.123
R116 a_193_47.t1 a_193_47.n1 27.295
R117 a_193_47.n0 a_193_47.t3 25.846
R118 a_193_47.n0 a_193_47.t2 24.923
R119 a_193_47.n1 a_193_47.t0 21.28
C0 Y VGND 0.33fF
C1 A1 Y 0.10fF
C2 VPWR Y 0.35fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__mux2i_4.ext - technology: sky130A

.subckt sky130_fd_sc_hd__mux2i_4 S A1 A0 Y VGND VPWR VNB VPB
X0 Y.t3 A1.t0 a_445_47.t3 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 Y.t2 A1.t1 a_445_47.t2 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 VPWR.t3 a_1191_21.t2 a_445_297.t7 VPB.t11 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 a_445_297.t3 A1.t2 Y.t5 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 Y.t8 A0.t0 a_109_297.t3 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 a_445_297.t6 a_1191_21.t3 VPWR.t2 VPB.t10 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 a_1191_21.t0 S.t0 VGND.t8 VNB.t14 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 VPWR.t1 a_1191_21.t4 a_445_297.t5 VPB.t9 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 a_445_47.t6 S.t1 VGND.t7 VNB.t15 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 a_109_297.t2 A0.t1 Y.t9 VPB.t5 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 a_445_297.t4 a_1191_21.t5 VPWR.t0 VPB.t8 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 a_445_47.t7 S.t2 VGND.t6 VNB.t16 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 a_109_47.t3 a_1191_21.t6 VGND.t3 VNB.t8 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 Y.t10 A0.t2 a_109_297.t1 VPB.t6 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14 Y.t11 A0.t3 a_109_47.t7 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X15 Y.t12 A0.t4 a_109_47.t6 VNB.t5 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X16 a_1191_21.t1 S.t3 VPWR.t8 VPB.t16 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17 VGND.t5 S.t4 a_445_47.t4 VNB.t12 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X18 Y.t7 A1.t3 a_445_297.t2 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X19 VGND.t4 S.t5 a_445_47.t5 VNB.t13 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X20 VGND.t2 a_1191_21.t7 a_109_47.t2 VNB.t9 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X21 a_109_47.t5 A0.t5 Y.t13 VNB.t6 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X22 a_445_47.t1 A1.t4 Y.t1 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X23 a_445_297.t1 A1.t5 Y.t6 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X24 VPWR.t4 S.t6 a_109_297.t4 VPB.t12 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X25 a_445_47.t0 A1.t6 Y.t0 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X26 VGND.t1 a_1191_21.t8 a_109_47.t1 VNB.t10 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X27 Y.t4 A1.t7 a_445_297.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X28 a_109_297.t5 S.t7 VPWR.t5 VPB.t13 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X29 VPWR.t6 S.t8 a_109_297.t6 VPB.t14 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X30 a_109_47.t0 a_1191_21.t9 VGND.t0 VNB.t11 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X31 a_109_297.t0 A0.t6 Y.t14 VPB.t7 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X32 a_109_297.t7 S.t9 VPWR.t7 VPB.t15 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X33 a_109_47.t4 A0.t7 Y.t15 VNB.t7 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
R0 A1.n0 A1.t3 212.079
R1 A1.n2 A1.t5 212.079
R2 A1.n3 A1.t7 212.079
R3 A1.n4 A1.t2 212.079
R4 A1.n0 A1.t1 139.779
R5 A1.n2 A1.t6 139.779
R6 A1.n3 A1.t0 139.779
R7 A1.n4 A1.t4 139.779
R8 A1.n11 A1.n1 76
R9 A1.n10 A1.n9 76
R10 A1.n8 A1.n7 76
R11 A1.n6 A1.n5 76
R12 A1.n9 A1.n8 49.66
R13 A1.n5 A1.n3 48.2
R14 A1.n1 A1.n0 21.909
R15 A1.n11 A1.n10 13.187
R16 A1.n5 A1.n4 13.145
R17 A1.n7 A1 12.8
R18 A1.n9 A1.n2 10.224
R19 A1.n6 A1 9.696
R20 A1 A1.n6 8.145
R21 A1.n7 A1 5.042
R22 A1 A1.n11 4.266
R23 A1.n8 A1.n3 1.46
R24 A1.n10 A1 0.387
R25 a_445_47.n2 a_445_47.n1 173.441
R26 a_445_47.n4 a_445_47.n3 155.747
R27 a_445_47.n2 a_445_47.n0 110.194
R28 a_445_47.n4 a_445_47.n2 102.4
R29 a_445_47.n5 a_445_47.n4 92.5
R30 a_445_47.n3 a_445_47.t3 24.923
R31 a_445_47.n3 a_445_47.t1 24.923
R32 a_445_47.n0 a_445_47.t5 24.923
R33 a_445_47.n0 a_445_47.t7 24.923
R34 a_445_47.n1 a_445_47.t4 24.923
R35 a_445_47.n1 a_445_47.t6 24.923
R36 a_445_47.n5 a_445_47.t2 24.923
R37 a_445_47.t0 a_445_47.n5 24.923
R38 Y.n1 Y.t7 624.727
R39 Y.n6 Y.t14 561.48
R40 Y.n1 Y.n0 292.5
R41 Y.n3 Y.n2 292.5
R42 Y.n5 Y.n4 292.5
R43 Y.n8 Y.t2 229.593
R44 Y.n13 Y.t15 166.346
R45 Y.n8 Y.n7 92.5
R46 Y.n10 Y.n9 92.5
R47 Y.n12 Y.n11 92.5
R48 Y.n3 Y.n1 63.247
R49 Y.n5 Y.n3 63.247
R50 Y.n10 Y.n8 63.247
R51 Y.n12 Y.n10 63.247
R52 Y.n6 Y.n5 58.729
R53 Y.n13 Y.n12 58.729
R54 Y.n4 Y.t9 26.595
R55 Y.n4 Y.t10 26.595
R56 Y.n2 Y.t5 26.595
R57 Y.n2 Y.t8 26.595
R58 Y.n0 Y.t6 26.595
R59 Y.n0 Y.t4 26.595
R60 Y.n11 Y.t13 24.923
R61 Y.n11 Y.t11 24.923
R62 Y.n9 Y.t1 24.923
R63 Y.n9 Y.t12 24.923
R64 Y.n7 Y.t0 24.923
R65 Y.n7 Y.t3 24.923
R66 Y Y.n13 20.764
R67 Y Y.n6 12.231
R68 VNB VNB.t7 6053.91
R69 VNB.t2 VNB.t16 4545.05
R70 VNB.t11 VNB.t10 2296.7
R71 VNB.t10 VNB.t14 2248.35
R72 VNB.t9 VNB.t11 2030.77
R73 VNB.t8 VNB.t9 2030.77
R74 VNB.t12 VNB.t8 2030.77
R75 VNB.t15 VNB.t12 2030.77
R76 VNB.t13 VNB.t15 2030.77
R77 VNB.t16 VNB.t13 2030.77
R78 VNB.t0 VNB.t2 2030.77
R79 VNB.t3 VNB.t0 2030.77
R80 VNB.t1 VNB.t3 2030.77
R81 VNB.t5 VNB.t1 2030.77
R82 VNB.t6 VNB.t5 2030.77
R83 VNB.t4 VNB.t6 2030.77
R84 VNB.t7 VNB.t4 2030.77
R85 a_1191_21.t1 a_1191_21.n5 260.17
R86 a_1191_21.n3 a_1191_21.t2 212.079
R87 a_1191_21.n2 a_1191_21.t3 212.079
R88 a_1191_21.n1 a_1191_21.t4 212.079
R89 a_1191_21.n0 a_1191_21.t5 212.079
R90 a_1191_21.n5 a_1191_21.t0 172.868
R91 a_1191_21.n3 a_1191_21.t8 139.779
R92 a_1191_21.n2 a_1191_21.t9 139.779
R93 a_1191_21.n1 a_1191_21.t7 139.779
R94 a_1191_21.n0 a_1191_21.t6 139.779
R95 a_1191_21.n5 a_1191_21.n4 103.845
R96 a_1191_21.n2 a_1191_21.n1 61.345
R97 a_1191_21.n1 a_1191_21.n0 61.345
R98 a_1191_21.n4 a_1191_21.n3 30.394
R99 a_1191_21.n4 a_1191_21.n2 27.051
R100 a_445_297.n5 a_445_297.n4 355.747
R101 a_445_297.n4 a_445_297.n3 292.5
R102 a_445_297.n4 a_445_297.n2 228.894
R103 a_445_297.n2 a_445_297.n0 213.435
R104 a_445_297.n2 a_445_297.n1 150.188
R105 a_445_297.n0 a_445_297.t7 37.43
R106 a_445_297.n3 a_445_297.t2 26.595
R107 a_445_297.n3 a_445_297.t1 26.595
R108 a_445_297.n1 a_445_297.t5 26.595
R109 a_445_297.n1 a_445_297.t4 26.595
R110 a_445_297.n0 a_445_297.t6 26.595
R111 a_445_297.n5 a_445_297.t0 26.595
R112 a_445_297.t3 a_445_297.n5 26.595
R113 VPWR.n0 VPWR.t7 576.219
R114 VPWR.n4 VPWR.n3 310.785
R115 VPWR.n2 VPWR.n1 307.239
R116 VPWR.n8 VPWR.n7 307.239
R117 VPWR.n13 VPWR.n12 307.239
R118 VPWR.n3 VPWR.t3 35.46
R119 VPWR.n3 VPWR.t8 26.595
R120 VPWR.n1 VPWR.t2 26.595
R121 VPWR.n1 VPWR.t1 26.595
R122 VPWR.n7 VPWR.t0 26.595
R123 VPWR.n7 VPWR.t4 26.595
R124 VPWR.n12 VPWR.t5 26.595
R125 VPWR.n12 VPWR.t6 26.595
R126 VPWR.n17 VPWR.n0 9.034
R127 VPWR.n16 VPWR.n15 4.65
R128 VPWR.n6 VPWR.n5 4.65
R129 VPWR.n9 VPWR.n8 4.65
R130 VPWR.n11 VPWR.n10 4.65
R131 VPWR.n14 VPWR.n13 4.65
R132 VPWR.n4 VPWR.n2 3.863
R133 VPWR VPWR.n17 0.962
R134 VPWR.n6 VPWR.n4 0.225
R135 VPWR.n17 VPWR.n16 0.134
R136 VPWR.n9 VPWR.n6 0.119
R137 VPWR.n11 VPWR.n9 0.119
R138 VPWR.n14 VPWR.n11 0.119
R139 VPWR.n16 VPWR.n14 0.119
R140 VPB.t2 VPB.t15 556.386
R141 VPB.t10 VPB.t11 281.152
R142 VPB.t11 VPB.t16 275.233
R143 VPB.t9 VPB.t10 248.598
R144 VPB.t8 VPB.t9 248.598
R145 VPB.t12 VPB.t8 248.598
R146 VPB.t13 VPB.t12 248.598
R147 VPB.t14 VPB.t13 248.598
R148 VPB.t15 VPB.t14 248.598
R149 VPB.t1 VPB.t2 248.598
R150 VPB.t0 VPB.t1 248.598
R151 VPB.t3 VPB.t0 248.598
R152 VPB.t4 VPB.t3 248.598
R153 VPB.t5 VPB.t4 248.598
R154 VPB.t6 VPB.t5 248.598
R155 VPB.t7 VPB.t6 248.598
R156 VPB VPB.t7 189.408
R157 A0.n0 A0.t0 212.079
R158 A0.n1 A0.t1 212.079
R159 A0.n2 A0.t2 212.079
R160 A0.n5 A0.t6 212.079
R161 A0.n0 A0.t4 139.779
R162 A0.n1 A0.t5 139.779
R163 A0.n2 A0.t3 139.779
R164 A0.n5 A0.t7 139.779
R165 A0.n4 A0.n3 76
R166 A0.n7 A0.n6 76
R167 A0.n1 A0.n0 61.345
R168 A0.n3 A0.n1 47.469
R169 A0.n6 A0.n5 25.56
R170 A0.n3 A0.n2 13.875
R171 A0.n7 A0.n4 13.187
R172 A0.n4 A0 11.578
R173 A0 A0.n7 1.357
R174 a_109_297.n4 a_109_297.n3 355.747
R175 a_109_297.n2 a_109_297.n0 355.747
R176 a_109_297.n2 a_109_297.n1 292.5
R177 a_109_297.n5 a_109_297.n4 292.5
R178 a_109_297.n4 a_109_297.n2 228.894
R179 a_109_297.n3 a_109_297.t1 26.595
R180 a_109_297.n3 a_109_297.t0 26.595
R181 a_109_297.n1 a_109_297.t6 26.595
R182 a_109_297.n1 a_109_297.t7 26.595
R183 a_109_297.n0 a_109_297.t4 26.595
R184 a_109_297.n0 a_109_297.t5 26.595
R185 a_109_297.t3 a_109_297.n5 26.595
R186 a_109_297.n5 a_109_297.t2 26.595
R187 S S.n0 259.907
R188 S.n0 S.t3 241.534
R189 S.n1 S.t6 212.079
R190 S.n4 S.t7 212.079
R191 S.n9 S.t8 212.079
R192 S.n5 S.t9 212.079
R193 S.n0 S.t0 169.234
R194 S.n1 S.t4 139.779
R195 S.n4 S.t1 139.779
R196 S.n9 S.t5 139.779
R197 S.n5 S.t2 139.779
R198 S.n6 S.n5 103.751
R199 S.n13 S.n2 76
R200 S.n12 S.n11 76
R201 S.n8 S.n7 76
R202 S.n11 S.n10 49.66
R203 S.n4 S.n2 48.2
R204 S.n9 S.n8 39.436
R205 S.n8 S.n5 21.909
R206 S.n12 S.n3 20.241
R207 S.n6 S 18.455
R208 S.n13 S 17.265
R209 S.n7 S 16.074
R210 S.n2 S.n1 13.145
R211 S.n7 S 11.311
R212 S.n10 S.n9 10.224
R213 S S.n13 10.12
R214 S S.n6 8.93
R215 S S.n3 4.167
R216 S S.n12 2.976
R217 S.n11 S.n4 1.46
R218 VGND.n0 VGND.t6 190.315
R219 VGND.n3 VGND.n2 111.956
R220 VGND.n4 VGND.n1 110.793
R221 VGND.n8 VGND.n7 109.238
R222 VGND.n13 VGND.n12 107.239
R223 VGND.n1 VGND.t1 33.23
R224 VGND.n1 VGND.t8 24.923
R225 VGND.n2 VGND.t0 24.923
R226 VGND.n2 VGND.t2 24.923
R227 VGND.n7 VGND.t3 24.923
R228 VGND.n7 VGND.t5 24.923
R229 VGND.n12 VGND.t7 24.923
R230 VGND.n12 VGND.t4 24.923
R231 VGND.n17 VGND.n0 9.034
R232 VGND.n6 VGND.n5 4.65
R233 VGND.n9 VGND.n8 4.65
R234 VGND.n11 VGND.n10 4.65
R235 VGND.n14 VGND.n13 4.65
R236 VGND.n16 VGND.n15 4.65
R237 VGND.n4 VGND.n3 3.916
R238 VGND VGND.n17 0.962
R239 VGND.n6 VGND.n4 0.218
R240 VGND.n17 VGND.n16 0.134
R241 VGND.n9 VGND.n6 0.119
R242 VGND.n11 VGND.n9 0.119
R243 VGND.n14 VGND.n11 0.119
R244 VGND.n16 VGND.n14 0.119
R245 a_109_47.n8 a_109_47.n0 150.462
R246 a_109_47.n2 a_109_47.n1 149.037
R247 a_109_47.n9 a_109_47.n8 114.077
R248 a_109_47.n0 a_109_47.t1 35.076
R249 a_109_47.n1 a_109_47.t7 24.923
R250 a_109_47.n1 a_109_47.t4 24.923
R251 a_109_47.n0 a_109_47.t0 24.923
R252 a_109_47.n9 a_109_47.t2 24.923
R253 a_109_47.t3 a_109_47.n9 24.923
R254 a_109_47.n4 a_109_47.t5 17.538
R255 a_109_47.n6 a_109_47.t6 16.615
R256 a_109_47.n8 a_109_47.n7 12.146
R257 a_109_47.n7 a_109_47.n6 9.3
R258 a_109_47.n6 a_109_47.n5 8.307
R259 a_109_47.n5 a_109_47.n4 7.384
R260 a_109_47.n7 a_109_47.n3 2.057
R261 a_109_47.n3 a_109_47.n2 1.828
C0 VPB VPWR 0.16fF
C1 Y VPWR 0.54fF
C2 Y VGND 0.50fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__mux4_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__mux4_1 S0 A1 X S1 A2 A0 A3 VGND VPWR VNB VPB
X0 a_277_47.t4 a_247_21.t2 a_27_413.t1 VPB.t12 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1 VGND.t6 S0.t0 a_247_21.t1 VNB.t12 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 a_834_97.t1 a_247_21.t3 a_750_97.t2 VNB.t9 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3 VGND.t0 A3.t0 a_668_97.t0 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 a_1290_413.t1 S1.t0 VPWR.t1 VPB.t8 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 a_834_97.t0 A2.t0 VGND.t1 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 a_750_97.t5 S0.t1 a_757_363.t1 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7 a_27_47.t1 S0.t2 a_277_47.t1 VNB.t11 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 X.t0 a_1478_413.t4 VGND.t4 VNB.t5 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 VPWR.t5 A1.t0 a_27_413.t0 VPB.t10 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10 VPWR.t6 S0.t3 a_247_21.t0 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11 X.t1 a_1478_413.t5 VPWR.t3 VPB.t7 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 a_193_47.t0 A0.t0 VGND.t2 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13 a_750_97.t0 a_1290_413.t2 a_1478_413.t1 VPB.t5 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14 a_1478_413.t2 S1.t1 a_277_47.t3 VPB.t9 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15 a_1290_413.t0 S1.t2 VGND.t5 VNB.t7 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16 a_277_47.t5 a_247_21.t4 a_193_47.t1 VNB.t8 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17 a_750_97.t4 S0.t4 a_668_97.t1 VNB.t10 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18 a_923_363.t1 a_247_21.t5 a_750_97.t3 VPB.t11 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19 a_757_363.t0 A2.t1 VPWR.t0 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20 VPWR.t4 A3.t1 a_923_363.t0 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21 a_277_47.t2 a_1290_413.t3 a_1478_413.t0 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22 a_193_413.t0 A0.t1 VPWR.t2 VPB.t6 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23 a_193_413.t1 S0.t5 a_277_47.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24 VGND.t3 A1.t1 a_27_47.t0 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X25 a_1478_413.t3 S1.t3 a_750_97.t1 VNB.t6 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
R0 a_247_21.n1 a_247_21.t4 404.879
R1 a_247_21.n3 a_247_21.n0 343.846
R2 a_247_21.n2 a_247_21.t5 287.023
R3 a_247_21.n1 a_247_21.t2 221.72
R4 a_247_21.n0 a_247_21.n1 186.854
R5 a_247_21.n0 a_247_21.t1 152.226
R6 a_247_21.n2 a_247_21.t3 145.091
R7 a_247_21.n3 a_247_21.t0 41.708
R8 a_247_21.n4 a_247_21.n3 35.46
R9 a_247_21.n0 a_247_21.n2 17.628
R10 a_27_413.t0 a_27_413.t1 839.265
R11 a_277_47.n0 a_277_47.t3 465.413
R12 a_277_47.n3 a_277_47.n2 398.557
R13 a_277_47.n0 a_277_47.t2 151.497
R14 a_277_47.n2 a_277_47.n1 103.532
R15 a_277_47.n1 a_277_47.t5 74.114
R16 a_277_47.t0 a_277_47.n3 63.321
R17 a_277_47.n3 a_277_47.t4 63.321
R18 a_277_47.n1 a_277_47.t1 37.143
R19 a_277_47.n2 a_277_47.n0 9.475
R20 VPB.t5 VPB.t7 822.741
R21 VPB.t8 VPB.t9 556.386
R22 VPB.t4 VPB.t8 556.386
R23 VPB.t0 VPB.t1 556.386
R24 VPB.t6 VPB.t12 556.386
R25 VPB.t1 VPB.t2 550.467
R26 VPB.t9 VPB.t5 287.071
R27 VPB.t11 VPB.t3 281.152
R28 VPB.t3 VPB.t4 248.598
R29 VPB.t2 VPB.t11 248.598
R30 VPB.t12 VPB.t0 248.598
R31 VPB.t10 VPB.t6 248.598
R32 VPB VPB.t10 192.367
R33 S0.t0 S0.t2 547.873
R34 S0.n0 S0.t1 377.24
R35 S0.n1 S0.t5 223.326
R36 S0.n0 S0.t3 173.996
R37 S0.n3 S0.t4 130.27
R38 S0.n2 S0.t0 123.428
R39 S0 S0.n3 87.306
R40 S0.n2 S0.n1 41.375
R41 S0.n3 S0.n2 24.751
R42  S0 14.506
R43 S0.n1 S0.n0 1.784
R44 VGND.n1 VGND.t4 202.815
R45 VGND.n16 VGND.t6 159.319
R46 VGND.n0 VGND.t5 145.81
R47 VGND.n5 VGND.n4 114.711
R48 VGND.n27 VGND.n26 107.239
R49 VGND.n4 VGND.t1 38.571
R50 VGND.n4 VGND.t0 38.571
R51 VGND.n26 VGND.t2 38.571
R52 VGND.n26 VGND.t3 38.571
R53 VGND.n3 VGND.n2 4.65
R54 VGND.n7 VGND.n6 4.65
R55 VGND.n9 VGND.n8 4.65
R56 VGND.n11 VGND.n10 4.65
R57 VGND.n13 VGND.n12 4.65
R58 VGND.n15 VGND.n14 4.65
R59 VGND.n17 VGND.n16 4.65
R60 VGND.n19 VGND.n18 4.65
R61 VGND.n21 VGND.n20 4.65
R62 VGND.n23 VGND.n22 4.65
R63 VGND.n25 VGND.n24 4.65
R64 VGND.n6 VGND.n5 4.141
R65 VGND.n1 VGND.n0 3.992
R66 VGND.n28 VGND.n27 3.932
R67 VGND.n3 VGND.n1 0.138
R68 VGND.n28 VGND.n25 0.137
R69 VGND VGND.n28 0.123
R70 VGND.n7 VGND.n3 0.119
R71 VGND.n9 VGND.n7 0.119
R72 VGND.n11 VGND.n9 0.119
R73 VGND.n13 VGND.n11 0.119
R74 VGND.n15 VGND.n13 0.119
R75 VGND.n17 VGND.n15 0.119
R76 VGND.n19 VGND.n17 0.119
R77 VGND.n21 VGND.n19 0.119
R78 VGND.n23 VGND.n21 0.119
R79 VGND.n25 VGND.n23 0.119
R80 VNB VNB.t4 6470.59
R81 VNB.t11 VNB.t12 6086.94
R82 VNB.t12 VNB.t10 6085.86
R83 VNB.t7 VNB.t6 6082.35
R84 VNB.t1 VNB.t7 6082.35
R85 VNB.t9 VNB.t0 6017.65
R86 VNB.t2 VNB.t5 5270.33
R87 VNB.t6 VNB.t2 4158.57
R88 VNB.t0 VNB.t1 2717.65
R89 VNB.t10 VNB.t9 2717.65
R90 VNB.t3 VNB.t8 2717.65
R91 VNB.t4 VNB.t3 2717.65
R92 VNB.t8 VNB.t11 2395.55
R93 a_750_97.t0 a_750_97.n3 373.822
R94 a_750_97.n2 a_750_97.n0 299.093
R95 a_750_97.n3 a_750_97.t1 255.452
R96 a_750_97.n2 a_750_97.n1 177.693
R97 a_750_97.n0 a_750_97.t3 63.321
R98 a_750_97.n0 a_750_97.t5 63.321
R99 a_750_97.n1 a_750_97.t2 38.571
R100 a_750_97.n1 a_750_97.t4 38.571
R101 a_750_97.n3 a_750_97.n2 12.081
R102 a_834_97.t0 a_834_97.t1 370.715
R103 A3.n0 A3.t1 310.456
R104 A3.n0 A3.t0 220.483
R105 A3.n1 A3.n0 76
R106  A3.n1 11.755
R107 A3.n1 A3 6.008
R108 a_668_97.n0 a_668_97.t1 337.927
R109 a_668_97.n0 a_668_97.t0 30
R110 S1.n1 S1.t0 322.745
R111 S1.n0 S1.t1 305.266
R112 S1.n1 S1.t2 194.212
R113 S1.n0 S1.t3 179.823
R114 S1.n1 S1.n0 126.803
R115 S1 S1.n1 78.427
R116 VPWR.n1 VPWR.t3 580.338
R117 VPWR.n13 VPWR.t6 372.663
R118 VPWR.n0 VPWR.t1 369.718
R119 VPWR.n5 VPWR.n4 307.239
R120 VPWR.n26 VPWR.n25 307.239
R121 VPWR.n4 VPWR.t0 63.321
R122 VPWR.n4 VPWR.t4 63.321
R123 VPWR.n25 VPWR.t2 63.321
R124 VPWR.n25 VPWR.t5 63.321
R125 VPWR.n3 VPWR.n2 4.65
R126 VPWR.n6 VPWR.n5 4.65
R127 VPWR.n8 VPWR.n7 4.65
R128 VPWR.n10 VPWR.n9 4.65
R129 VPWR.n12 VPWR.n11 4.65
R130 VPWR.n14 VPWR.n13 4.65
R131 VPWR.n16 VPWR.n15 4.65
R132 VPWR.n18 VPWR.n17 4.65
R133 VPWR.n20 VPWR.n19 4.65
R134 VPWR.n22 VPWR.n21 4.65
R135 VPWR.n24 VPWR.n23 4.65
R136 VPWR.n1 VPWR.n0 4.006
R137 VPWR.n27 VPWR.n26 3.932
R138 VPWR.n3 VPWR.n1 0.138
R139 VPWR.n27 VPWR.n24 0.137
R140 VPWR VPWR.n27 0.123
R141 VPWR.n6 VPWR.n3 0.119
R142 VPWR.n8 VPWR.n6 0.119
R143 VPWR.n10 VPWR.n8 0.119
R144 VPWR.n12 VPWR.n10 0.119
R145 VPWR.n14 VPWR.n12 0.119
R146 VPWR.n16 VPWR.n14 0.119
R147 VPWR.n18 VPWR.n16 0.119
R148 VPWR.n20 VPWR.n18 0.119
R149 VPWR.n22 VPWR.n20 0.119
R150 VPWR.n24 VPWR.n22 0.119
R151 a_1290_413.n1 a_1290_413.t1 435.74
R152 a_1290_413.n0 a_1290_413.t2 312.227
R153 a_1290_413.t0 a_1290_413.n1 180.772
R154 a_1290_413.n1 a_1290_413.n0 149.581
R155 a_1290_413.n0 a_1290_413.t3 115.68
R156 A2.n0 A2.t1 315.441
R157 A2.n0 A2.t0 225.468
R158 A2 A2.n0 80.335
R159 a_757_363.t0 a_757_363.t1 901.602
R160 a_27_47.t0 a_27_47.t1 434.563
R161 a_1478_413.n2 a_1478_413.n0 481.052
R162 a_1478_413.n1 a_1478_413.t5 233.573
R163 a_1478_413.n3 a_1478_413.n2 227.274
R164 a_1478_413.n1 a_1478_413.t4 161.273
R165 a_1478_413.n0 a_1478_413.t1 140.84
R166 a_1478_413.t0 a_1478_413.n3 121.849
R167 a_1478_413.n3 a_1478_413.t3 118.571
R168 a_1478_413.n2 a_1478_413.n1 76
R169 a_1478_413.n0 a_1478_413.t2 60.976
R170 X X.t1 556.526
R171 X X.t0 174.099
R172 A1.n0 A1.t0 334.721
R173 A1.n0 A1.t1 206.188
R174 A1.n1 A1.n0 76
R175 A1.n1 A1 10.573
R176 A1 A1.n1 2.04
R177 A0.n0 A0.t1 334.721
R178 A0.n0 A0.t0 206.188
R179 A0.n1 A0.n0 76
R180 A0.n1 A0 8.386
R181 A0 A0.n1 1.618
R182 a_193_47.t0 a_193_47.t1 77.142
R183 a_923_363.t0 a_923_363.t1 204.173
R184 a_193_413.t0 a_193_413.t1 841.368
C0 VPB S0 0.11fF
C1 A3 A2 0.20fF
C2 VPB VPWR 0.20fF
C3 A1 A0 0.17fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__mux4_2.ext - technology: sky130A

.subckt sky130_fd_sc_hd__mux4_2 VGND VPWR X S0 A2 A3 S1 A1 A0 VNB VPB
X0 a_600_345.t1 S1.t0 VPWR.t6 VPB.t12 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1 a_788_316.t2 S1.t1 a_288_47.t5 VNB.t13 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 VPWR.t2 A3.t0 a_372_413.t1 VPB.t5 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X3 a_872_316.t2 a_600_345.t2 a_788_316.t1 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 VPWR.t0 S0.t0 a_27_47.t1 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X5 a_1279_413.t0 S0.t1 a_872_316.t0 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 VGND.t3 a_788_316.t4 X.t1 VNB.t9 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 a_1060_369.t0 A1.t0 VPWR.t1 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X8 a_872_316.t4 a_27_47.t2 a_1060_369.t1 VPB.t7 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9 a_1281_47.t1 a_27_47.t3 a_872_316.t3 VNB.t6 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X10 a_193_47.t1 A2.t0 VGND.t5 VNB.t11 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11 a_1064_47.t1 A1.t1 VGND.t0 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12 a_872_316.t5 S1.t2 a_788_316.t3 VPB.t11 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=540000u l=150000u
X13 a_872_316.t1 S0.t2 a_1064_47.t0 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X14 X.t0 a_788_316.t5 VGND.t2 VNB.t8 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X15 a_788_316.t0 a_600_345.t3 a_288_47.t2 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=540000u l=150000u
X16 a_372_413.t0 a_27_47.t4 a_288_47.t3 VPB.t6 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17 VGND.t7 A3.t1 a_397_47.t1 VNB.t5 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18 a_600_345.t0 S1.t3 VGND.t6 VNB.t12 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19 a_193_369.t1 A2.t1 VPWR.t5 VPB.t10 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X20 VPWR.t3 a_788_316.t6 X.t3 VPB.t8 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X21 a_288_47.t0 S0.t3 a_193_369.t0 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22 a_397_47.t0 S0.t4 a_288_47.t1 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X23 VGND.t4 A0.t0 a_1281_47.t0 VNB.t10 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24 a_288_47.t4 a_27_47.t5 a_193_47.t0 VNB.t7 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X25 X.t2 a_788_316.t7 VPWR.t4 VPB.t9 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X26 VGND.t1 S0.t5 a_27_47.t0 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X27 VPWR.t7 A0.t1 a_1279_413.t1 VPB.t13 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
R0 S1.t0 S1.t2 769.592
R1 S1.n0 S1.t1 367.926
R2 S1.n1 S1.t0 350.711
R3 S1.n0 S1.t3 112.237
R4 S1.n2 S1.n1 76
R5 S1.n1 S1.n0 34.428
R6 S1.n2 S1 7.724
R7 S1 S1.n2 7.282
R8 VPWR.n11 VPWR.t1 351.862
R9 VPWR.n22 VPWR.n21 320.326
R10 VPWR.n32 VPWR.n31 307.239
R11 VPWR.n1 VPWR.n0 174.594
R12 VPWR.n2 VPWR.t3 172.632
R13 VPWR.n0 VPWR.t7 61.562
R14 VPWR.n21 VPWR.t6 41.554
R15 VPWR.n21 VPWR.t2 41.554
R16 VPWR.n31 VPWR.t5 41.554
R17 VPWR.n31 VPWR.t0 41.554
R18 VPWR.n0 VPWR.t4 30.594
R19 VPWR.n2 VPWR.n1 6.331
R20 VPWR.n23 VPWR.n22 4.894
R21 VPWR.n4 VPWR.n3 4.65
R22 VPWR.n6 VPWR.n5 4.65
R23 VPWR.n8 VPWR.n7 4.65
R24 VPWR.n10 VPWR.n9 4.65
R25 VPWR.n12 VPWR.n11 4.65
R26 VPWR.n14 VPWR.n13 4.65
R27 VPWR.n16 VPWR.n15 4.65
R28 VPWR.n18 VPWR.n17 4.65
R29 VPWR.n20 VPWR.n19 4.65
R30 VPWR.n24 VPWR.n23 4.65
R31 VPWR.n26 VPWR.n25 4.65
R32 VPWR.n28 VPWR.n27 4.65
R33 VPWR.n30 VPWR.n29 4.65
R34 VPWR.n33 VPWR.n32 3.932
R35 VPWR.n4 VPWR.n2 0.2
R36 VPWR.n33 VPWR.n30 0.137
R37 VPWR VPWR.n33 0.123
R38 VPWR.n6 VPWR.n4 0.119
R39 VPWR.n8 VPWR.n6 0.119
R40 VPWR.n10 VPWR.n8 0.119
R41 VPWR.n12 VPWR.n10 0.119
R42 VPWR.n14 VPWR.n12 0.119
R43 VPWR.n16 VPWR.n14 0.119
R44 VPWR.n18 VPWR.n16 0.119
R45 VPWR.n20 VPWR.n18 0.119
R46 VPWR.n24 VPWR.n20 0.119
R47 VPWR.n26 VPWR.n24 0.119
R48 VPWR.n28 VPWR.n26 0.119
R49 VPWR.n30 VPWR.n28 0.119
R50 a_600_345.t1 a_600_345.n1 466.234
R51 a_600_345.n0 a_600_345.t2 337.934
R52 a_600_345.n1 a_600_345.t0 201.267
R53 a_600_345.n1 a_600_345.n0 159.903
R54 a_600_345.n0 a_600_345.t3 157.453
R55 VPB.t11 VPB.t3 556.386
R56 VPB.t12 VPB.t4 556.386
R57 VPB.t6 VPB.t5 426.168
R58 VPB.t3 VPB.t7 399.532
R59 VPB.t1 VPB.t13 298.909
R60 VPB.t13 VPB.t9 287.071
R61 VPB.t10 VPB.t2 281.152
R62 VPB.t9 VPB.t8 248.598
R63 VPB.t7 VPB.t1 248.598
R64 VPB.t4 VPB.t11 248.598
R65 VPB.t5 VPB.t12 248.598
R66 VPB.t2 VPB.t6 248.598
R67 VPB.t0 VPB.t10 248.598
R68 VPB VPB.t0 192.367
R69 a_288_47.t2 a_288_47.n3 341.75
R70 a_288_47.n2 a_288_47.n1 329.77
R71 a_288_47.n2 a_288_47.n0 244.968
R72 a_288_47.n3 a_288_47.t5 233.798
R73 a_288_47.n0 a_288_47.t1 66.666
R74 a_288_47.n0 a_288_47.t4 65
R75 a_288_47.n1 a_288_47.t3 63.321
R76 a_288_47.n1 a_288_47.t0 63.321
R77 a_288_47.n3 a_288_47.n2 30.883
R78 a_788_316.n5 a_788_316.n4 292.5
R79 a_788_316.n4 a_788_316.n2 228.38
R80 a_788_316.n0 a_788_316.t6 212.079
R81 a_788_316.n1 a_788_316.t7 212.079
R82 a_788_316.n4 a_788_316.n3 174.352
R83 a_788_316.n0 a_788_316.t4 139.779
R84 a_788_316.n1 a_788_316.t5 139.779
R85 a_788_316.n2 a_788_316.n0 56.963
R86 a_788_316.n5 a_788_316.t3 49.25
R87 a_788_316.t0 a_788_316.n5 49.25
R88 a_788_316.n3 a_788_316.t2 40
R89 a_788_316.n3 a_788_316.t1 38.571
R90 a_788_316.n2 a_788_316.n1 4.381
R91 VNB VNB.t2 6470.59
R92 VNB.t12 VNB.t13 6147.06
R93 VNB.t4 VNB.t3 6082.35
R94 VNB.t0 VNB.t6 3558.82
R95 VNB.t7 VNB.t1 3526.47
R96 VNB.t5 VNB.t12 3494.12
R97 VNB.t3 VNB.t0 3461.76
R98 VNB.t1 VNB.t5 3105.88
R99 VNB.t6 VNB.t10 3073.53
R100 VNB.t11 VNB.t7 3073.53
R101 VNB.t13 VNB.t4 2750
R102 VNB.t2 VNB.t11 2717.65
R103 VNB.t10 VNB.t8 2400.4
R104 VNB.t8 VNB.t9 2030.77
R105 A3.n0 A3.t0 313.804
R106 A3.n0 A3.t1 132.281
R107 A3.n1 A3.n0 76
R108 A3 A3.n1 8.52
R109 A3.n1 A3 5.632
R110 a_372_413.t1 a_372_413.t0 245.006
R111 a_372_413.n0 a_372_413.t1 101.896
R112 a_872_316.n2 a_872_316.n0 376.828
R113 a_872_316.t5 a_872_316.n3 347.139
R114 a_872_316.n2 a_872_316.n1 223.887
R115 a_872_316.n3 a_872_316.t2 220.887
R116 a_872_316.n1 a_872_316.t3 66.666
R117 a_872_316.n1 a_872_316.t1 66.666
R118 a_872_316.n0 a_872_316.t0 63.321
R119 a_872_316.n0 a_872_316.t4 63.321
R120 a_872_316.n3 a_872_316.n2 62.117
R121 S0.n1 S0.t4 445.045
R122 S0.n5 S0.t2 432.192
R123 S0.n7 S0.t0 287.994
R124 S0.n2 S0.t3 258.42
R125 S0.n5 S0.t1 254.388
R126 S0.n7 S0.t5 194.808
R127 S0.n6 S0.n5 90.486
R128 S0.n8 S0.n7 76
R129 S0 S0.n8 20.266
R130 S0.n4 S0.n3 18.793
R131 S0.n3 S0.n1 14.46
R132 S0 S0.n6 11.432
R133 S0.n3 S0.n2 6.159
R134 S0.n4 S0.n0 6.023
R135 S0.n6 S0.n4 4.518
R136 S0.n8 S0 3.911
R137 a_27_47.t1 a_27_47.n3 370.947
R138 a_27_47.n0 a_27_47.t5 246.293
R139 a_27_47.n3 a_27_47.t0 244.313
R140 a_27_47.n1 a_27_47.t3 241.28
R141 a_27_47.n0 a_27_47.t4 224.251
R142 a_27_47.n1 a_27_47.t2 146.443
R143 a_27_47.n3 a_27_47.n2 67.388
R144 a_27_47.n2 a_27_47.n1 11.44
R145 a_27_47.n2 a_27_47.n0 4.894
R146 a_1279_413.n0 a_1279_413.t0 100.845
R147 a_1279_413.n1 a_1279_413.n0 77.392
R148 a_1279_413.n0 a_1279_413.t1 33.965
R149 X.n1 X.n0 145.944
R150 X.n4 X.n3 92.5
R151 X.n4 X 81.392
R152 X.n0 X.t3 26.595
R153 X.n0 X.t2 26.595
R154 X.n3 X.t1 24.923
R155 X.n3 X.t0 24.923
R156 X.n2 X.n1 5.792
R157 X.n1 X 3.194
R158 X X.n2 2.064
R159 X.n2 X 1.56
R160 X X.n4 0.193
R161 VGND.n11 VGND.t0 145.81
R162 VGND.n1 VGND.n0 119.1
R163 VGND.n2 VGND.t3 113.05
R164 VGND.n22 VGND.n21 107.239
R165 VGND.n31 VGND.n30 107.239
R166 VGND.n0 VGND.t4 62.351
R167 VGND.n21 VGND.t6 57.142
R168 VGND.n21 VGND.t7 54.285
R169 VGND.n30 VGND.t5 38.571
R170 VGND.n30 VGND.t1 38.571
R171 VGND.n0 VGND.t2 24.924
R172 VGND.n4 VGND.n3 4.65
R173 VGND.n6 VGND.n5 4.65
R174 VGND.n8 VGND.n7 4.65
R175 VGND.n10 VGND.n9 4.65
R176 VGND.n12 VGND.n11 4.65
R177 VGND.n14 VGND.n13 4.65
R178 VGND.n16 VGND.n15 4.65
R179 VGND.n18 VGND.n17 4.65
R180 VGND.n20 VGND.n19 4.65
R181 VGND.n23 VGND.n22 4.65
R182 VGND.n25 VGND.n24 4.65
R183 VGND.n27 VGND.n26 4.65
R184 VGND.n29 VGND.n28 4.65
R185 VGND.n32 VGND.n31 3.932
R186 VGND.n2 VGND.n1 3.897
R187 VGND.n4 VGND.n2 0.224
R188 VGND.n32 VGND.n29 0.137
R189 VGND VGND.n32 0.123
R190 VGND.n6 VGND.n4 0.119
R191 VGND.n8 VGND.n6 0.119
R192 VGND.n10 VGND.n8 0.119
R193 VGND.n12 VGND.n10 0.119
R194 VGND.n14 VGND.n12 0.119
R195 VGND.n16 VGND.n14 0.119
R196 VGND.n18 VGND.n16 0.119
R197 VGND.n20 VGND.n18 0.119
R198 VGND.n23 VGND.n20 0.119
R199 VGND.n25 VGND.n23 0.119
R200 VGND.n27 VGND.n25 0.119
R201 VGND.n29 VGND.n27 0.119
R202 A1.n0 A1.t0 266.138
R203 A1.n0 A1.t1 217.938
R204 A1 A1.n0 80.324
R205 a_1060_369.t0 a_1060_369.t1 226.095
R206 a_1281_47.t0 a_1281_47.t1 93.059
R207 A2.n0 A2.t1 372.865
R208 A2.n0 A2.t0 132.281
R209 A2 A2.n0 81.624
R210 a_193_47.n0 a_193_47.t0 66.666
R211 a_193_47.n0 a_193_47.t1 26.393
R212 a_193_47.n1 a_193_47.n0 14.4
R213 a_1064_47.n0 a_1064_47.t0 76.666
R214 a_1064_47.n0 a_1064_47.t1 27.339
R215 a_1064_47.n1 a_1064_47.n0 11.612
R216 a_397_47.t1 a_397_47.t0 93.516
R217 a_193_369.t1 a_193_369.t0 132.285
R218 A0.n0 A0.t1 299.374
R219 A0.n0 A0.t0 206.188
R220 A0 A0.n0 105.005
C0 A0 VGND 0.11fF
C1 VPWR X 0.28fF
C2 A3 S1 0.18fF
C3 S0 VGND 0.24fF
C4 VPB VPWR 0.18fF
C5 S0 A2 0.15fF
C6 S0 VPWR 0.10fF
C7 VGND X 0.20fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__mux4_4.ext - technology: sky130A

.subckt sky130_fd_sc_hd__mux4_4 VGND VPWR X S0 A2 A3 S1 A1 A0 VNB VPB
X0 X.t7 a_789_316.t4 VGND.t7 VNB.t13 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 X.t3 a_789_316.t5 VPWR.t7 VPB.t13 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 VPWR.t2 A0.t0 a_1280_413.t1 VPB.t6 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X3 a_873_316.t5 a_601_345.t2 a_789_316.t2 VNB.t5 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 a_601_345.t0 S1.t0 VPWR.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X5 VPWR.t1 S0.t0 a_27_47.t0 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X6 VGND.t6 a_789_316.t6 X.t6 VNB.t12 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 VGND.t5 a_789_316.t7 X.t5 VNB.t11 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 VPWR.t3 A3.t0 a_373_413.t0 VPB.t7 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X9 a_1282_47.t0 a_27_47.t2 a_873_316.t3 VNB.t8 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X10 a_1280_413.t0 S0.t1 a_873_316.t1 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11 a_1065_47.t1 A1.t0 VGND.t9 VNB.t15 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12 a_193_47.t0 A2.t0 VGND.t8 VNB.t14 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13 a_873_316.t2 S0.t2 a_1065_47.t0 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X14 X.t4 a_789_316.t8 VGND.t4 VNB.t10 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X15 a_1061_369.t0 A1.t1 VPWR.t9 VPB.t15 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X16 a_873_316.t4 a_27_47.t3 a_1061_369.t1 VPB.t8 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17 VPWR.t6 a_789_316.t9 X.t2 VPB.t12 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X18 X.t1 a_789_316.t10 VPWR.t5 VPB.t11 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X19 VGND.t3 A3.t1 a_398_47.t1 VNB.t7 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20 a_601_345.t1 S1.t1 VGND.t0 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21 a_873_316.t0 S1.t2 a_789_316.t0 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=540000u l=150000u
X22 a_193_369.t0 A2.t1 VPWR.t8 VPB.t14 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X23 a_789_316.t3 a_601_345.t3 a_288_47.t5 VPB.t5 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=540000u l=150000u
X24 a_398_47.t0 S0.t3 a_288_47.t1 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X25 VGND.t2 A0.t1 a_1282_47.t1 VNB.t6 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X26 a_373_413.t1 a_27_47.t4 a_288_47.t3 VPB.t9 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X27 a_288_47.t4 a_27_47.t5 a_193_47.t1 VNB.t9 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X28 VPWR.t4 a_789_316.t11 X.t0 VPB.t10 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X29 a_288_47.t0 S0.t4 a_193_369.t1 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X30 VGND.t1 S0.t5 a_27_47.t1 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X31 a_789_316.t1 S1.t3 a_288_47.t2 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
R0 a_789_316.n7 a_789_316.n6 292.5
R1 a_789_316.n6 a_789_316.n4 228.38
R2 a_789_316.n0 a_789_316.t9 212.079
R3 a_789_316.n1 a_789_316.t10 212.079
R4 a_789_316.n2 a_789_316.t11 212.079
R5 a_789_316.n3 a_789_316.t5 212.079
R6 a_789_316.n6 a_789_316.n5 174.352
R7 a_789_316.n0 a_789_316.t6 139.779
R8 a_789_316.n1 a_789_316.t4 139.779
R9 a_789_316.n2 a_789_316.t7 139.779
R10 a_789_316.n3 a_789_316.t8 139.779
R11 a_789_316.n2 a_789_316.n1 73.03
R12 a_789_316.n1 a_789_316.n0 61.345
R13 a_789_316.n4 a_789_316.n2 56.963
R14 a_789_316.t0 a_789_316.n7 49.25
R15 a_789_316.n7 a_789_316.t3 49.25
R16 a_789_316.n5 a_789_316.t1 40
R17 a_789_316.n5 a_789_316.t2 38.571
R18 a_789_316.n4 a_789_316.n3 4.381
R19 VGND.n16 VGND.t9 145.81
R20 VGND.n6 VGND.n5 119.1
R21 VGND.n2 VGND.t6 112.579
R22 VGND.n27 VGND.n26 107.239
R23 VGND.n36 VGND.n35 107.239
R24 VGND.n1 VGND.n0 69.685
R25 VGND.n5 VGND.t2 62.351
R26 VGND.n26 VGND.t0 57.142
R27 VGND.n26 VGND.t3 54.285
R28 VGND.n0 VGND.t5 39.692
R29 VGND.n35 VGND.t8 38.571
R30 VGND.n35 VGND.t1 38.571
R31 VGND.n5 VGND.t4 24.924
R32 VGND.n0 VGND.t7 24.923
R33 VGND.n4 VGND.n3 4.65
R34 VGND.n7 VGND.n6 4.65
R35 VGND.n9 VGND.n8 4.65
R36 VGND.n11 VGND.n10 4.65
R37 VGND.n13 VGND.n12 4.65
R38 VGND.n15 VGND.n14 4.65
R39 VGND.n17 VGND.n16 4.65
R40 VGND.n19 VGND.n18 4.65
R41 VGND.n21 VGND.n20 4.65
R42 VGND.n23 VGND.n22 4.65
R43 VGND.n25 VGND.n24 4.65
R44 VGND.n28 VGND.n27 4.65
R45 VGND.n30 VGND.n29 4.65
R46 VGND.n32 VGND.n31 4.65
R47 VGND.n34 VGND.n33 4.65
R48 VGND.n37 VGND.n36 3.932
R49 VGND.n2 VGND.n1 3.888
R50 VGND.n4 VGND.n2 0.225
R51 VGND.n37 VGND.n34 0.137
R52 VGND VGND.n37 0.121
R53 VGND.n7 VGND.n4 0.119
R54 VGND.n9 VGND.n7 0.119
R55 VGND.n11 VGND.n9 0.119
R56 VGND.n13 VGND.n11 0.119
R57 VGND.n15 VGND.n13 0.119
R58 VGND.n17 VGND.n15 0.119
R59 VGND.n19 VGND.n17 0.119
R60 VGND.n21 VGND.n19 0.119
R61 VGND.n23 VGND.n21 0.119
R62 VGND.n25 VGND.n23 0.119
R63 VGND.n28 VGND.n25 0.119
R64 VGND.n30 VGND.n28 0.119
R65 VGND.n32 VGND.n30 0.119
R66 VGND.n34 VGND.n32 0.119
R67 X.n0 X 298.998
R68 X.n7 X.n0 292.5
R69 X.n3 X.n1 180.079
R70 X.n3 X.n2 124.5
R71 X.n5 X.n4 92.5
R72 X.n6 X.n3 36
R73 X.n0 X.t2 26.595
R74 X.n0 X.t1 26.595
R75 X.n1 X.t0 26.595
R76 X.n1 X.t3 26.595
R77 X.n4 X.t6 24.923
R78 X.n4 X.t7 24.923
R79 X.n2 X.t5 24.923
R80 X.n2 X.t4 24.923
R81 X X.n6 10.24
R82 X.n7 X 8.467
R83 X X.n5 8.073
R84 X.n5 X 5.316
R85 X X.n7 4.923
R86 X.n6 X 3.15
R87 VNB VNB.t4 6438.23
R88 VNB.t0 VNB.t1 6147.06
R89 VNB.t5 VNB.t15 6082.35
R90 VNB.t2 VNB.t8 3558.82
R91 VNB.t9 VNB.t3 3558.82
R92 VNB.t7 VNB.t0 3494.12
R93 VNB.t15 VNB.t2 3461.76
R94 VNB.t3 VNB.t7 3105.88
R95 VNB.t8 VNB.t6 3073.53
R96 VNB.t14 VNB.t9 3073.53
R97 VNB.t1 VNB.t5 2750
R98 VNB.t4 VNB.t14 2717.65
R99 VNB.t11 VNB.t13 2417.58
R100 VNB.t6 VNB.t10 2400.4
R101 VNB.t13 VNB.t12 2030.77
R102 VNB.t10 VNB.t11 2030.77
R103 VPWR.n17 VPWR.t9 354.459
R104 VPWR.n28 VPWR.n27 320.326
R105 VPWR.n38 VPWR.n37 307.239
R106 VPWR.n6 VPWR.n5 174.594
R107 VPWR.n2 VPWR.t6 171.616
R108 VPWR.n1 VPWR.n0 126.121
R109 VPWR.n5 VPWR.t2 61.562
R110 VPWR.n0 VPWR.t4 42.355
R111 VPWR.n27 VPWR.t0 41.554
R112 VPWR.n27 VPWR.t3 41.554
R113 VPWR.n37 VPWR.t8 41.554
R114 VPWR.n37 VPWR.t1 41.554
R115 VPWR.n5 VPWR.t7 30.594
R116 VPWR.n0 VPWR.t5 26.595
R117 VPWR.n29 VPWR.n28 5.27
R118 VPWR.n4 VPWR.n3 4.65
R119 VPWR.n8 VPWR.n7 4.65
R120 VPWR.n10 VPWR.n9 4.65
R121 VPWR.n12 VPWR.n11 4.65
R122 VPWR.n14 VPWR.n13 4.65
R123 VPWR.n16 VPWR.n15 4.65
R124 VPWR.n18 VPWR.n17 4.65
R125 VPWR.n20 VPWR.n19 4.65
R126 VPWR.n22 VPWR.n21 4.65
R127 VPWR.n24 VPWR.n23 4.65
R128 VPWR.n26 VPWR.n25 4.65
R129 VPWR.n30 VPWR.n29 4.65
R130 VPWR.n32 VPWR.n31 4.65
R131 VPWR.n34 VPWR.n33 4.65
R132 VPWR.n36 VPWR.n35 4.65
R133 VPWR.n39 VPWR.n38 3.932
R134 VPWR.n2 VPWR.n1 3.888
R135 VPWR.n7 VPWR.n6 1.882
R136 VPWR.n4 VPWR.n2 0.225
R137 VPWR.n39 VPWR.n36 0.137
R138 VPWR VPWR.n39 0.121
R139 VPWR.n8 VPWR.n4 0.119
R140 VPWR.n10 VPWR.n8 0.119
R141 VPWR.n12 VPWR.n10 0.119
R142 VPWR.n14 VPWR.n12 0.119
R143 VPWR.n16 VPWR.n14 0.119
R144 VPWR.n18 VPWR.n16 0.119
R145 VPWR.n20 VPWR.n18 0.119
R146 VPWR.n22 VPWR.n20 0.119
R147 VPWR.n24 VPWR.n22 0.119
R148 VPWR.n26 VPWR.n24 0.119
R149 VPWR.n30 VPWR.n26 0.119
R150 VPWR.n32 VPWR.n30 0.119
R151 VPWR.n34 VPWR.n32 0.119
R152 VPWR.n36 VPWR.n34 0.119
R153 VPB.t1 VPB.t15 556.386
R154 VPB.t0 VPB.t5 556.386
R155 VPB.t9 VPB.t7 426.168
R156 VPB.t15 VPB.t8 399.532
R157 VPB.t3 VPB.t6 298.909
R158 VPB.t10 VPB.t11 295.95
R159 VPB.t6 VPB.t13 287.071
R160 VPB.t14 VPB.t4 284.112
R161 VPB.t11 VPB.t12 248.598
R162 VPB.t13 VPB.t10 248.598
R163 VPB.t8 VPB.t3 248.598
R164 VPB.t5 VPB.t1 248.598
R165 VPB.t7 VPB.t0 248.598
R166 VPB.t4 VPB.t9 248.598
R167 VPB.t2 VPB.t14 248.598
R168 VPB VPB.t2 189.408
R169 A0.n0 A0.t0 299.374
R170 A0.n0 A0.t1 206.188
R171 A0 A0.n0 105.005
R172 a_1280_413.n0 a_1280_413.t0 100.845
R173 a_1280_413.n1 a_1280_413.n0 77.392
R174 a_1280_413.n0 a_1280_413.t1 33.965
R175 a_601_345.t0 a_601_345.n1 466.234
R176 a_601_345.n0 a_601_345.t2 337.934
R177 a_601_345.n1 a_601_345.t1 201.267
R178 a_601_345.n1 a_601_345.n0 159.903
R179 a_601_345.n0 a_601_345.t3 157.453
R180 a_873_316.n2 a_873_316.n0 376.828
R181 a_873_316.t0 a_873_316.n3 347.139
R182 a_873_316.n2 a_873_316.n1 223.887
R183 a_873_316.n3 a_873_316.t5 220.887
R184 a_873_316.n1 a_873_316.t3 66.666
R185 a_873_316.n1 a_873_316.t2 66.666
R186 a_873_316.n0 a_873_316.t1 63.321
R187 a_873_316.n0 a_873_316.t4 63.321
R188 a_873_316.n3 a_873_316.n2 62.117
R189 S1.t0 S1.t2 769.592
R190 S1.n0 S1.t3 367.926
R191 S1.n1 S1.t0 350.711
R192 S1.n0 S1.t1 112.237
R193 S1.n2 S1.n1 76
R194 S1.n1 S1.n0 34.428
R195 S1.n2 S1 7.724
R196 S1 S1.n2 7.282
R197 S0.n1 S0.t3 445.045
R198 S0.n5 S0.t2 432.192
R199 S0.n7 S0.t0 287.994
R200 S0.n2 S0.t4 258.42
R201 S0.n5 S0.t1 254.388
R202 S0.n7 S0.t5 194.808
R203 S0.n6 S0.n5 90.486
R204 S0.n8 S0.n7 76
R205 S0 S0.n8 20.266
R206 S0.n4 S0.n3 18.793
R207 S0.n3 S0.n1 14.46
R208 S0 S0.n6 11.432
R209 S0.n3 S0.n2 6.159
R210 S0.n4 S0.n0 6.023
R211 S0.n6 S0.n4 4.518
R212 S0.n8 S0 3.911
R213 a_27_47.t0 a_27_47.n3 368.312
R214 a_27_47.n0 a_27_47.t5 245.944
R215 a_27_47.n3 a_27_47.t1 242.129
R216 a_27_47.n1 a_27_47.t2 241.28
R217 a_27_47.n0 a_27_47.t4 224.251
R218 a_27_47.n1 a_27_47.t3 146.443
R219 a_27_47.n3 a_27_47.n2 67.388
R220 a_27_47.n2 a_27_47.n1 11.44
R221 a_27_47.n2 a_27_47.n0 4.894
R222 A3.n0 A3.t0 313.804
R223 A3.n0 A3.t1 132.281
R224 A3.n1 A3.n0 76
R225 A3 A3.n1 8.52
R226 A3.n1 A3 5.632
R227 a_373_413.t0 a_373_413.t1 245.006
R228 a_373_413.n0 a_373_413.t0 101.896
R229 a_1282_47.t1 a_1282_47.t0 93.059
R230 A1.n0 A1.t1 282.237
R231 A1.n0 A1.t0 247.426
R232 A1 A1.n0 97.729
R233 a_1065_47.n0 a_1065_47.t0 76.666
R234 a_1065_47.n0 a_1065_47.t1 27.339
R235 a_1065_47.n1 a_1065_47.n0 11.612
R236 A2.n0 A2.t1 373.281
R237 A2.n0 A2.t0 132.281
R238 A2 A2.n0 81.624
R239 a_193_47.n0 a_193_47.t1 66.666
R240 a_193_47.n0 a_193_47.t0 26.393
R241 a_193_47.n1 a_193_47.n0 14.4
R242 a_1061_369.t0 a_1061_369.t1 226.095
R243 a_398_47.t1 a_398_47.t0 93.516
R244 a_193_369.t0 a_193_369.t1 134.63
R245 a_288_47.t5 a_288_47.n3 341.75
R246 a_288_47.n2 a_288_47.n1 329.77
R247 a_288_47.n2 a_288_47.n0 244.968
R248 a_288_47.n3 a_288_47.t2 233.964
R249 a_288_47.n0 a_288_47.t1 66.666
R250 a_288_47.n0 a_288_47.t4 66.666
R251 a_288_47.n1 a_288_47.t3 63.321
R252 a_288_47.n1 a_288_47.t0 63.321
R253 a_288_47.n3 a_288_47.n2 31.496
C0 VGND VPWR 0.11fF
C1 VGND X 0.49fF
C2 A3 S1 0.18fF
C3 X VPWR 0.67fF
C4 S0 A2 0.15fF
C5 VPB VPWR 0.19fF
C6 VGND S0 0.24fF
C7 A0 VGND 0.11fF
C8 S0 VPWR 0.10fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__nand2_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__nand2_1 Y B A VGND VPWR VNB VPB
X0 VPWR.t0 A.t0 Y.t1 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 Y.t0 A.t1 a_113_47.t1 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 a_113_47.t0 B.t0 VGND.t0 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 Y.t2 B.t1 VPWR.t1 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
R0 A.n0 A.t0 230.154
R1 A.n0 A.t1 157.854
R2 A A.n0 78.101
R3 Y Y.n0 139.93
R4 Y.n1 Y.t0 94.258
R5 Y.n0 Y.t1 26.595
R6 Y.n0 Y.t2 26.595
R7 Y.n1 Y 16.564
R8 Y Y.n1 9.035
R9 Y.n1 Y 1.726
R10 VPWR.n0 VPWR.t0 155.759
R11 VPWR.n0 VPWR.t1 153.591
R12 VPWR VPWR.n0 0.128
R13 VPB.t1 VPB.t0 248.598
R14 VPB VPB.t1 207.165
R15 a_113_47.t0 a_113_47.t1 49.846
R16 VNB VNB.t0 6198.96
R17 VNB.t0 VNB.t1 2030.77
R18 B.n0 B.t1 229.368
R19 B.n0 B.t0 157.068
R20 B B.n0 81.925
R21 VGND VGND.t0 108.644
C0 Y VGND 0.21fF
C1 A Y 0.11fF
C2 VPWR Y 0.38fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__nand2_2.ext - technology: sky130A

.subckt sky130_fd_sc_hd__nand2_2 Y A B VGND VPWR VNB VPB
X0 VPWR.t3 A.t0 Y.t4 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 Y.t3 A.t1 VPWR.t2 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 VPWR.t0 B.t0 Y.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 a_27_47.t3 B.t1 VGND.t1 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 a_27_47.t1 A.t2 Y.t5 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 Y.t2 A.t3 a_27_47.t0 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 Y.t1 B.t2 VPWR.t1 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 VGND.t0 B.t3 a_27_47.t2 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
R0 A.n0 A.t0 212.079
R1 A.n1 A.t1 212.079
R2 A.n0 A.t2 139.779
R3 A.n1 A.t3 139.779
R4 A.n3 A.n2 76
R5 A.n2 A.n0 30.672
R6 A.n2 A.n1 30.672
R7  A.n3 23.04
R8 A.n3 A 0.512
R9 Y.n3 Y.n1 146.035
R10 Y.n4 Y.n0 113.748
R11 Y.n3 Y.n2 107.635
R12 Y.n1 Y.t0 26.595
R13 Y.n1 Y.t1 26.595
R14 Y.n2 Y.t4 26.595
R15 Y.n2 Y.t3 26.595
R16 Y Y.n3 24.994
R17 Y.n0 Y.t5 24.923
R18 Y.n0 Y.t2 24.923
R19 Y.n4 Y 14.857
R20 Y Y.n4 0.685
R21 VPWR.n2 VPWR.t3 200.022
R22 VPWR.n1 VPWR.n0 174.594
R23 VPWR.n5 VPWR.t1 151.631
R24 VPWR.n0 VPWR.t2 26.595
R25 VPWR.n0 VPWR.t0 26.595
R26 VPWR.n2 VPWR.n1 7.817
R27 VPWR.n4 VPWR.n3 4.65
R28 VPWR.n6 VPWR.n5 4.65
R29 VPWR.n4 VPWR.n2 0.218
R30 VPWR.n6 VPWR.n4 0.119
R31 VPWR VPWR.n6 0.02
R32 VPB.t2 VPB.t3 248.598
R33 VPB.t0 VPB.t2 248.598
R34 VPB.t1 VPB.t0 248.598
R35 VPB VPB.t1 189.408
R36 B.n0 B.t0 212.079
R37 B.n1 B.t2 212.079
R38 B.n0 B.t1 139.779
R39 B.n1 B.t3 139.779
R40 B B.n2 79.584
R41 B.n2 B.n0 30.672
R42 B.n2 B.n1 30.672
R43  B 23.552
R44 VGND VGND.n0 119.177
R45 VGND.n0 VGND.t1 24.923
R46 VGND.n0 VGND.t0 24.923
R47 a_27_47.t1 a_27_47.n1 229.699
R48 a_27_47.n1 a_27_47.t2 141.802
R49 a_27_47.n1 a_27_47.n0 42.273
R50 a_27_47.n0 a_27_47.t0 24.923
R51 a_27_47.n0 a_27_47.t3 24.923
R52 VNB VNB.t2 6053.91
R53 VNB.t0 VNB.t1 2030.77
R54 VNB.t3 VNB.t0 2030.77
R55 VNB.t2 VNB.t3 2030.77
C0 VPWR Y 0.72fF
C1 A Y 0.32fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__nand2_4.ext - technology: sky130A

.subckt sky130_fd_sc_hd__nand2_4 Y A B VGND VPWR VNB VPB
X0 a_27_47.t7 A.t0 Y.t7 VNB.t7 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 a_27_47.t6 A.t1 Y.t6 VNB.t6 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 Y.t11 A.t2 VPWR.t7 VPB.t7 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 VPWR.t1 B.t0 Y.t1 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 Y.t2 B.t1 VPWR.t2 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 VPWR.t3 B.t2 Y.t3 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 a_27_47.t2 B.t3 VGND.t3 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 a_27_47.t3 B.t4 VGND.t2 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 VPWR.t6 A.t3 Y.t10 VPB.t6 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 VGND.t1 B.t5 a_27_47.t0 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 Y.t5 A.t4 a_27_47.t5 VNB.t5 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 Y.t9 A.t5 VPWR.t5 VPB.t5 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 Y.t4 A.t6 a_27_47.t4 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 VPWR.t4 A.t7 Y.t8 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14 Y.t0 B.t6 VPWR.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 VGND.t0 B.t7 a_27_47.t1 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
R0 A.n0 A.t3 212.079
R1 A.n3 A.t5 212.079
R2 A.n5 A.t7 212.079
R3 A.n4 A.t2 212.079
R4 A.n0 A.t1 139.779
R5 A.n3 A.t6 139.779
R6 A.n5 A.t0 139.779
R7 A.n4 A.t4 139.779
R8 A A.n6 82.656
R9 A.n2 A.n1 76
R10 A.n5 A.n4 61.345
R11 A.n1 A.n0 30.672
R12 A.n6 A.n3 30.672
R13 A.n6 A.n5 30.672
R14 A  23.552
R15 A A.n2 14.848
R16 A.n2 A 8.704
R17 Y.n2 Y.n0 158.458
R18 Y.n9 Y.n7 149.347
R19 Y.n5 Y.n3 146.035
R20 Y.n5 Y.n4 107.635
R21 Y.n2 Y.n1 104.452
R22 Y.n9 Y.n8 92.5
R23 Y.n1 Y.t8 26.595
R24 Y.n1 Y.t11 26.595
R25 Y.n3 Y.t3 26.595
R26 Y.n3 Y.t0 26.595
R27 Y.n4 Y.t1 26.595
R28 Y.n4 Y.t2 26.595
R29 Y.n0 Y.t10 26.595
R30 Y.n0 Y.t9 26.595
R31 Y.n7 Y.t6 24.923
R32 Y.n7 Y.t4 24.923
R33 Y.n8 Y.t7 24.923
R34 Y.n8 Y.t5 24.923
R35 Y Y.n5 22.964
R36 Y Y.n9 18.893
R37 Y.n6 Y.n2 13.929
R38 Y.n6 Y 13.929
R39 Y Y.n6 1.196
R40 a_27_47.t6 a_27_47.n5 136.83
R41 a_27_47.n2 a_27_47.t1 126.176
R42 a_27_47.n5 a_27_47.n0 92.5
R43 a_27_47.n5 a_27_47.n4 54.999
R44 a_27_47.n2 a_27_47.n1 52.818
R45 a_27_47.n4 a_27_47.n2 46.921
R46 a_27_47.n4 a_27_47.n3 42.273
R47 a_27_47.n0 a_27_47.t4 24.923
R48 a_27_47.n0 a_27_47.t7 24.923
R49 a_27_47.n3 a_27_47.t5 24.923
R50 a_27_47.n3 a_27_47.t3 24.923
R51 a_27_47.n1 a_27_47.t0 24.923
R52 a_27_47.n1 a_27_47.t2 24.923
R53 VNB VNB.t1 6053.91
R54 VNB.t4 VNB.t6 2030.77
R55 VNB.t7 VNB.t4 2030.77
R56 VNB.t5 VNB.t7 2030.77
R57 VNB.t3 VNB.t5 2030.77
R58 VNB.t0 VNB.t3 2030.77
R59 VNB.t2 VNB.t0 2030.77
R60 VNB.t1 VNB.t2 2030.77
R61 VPWR.n2 VPWR.t6 202.393
R62 VPWR.n12 VPWR.n11 174.594
R63 VPWR.n6 VPWR.n5 174.594
R64 VPWR.n1 VPWR.n0 174.594
R65 VPWR.n17 VPWR.t0 152.162
R66 VPWR.n11 VPWR.t2 26.595
R67 VPWR.n11 VPWR.t3 26.595
R68 VPWR.n5 VPWR.t7 26.595
R69 VPWR.n5 VPWR.t1 26.595
R70 VPWR.n0 VPWR.t5 26.595
R71 VPWR.n0 VPWR.t4 26.595
R72 VPWR.n2 VPWR.n1 19.667
R73 VPWR.n7 VPWR.n6 9.788
R74 VPWR.n4 VPWR.n3 4.65
R75 VPWR.n8 VPWR.n7 4.65
R76 VPWR.n10 VPWR.n9 4.65
R77 VPWR.n14 VPWR.n13 4.65
R78 VPWR.n16 VPWR.n15 4.65
R79 VPWR.n18 VPWR.n17 4.65
R80 VPWR.n13 VPWR.n12 3.764
R81 VPWR.n4 VPWR.n2 0.414
R82 VPWR.n8 VPWR.n4 0.119
R83 VPWR.n10 VPWR.n8 0.119
R84 VPWR.n14 VPWR.n10 0.119
R85 VPWR.n16 VPWR.n14 0.119
R86 VPWR.n18 VPWR.n16 0.119
R87 VPWR VPWR.n18 0.02
R88 VPB.t5 VPB.t6 248.598
R89 VPB.t4 VPB.t5 248.598
R90 VPB.t7 VPB.t4 248.598
R91 VPB.t1 VPB.t7 248.598
R92 VPB.t2 VPB.t1 248.598
R93 VPB.t3 VPB.t2 248.598
R94 VPB.t0 VPB.t3 248.598
R95 VPB VPB.t0 189.408
R96 B.n0 B.t0 212.079
R97 B.n2 B.t1 212.079
R98 B.n6 B.t2 212.079
R99 B.n7 B.t6 212.079
R100 B.n0 B.t4 139.779
R101 B.n2 B.t5 139.779
R102 B.n6 B.t3 139.779
R103 B.n7 B.t7 139.779
R104 B.n5 B.n4 76
R105 B.n9 B.n8 76
R106 B.n1 B.n0 30.672
R107 B.n2 B.n1 30.672
R108 B.n5 B.n2 30.672
R109 B.n6 B.n5 30.672
R110 B.n8 B.n6 30.672
R111 B.n8 B.n7 30.672
R112 B.n4 B.n3 21.504
R113 B.n9 B 19.968
R114 B B.n10 17.152
R115 B.n10 B 6.4
R116 B B.n9 3.584
R117 B.n4 B 1.536
R118 B.n3 B 0.512
R119 VGND.n2 VGND.n0 122.93
R120 VGND.n2 VGND.n1 118.929
R121 VGND.n0 VGND.t2 24.923
R122 VGND.n0 VGND.t1 24.923
R123 VGND.n1 VGND.t3 24.923
R124 VGND.n1 VGND.t0 24.923
R125 VGND VGND.n2 0.249
C0 Y B 0.26fF
C1 VPWR Y 1.29fF
C2 Y A 0.29fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__nand2_8.ext - technology: sky130A

.subckt sky130_fd_sc_hd__nand2_8 A B Y VGND VPWR VNB VPB
X0 a_27_47.t15 B.t0 VGND.t7 VNB.t15 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 Y.t15 A.t0 VPWR.t15 VPB.t15 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 a_27_47.t14 B.t1 VGND.t6 VNB.t14 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 a_27_47.t5 A.t1 Y.t23 VNB.t5 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 a_27_47.t6 A.t2 Y.t22 VNB.t6 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 Y.t7 B.t2 VPWR.t7 VPB.t7 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 VPWR.t6 B.t3 Y.t6 VPB.t6 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 Y.t21 A.t3 a_27_47.t7 VNB.t7 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 Y.t20 A.t4 a_27_47.t2 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 Y.t19 A.t5 a_27_47.t3 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 Y.t5 B.t4 VPWR.t5 VPB.t5 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 VPWR.t14 A.t6 Y.t14 VPB.t14 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 Y.t13 A.t7 VPWR.t13 VPB.t13 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13 VPWR.t4 B.t5 Y.t4 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14 VPWR.t12 A.t8 Y.t12 VPB.t12 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 a_27_47.t13 B.t6 VGND.t5 VNB.t13 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X16 a_27_47.t12 B.t7 VGND.t4 VNB.t12 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X17 a_27_47.t4 A.t9 Y.t18 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X18 Y.t11 A.t10 VPWR.t11 VPB.t11 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X19 VPWR.t3 B.t8 Y.t3 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X20 VGND.t3 B.t9 a_27_47.t11 VNB.t11 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X21 VGND.t2 B.t10 a_27_47.t10 VNB.t10 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X22 Y.t2 B.t11 VPWR.t2 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X23 VPWR.t10 A.t11 Y.t10 VPB.t10 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X24 VGND.t1 B.t12 a_27_47.t9 VNB.t9 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X25 Y.t17 A.t12 a_27_47.t0 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X26 VPWR.t1 B.t13 Y.t1 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X27 Y.t9 A.t13 VPWR.t9 VPB.t9 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X28 Y.t0 B.t14 VPWR.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X29 VPWR.t8 A.t14 Y.t8 VPB.t8 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X30 VGND.t0 B.t15 a_27_47.t8 VNB.t8 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X31 a_27_47.t1 A.t15 Y.t16 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
R0 B.n1 B.t8 221.719
R1 B.n3 B.t11 221.719
R2 B.n0 B.t13 221.719
R3 B.n8 B.t2 221.719
R4 B.n17 B.t3 221.719
R5 B.n18 B.t4 221.719
R6 B.n14 B.t5 221.719
R7 B.n11 B.t14 221.719
R8 B.n1 B.t1 149.419
R9 B.n3 B.t12 149.419
R10 B.n0 B.t0 149.419
R11 B.n8 B.t10 149.419
R12 B.n17 B.t7 149.419
R13 B.n18 B.t9 149.419
R14 B.n14 B.t6 149.419
R15 B.n11 B.t15 149.419
R16 B.n2 B 92.872
R17 B.n5 B.n4 76
R18 B.n7 B.n6 76
R19 B.n10 B.n9 76
R20 B.n20 B.n19 76
R21 B.n16 B.n15 76
R22 B.n13 B.n12 76
R23 B.n14 B.n13 38.381
R24 B.n2 B.n1 37.488
R25 B.n3 B.n2 37.488
R26 B.n4 B.n3 37.488
R27 B.n4 B.n0 37.488
R28 B.n7 B.n0 37.488
R29 B.n8 B.n7 37.488
R30 B.n9 B.n8 37.488
R31 B.n19 B.n17 37.488
R32 B.n19 B.n18 37.488
R33 B.n15 B.n14 37.488
R34 B.n13 B.n11 36.596
R35 B.n20 B.n16 24.436
R36 B B.n10 23.854
R37 B.n12 B 22.981
R38 B.n6 B 21.527
R39 B B.n5 19.2
R40 B.n5 B 7.563
R41 B.n6 B 5.236
R42 B.n12 B 3.781
R43 B.n10 B 2.909
R44 B.n16 B 1.745
R45 B B.n20 0.581
R46 VGND.n3 VGND.n0 126.758
R47 VGND.n2 VGND.n1 116.217
R48 VGND.n7 VGND.n6 116.217
R49 VGND.n13 VGND.n12 116.217
R50 VGND.n0 VGND.t6 24.923
R51 VGND.n0 VGND.t1 24.923
R52 VGND.n1 VGND.t7 24.923
R53 VGND.n1 VGND.t2 24.923
R54 VGND.n6 VGND.t4 24.923
R55 VGND.n6 VGND.t3 24.923
R56 VGND.n12 VGND.t5 24.923
R57 VGND.n12 VGND.t0 24.923
R58 VGND.n3 VGND.n2 16.678
R59 VGND.n8 VGND.n7 6.776
R60 VGND.n5 VGND.n4 4.65
R61 VGND.n9 VGND.n8 4.65
R62 VGND.n11 VGND.n10 4.65
R63 VGND.n15 VGND.n14 4.65
R64 VGND.n14 VGND.n13 0.752
R65 VGND.n5 VGND.n3 0.395
R66 VGND.n9 VGND.n5 0.119
R67 VGND.n11 VGND.n9 0.119
R68 VGND.n15 VGND.n11 0.119
R69 VGND.n16 VGND.n15 0.119
R70 VGND VGND.n16 0.02
R71 a_27_47.n7 a_27_47.t4 135.406
R72 a_27_47.n1 a_27_47.t8 130.175
R73 a_27_47.n7 a_27_47.n6 92.5
R74 a_27_47.n9 a_27_47.n8 92.5
R75 a_27_47.n11 a_27_47.n10 92.5
R76 a_27_47.n1 a_27_47.n0 52.431
R77 a_27_47.n3 a_27_47.n2 52.431
R78 a_27_47.n5 a_27_47.n4 52.431
R79 a_27_47.n12 a_27_47.n11 51.51
R80 a_27_47.n12 a_27_47.n5 50.452
R81 a_27_47.n9 a_27_47.n7 46.747
R82 a_27_47.n11 a_27_47.n9 46.747
R83 a_27_47.n13 a_27_47.n12 42.273
R84 a_27_47.n3 a_27_47.n1 38.4
R85 a_27_47.n5 a_27_47.n3 38.4
R86 a_27_47.n0 a_27_47.t11 24.923
R87 a_27_47.n0 a_27_47.t13 24.923
R88 a_27_47.n2 a_27_47.t10 24.923
R89 a_27_47.n2 a_27_47.t12 24.923
R90 a_27_47.n4 a_27_47.t9 24.923
R91 a_27_47.n4 a_27_47.t15 24.923
R92 a_27_47.n10 a_27_47.t3 24.923
R93 a_27_47.n10 a_27_47.t6 24.923
R94 a_27_47.n8 a_27_47.t7 24.923
R95 a_27_47.n8 a_27_47.t1 24.923
R96 a_27_47.n6 a_27_47.t2 24.923
R97 a_27_47.n6 a_27_47.t5 24.923
R98 a_27_47.n13 a_27_47.t0 24.923
R99 a_27_47.t14 a_27_47.n13 24.923
R100 VNB VNB.t8 6053.91
R101 VNB.t2 VNB.t4 2030.77
R102 VNB.t5 VNB.t2 2030.77
R103 VNB.t7 VNB.t5 2030.77
R104 VNB.t1 VNB.t7 2030.77
R105 VNB.t3 VNB.t1 2030.77
R106 VNB.t6 VNB.t3 2030.77
R107 VNB.t0 VNB.t6 2030.77
R108 VNB.t14 VNB.t0 2030.77
R109 VNB.t9 VNB.t14 2030.77
R110 VNB.t15 VNB.t9 2030.77
R111 VNB.t10 VNB.t15 2030.77
R112 VNB.t12 VNB.t10 2030.77
R113 VNB.t11 VNB.t12 2030.77
R114 VNB.t13 VNB.t11 2030.77
R115 VNB.t8 VNB.t13 2030.77
R116 A.n0 A.t11 221.719
R117 A.n1 A.t13 221.719
R118 A.n3 A.t14 221.719
R119 A.n4 A.t0 221.719
R120 A.n14 A.t6 221.719
R121 A.n7 A.t7 221.719
R122 A.n9 A.t8 221.719
R123 A.n8 A.t10 221.719
R124 A.n0 A.t9 149.419
R125 A.n1 A.t4 149.419
R126 A.n3 A.t1 149.419
R127 A.n4 A.t3 149.419
R128 A.n14 A.t15 149.419
R129 A.n7 A.t5 149.419
R130 A.n9 A.t2 149.419
R131 A.n8 A.t12 149.419
R132 A.n2 A 76.64
R133 A.n6 A.n5 76
R134 A.n16 A.n15 76
R135 A.n13 A.n12 76
R136 A.n11 A.n10 76
R137 A.n1 A.n0 74.977
R138 A.n9 A.n8 74.977
R139 A.n2 A.n1 37.488
R140 A.n3 A.n2 37.488
R141 A.n5 A.n3 37.488
R142 A.n5 A.n4 37.488
R143 A.n15 A.n14 37.488
R144 A.n14 A.n13 37.488
R145 A.n13 A.n7 37.488
R146 A.n10 A.n7 37.488
R147 A.n10 A.n9 37.488
R148 A.n6 A 26.24
R149 A A.n16 23.68
R150 A.n12 A 21.12
R151 A A.n11 18.56
R152 A.n11 A 10.88
R153 A.n12 A 8.32
R154 A.n16 A 5.76
R155 A A.n6 3.2
R156 VPWR.n34 VPWR.n33 174.594
R157 VPWR.n28 VPWR.n27 174.594
R158 VPWR.n22 VPWR.n21 174.594
R159 VPWR.n18 VPWR.n17 174.594
R160 VPWR.n12 VPWR.n11 174.594
R161 VPWR.n6 VPWR.n5 174.594
R162 VPWR.n1 VPWR.n0 174.594
R163 VPWR.n2 VPWR.t10 168.009
R164 VPWR.n39 VPWR.t0 152.162
R165 VPWR.n33 VPWR.t5 26.595
R166 VPWR.n33 VPWR.t4 26.595
R167 VPWR.n27 VPWR.t7 26.595
R168 VPWR.n27 VPWR.t6 26.595
R169 VPWR.n21 VPWR.t2 26.595
R170 VPWR.n21 VPWR.t1 26.595
R171 VPWR.n17 VPWR.t11 26.595
R172 VPWR.n17 VPWR.t3 26.595
R173 VPWR.n11 VPWR.t13 26.595
R174 VPWR.n11 VPWR.t12 26.595
R175 VPWR.n5 VPWR.t15 26.595
R176 VPWR.n5 VPWR.t14 26.595
R177 VPWR.n0 VPWR.t9 26.595
R178 VPWR.n0 VPWR.t8 26.595
R179 VPWR.n23 VPWR.n22 15.811
R180 VPWR.n19 VPWR.n18 12.8
R181 VPWR.n29 VPWR.n28 9.788
R182 VPWR.n2 VPWR.n1 9.323
R183 VPWR.n13 VPWR.n12 6.776
R184 VPWR.n4 VPWR.n3 4.65
R185 VPWR.n8 VPWR.n7 4.65
R186 VPWR.n10 VPWR.n9 4.65
R187 VPWR.n14 VPWR.n13 4.65
R188 VPWR.n16 VPWR.n15 4.65
R189 VPWR.n20 VPWR.n19 4.65
R190 VPWR.n24 VPWR.n23 4.65
R191 VPWR.n26 VPWR.n25 4.65
R192 VPWR.n30 VPWR.n29 4.65
R193 VPWR.n32 VPWR.n31 4.65
R194 VPWR.n36 VPWR.n35 4.65
R195 VPWR.n38 VPWR.n37 4.65
R196 VPWR.n40 VPWR.n39 4.65
R197 VPWR.n35 VPWR.n34 3.764
R198 VPWR.n7 VPWR.n6 0.752
R199 VPWR.n4 VPWR.n2 0.218
R200 VPWR.n8 VPWR.n4 0.119
R201 VPWR.n10 VPWR.n8 0.119
R202 VPWR.n14 VPWR.n10 0.119
R203 VPWR.n16 VPWR.n14 0.119
R204 VPWR.n20 VPWR.n16 0.119
R205 VPWR.n24 VPWR.n20 0.119
R206 VPWR.n26 VPWR.n24 0.119
R207 VPWR.n30 VPWR.n26 0.119
R208 VPWR.n32 VPWR.n30 0.119
R209 VPWR.n36 VPWR.n32 0.119
R210 VPWR.n38 VPWR.n36 0.119
R211 VPWR.n40 VPWR.n38 0.119
R212 VPWR VPWR.n40 0.02
R213 Y.n2 Y.n0 140.856
R214 Y.n2 Y.n1 108.216
R215 Y.n4 Y.n3 108.216
R216 Y.n6 Y.n5 108.216
R217 Y.n11 Y.n10 108.216
R218 Y.n13 Y.n12 108.216
R219 Y.n15 Y.n14 108.216
R220 Y.n9 Y.n8 104.452
R221 Y.n23 Y.n22 92.5
R222 Y.n21 Y.n20 92.5
R223 Y.n19 Y.n18 92.5
R224 Y.n17 Y.n16 92.5
R225 Y.n11 Y.n9 43.2
R226 Y.n19 Y.n17 43.008
R227 Y.n21 Y.n19 43.008
R228 Y.n23 Y.n21 43.008
R229 Y.n17 Y.n15 34.598
R230 Y.n4 Y.n2 32.64
R231 Y.n6 Y.n4 32.64
R232 Y.n13 Y.n11 32.64
R233 Y.n15 Y.n13 32.64
R234 Y Y.n6 29.76
R235 Y.n14 Y.t10 26.595
R236 Y.n14 Y.t9 26.595
R237 Y.n8 Y.t12 26.595
R238 Y.n8 Y.t11 26.595
R239 Y.n0 Y.t4 26.595
R240 Y.n0 Y.t0 26.595
R241 Y.n1 Y.t6 26.595
R242 Y.n1 Y.t5 26.595
R243 Y.n3 Y.t1 26.595
R244 Y.n3 Y.t7 26.595
R245 Y.n5 Y.t3 26.595
R246 Y.n5 Y.t2 26.595
R247 Y.n10 Y.t14 26.595
R248 Y.n10 Y.t13 26.595
R249 Y.n12 Y.t8 26.595
R250 Y.n12 Y.t15 26.595
R251 Y.n16 Y.t18 24.923
R252 Y.n16 Y.t20 24.923
R253 Y.n18 Y.t23 24.923
R254 Y.n18 Y.t21 24.923
R255 Y.n20 Y.t16 24.923
R256 Y.n20 Y.t19 24.923
R257 Y.n22 Y.t22 24.923
R258 Y.n22 Y.t17 24.923
R259 Y Y.n23 11.985
R260 Y.n9 Y.n7 10.24
R261 Y.n7 Y 3.2
R262 Y Y.n7 0.533
R263 VPB.t9 VPB.t10 248.598
R264 VPB.t8 VPB.t9 248.598
R265 VPB.t15 VPB.t8 248.598
R266 VPB.t14 VPB.t15 248.598
R267 VPB.t13 VPB.t14 248.598
R268 VPB.t12 VPB.t13 248.598
R269 VPB.t11 VPB.t12 248.598
R270 VPB.t3 VPB.t11 248.598
R271 VPB.t2 VPB.t3 248.598
R272 VPB.t1 VPB.t2 248.598
R273 VPB.t7 VPB.t1 248.598
R274 VPB.t6 VPB.t7 248.598
R275 VPB.t5 VPB.t6 248.598
R276 VPB.t4 VPB.t5 248.598
R277 VPB.t0 VPB.t4 248.598
R278 VPB VPB.t0 189.408
C0 VPWR Y 2.62fF
C1 VPB B 0.11fF
C2 VPWR VGND 0.16fF
C3 B Y 0.56fF
C4 VPB A 0.10fF
C5 A Y 0.96fF
C6 VPB VPWR 0.15fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__nand2b_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__nand2b_1 Y A_N B VGND VPWR VNB VPB
X0 VGND.t0 A_N.t0 a_27_93.t0 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1 Y.t1 a_27_93.t2 a_206_47.t0 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 a_206_47.t1 B.t0 VGND.t1 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 VPWR.t2 a_27_93.t3 Y.t0 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 Y.t2 B.t1 VPWR.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 VPWR.t1 A_N.t1 a_27_93.t1 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
R0 A_N.n0 A_N.t1 137.175
R1 A_N.n0 A_N.t0 121.108
R2 A_N A_N.n0 82.666
R3 a_27_93.n1 a_27_93.t1 451.554
R4 a_27_93.n0 a_27_93.t3 236.179
R5 a_27_93.t0 a_27_93.n1 226.722
R6 a_27_93.n0 a_27_93.t2 163.879
R7 a_27_93.n1 a_27_93.n0 76
R8 VGND VGND.n0 113.387
R9 VGND.n0 VGND.t0 58.571
R10 VGND.n0 VGND.t1 24
R11 VNB VNB.t0 6053.91
R12 VNB.t0 VNB.t2 2345.05
R13 VNB.t2 VNB.t1 2030.77
R14 a_206_47.t0 a_206_47.t1 49.846
R15 Y Y.n0 192.636
R16 Y Y.t1 185.929
R17 Y.n0 Y.t0 26.595
R18 Y.n0 Y.t2 26.595
R19 B.n0 B.t1 236.179
R20 B.n0 B.t0 163.879
R21 B B.n0 92.533
R22 VPWR.n1 VPWR.t2 582.742
R23 VPWR.n1 VPWR.n0 175.074
R24 VPWR.n0 VPWR.t1 96.154
R25 VPWR.n0 VPWR.t0 25.61
R26 VPWR VPWR.n1 0.21
R27 VPB.t1 VPB.t0 287.071
R28 VPB.t0 VPB.t2 248.598
R29 VPB VPB.t1 189.408
C0 Y VGND 0.15fF
C1 VPWR Y 0.30fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__nand2b_2.ext - technology: sky130A

.subckt sky130_fd_sc_hd__nand2b_2 B Y A_N VGND VPWR VNB VPB
X0 Y.t5 B.t0 VPWR.t4 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 VGND.t2 A_N.t0 a_27_93.t1 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 VGND.t0 B.t1 a_229_47.t3 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 Y.t0 a_27_93.t2 a_229_47.t1 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 a_229_47.t0 a_27_93.t3 Y.t1 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 Y.t2 a_27_93.t4 VPWR.t1 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 VPWR.t2 a_27_93.t5 Y.t3 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 VPWR.t3 B.t2 Y.t4 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 a_229_47.t2 B.t3 VGND.t1 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 VPWR.t0 A_N.t1 a_27_93.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
R0 B.n0 B.t3 869.206
R1 B.n2 B.t0 232.43
R2 B.n1 B.t2 218.506
R3 B.n2 B.t1 149.419
R4 B.n0 B 88.888
R5 B.n4 B.n3 76
R6 B.n3 B.n1 37.01
R7 B.n1 B.n0 36.15
R8 B.n4 B 28.16
R9 B.n3 B.n2 26.777
R10 B B.n5 23.36
R11 B.n5  11.452
R12 B.n5  6.08
R13 B B.n4 1.28
R14 VPWR.n4 VPWR.n3 292.5
R15 VPWR.n1 VPWR.n0 292.5
R16 VPWR.n10 VPWR.n9 171.169
R17 VPWR.n2 VPWR.t3 149.888
R18 VPWR.n9 VPWR.t0 98.5
R19 VPWR.n0 VPWR.t4 38.415
R20 VPWR.n3 VPWR.t2 26.595
R21 VPWR.n9 VPWR.t1 25.61
R22 VPWR.n2 VPWR.n1 5.653
R23 VPWR.n6 VPWR.n5 4.65
R24 VPWR.n8 VPWR.n7 4.65
R25 VPWR.n11 VPWR.n10 4.031
R26 VPWR.n5 VPWR.n4 0.812
R27 VPWR.n6 VPWR.n2 0.217
R28 VPWR.n11 VPWR.n8 0.135
R29 VPWR VPWR.n11 0.124
R30 VPWR.n8 VPWR.n6 0.119
R31 Y.n2 Y.n0 165.001
R32 Y.n2 Y.n1 136.75
R33 Y Y.n3 94.557
R34 Y.n0 Y.t3 32.505
R35 Y.n0 Y.t2 32.505
R36 Y.n1 Y.t4 26.595
R37 Y.n1 Y.t5 26.595
R38 Y.n3 Y.t1 24.923
R39 Y.n3 Y.t0 24.923
R40 Y Y.n2 6.171
R41 VPB.t2 VPB.t4 485.358
R42 VPB.t0 VPB.t1 290.031
R43 VPB.t1 VPB.t2 284.112
R44 VPB.t4 VPB.t3 248.598
R45 VPB VPB.t0 189.408
R46 A_N.n0 A_N.t1 147.296
R47 A_N.n0 A_N.t0 131.229
R48 A_N A_N.n0 78.715
R49 a_27_93.t0 a_27_93.n3 355.821
R50 a_27_93.n2 a_27_93.t4 263.67
R51 a_27_93.n0 a_27_93.t3 224.396
R52 a_27_93.n1 a_27_93.t5 221.719
R53 a_27_93.n3 a_27_93.t1 191.654
R54 a_27_93.n0 a_27_93.t2 149.419
R55 a_27_93.n3 a_27_93.n2 144.232
R56 a_27_93.n2 a_27_93.n1 43.737
R57 a_27_93.n1 a_27_93.n0 7.14
R58 VGND.n1 VGND.t2 119.048
R59 VGND.n1 VGND.n0 117.414
R60 VGND.n0 VGND.t1 24.923
R61 VGND.n0 VGND.t0 24.923
R62 VGND VGND.n1 0.141
R63 VNB VNB.t4 6053.91
R64 VNB.t4 VNB.t1 4883.52
R65 VNB.t3 VNB.t2 2030.77
R66 VNB.t0 VNB.t3 2030.77
R67 VNB.t1 VNB.t0 2030.77
R68 a_229_47.t1 a_229_47.n1 140.155
R69 a_229_47.n1 a_229_47.t2 134.321
R70 a_229_47.n1 a_229_47.n0 42.273
R71 a_229_47.n0 a_229_47.t3 24.923
R72 a_229_47.n0 a_229_47.t0 24.923
C0 Y B 0.23fF
C1 Y VPWR 0.63fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__nand2b_4.ext - technology: sky130A

.subckt sky130_fd_sc_hd__nand2b_4 B A_N Y VGND VPWR VNB VPB
X0 VGND.t4 B.t0 a_215_47.t2 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 Y.t3 B.t1 VPWR.t4 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 Y.t4 a_27_47.t2 a_215_47.t4 VNB.t5 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 VGND.t3 B.t2 a_215_47.t1 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 Y.t5 a_27_47.t3 a_215_47.t5 VNB.t6 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 a_215_47.t6 a_27_47.t4 Y.t6 VNB.t7 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 a_215_47.t0 B.t3 VGND.t2 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 VPWR.t3 B.t4 Y.t2 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 VPWR.t5 a_27_47.t5 Y.t7 VPB.t5 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 Y.t1 B.t5 VPWR.t2 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 VPWR.t1 B.t6 Y.t0 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 Y.t8 a_27_47.t6 VPWR.t6 VPB.t6 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 VPWR.t7 a_27_47.t7 Y.t9 VPB.t7 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13 a_215_47.t3 B.t7 VGND.t1 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14 a_215_47.t7 a_27_47.t8 Y.t10 VNB.t8 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X15 Y.t11 a_27_47.t9 VPWR.t8 VPB.t8 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16 VPWR.t0 A_N.t0 a_27_47.t1 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17 VGND.t0 A_N.t1 a_27_47.t0 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
R0 B.n0 B.t4 221.719
R1 B.n4 B.t5 221.719
R2 B.n7 B.t6 221.719
R3 B.n8 B.t1 221.719
R4 B.n0 B.t3 149.419
R5 B.n4 B.t2 149.419
R6 B.n7 B.t7 149.419
R7 B.n8 B.t0 149.419
R8 B.n1 B.n0 118.844
R9 B B.n9 80.48
R10 B.n3 B.n2 76
R11 B.n6 B.n5 76
R12 B.n3 B.n0 38.381
R13 B.n9 B.n8 38.381
R14 B.n5 B.n4 37.488
R15 B.n4 B.n3 36.596
R16 B.n9 B.n7 36.596
R17 B B.n6 22.08
R18 B.n2 B 19.2
R19 B B.n1 18.88
R20 B.n1 B 10.56
R21 B.n2 B 10.24
R22 B.n6 B 7.36
R23 a_215_47.t0 a_215_47.n5 139.815
R24 a_215_47.n1 a_215_47.t4 136.83
R25 a_215_47.n1 a_215_47.n0 92.5
R26 a_215_47.n3 a_215_47.n1 55.913
R27 a_215_47.n5 a_215_47.n4 52.818
R28 a_215_47.n5 a_215_47.n3 46.921
R29 a_215_47.n3 a_215_47.n2 42.273
R30 a_215_47.n2 a_215_47.t6 27.692
R31 a_215_47.n2 a_215_47.t2 24.923
R32 a_215_47.n0 a_215_47.t5 24.923
R33 a_215_47.n0 a_215_47.t7 24.923
R34 a_215_47.n4 a_215_47.t1 24.923
R35 a_215_47.n4 a_215_47.t3 24.923
R36 VGND.n14 VGND.t0 200.519
R37 VGND.n3 VGND.n2 118.394
R38 VGND.n1 VGND.n0 114.711
R39 VGND.n2 VGND.t2 24.923
R40 VGND.n2 VGND.t3 24.923
R41 VGND.n0 VGND.t1 24.923
R42 VGND.n0 VGND.t4 24.923
R43 VGND.n3 VGND.n1 14.129
R44 VGND.n5 VGND.n4 4.65
R45 VGND.n7 VGND.n6 4.65
R46 VGND.n9 VGND.n8 4.65
R47 VGND.n11 VGND.n10 4.65
R48 VGND.n13 VGND.n12 4.65
R49 VGND.n15 VGND.n14 4.05
R50 VGND.n5 VGND.n3 0.305
R51 VGND.n15 VGND.n13 0.134
R52 VGND VGND.n15 0.124
R53 VGND.n7 VGND.n5 0.119
R54 VGND.n9 VGND.n7 0.119
R55 VGND.n11 VGND.n9 0.119
R56 VGND.n13 VGND.n11 0.119
R57 VNB VNB.t0 6053.91
R58 VNB.t0 VNB.t5 4545.05
R59 VNB.t7 VNB.t4 2103.3
R60 VNB.t3 VNB.t2 2030.77
R61 VNB.t1 VNB.t3 2030.77
R62 VNB.t4 VNB.t1 2030.77
R63 VNB.t6 VNB.t7 2030.77
R64 VNB.t8 VNB.t6 2030.77
R65 VNB.t5 VNB.t8 2030.77
R66 VPWR.n12 VPWR.n11 174.594
R67 VPWR.n6 VPWR.n5 174.594
R68 VPWR.n1 VPWR.n0 174.594
R69 VPWR.n17 VPWR.t0 172.344
R70 VPWR.n2 VPWR.t3 171.168
R71 VPWR.n17 VPWR.t8 125.866
R72 VPWR.n5 VPWR.t5 29.55
R73 VPWR.n11 VPWR.t6 26.595
R74 VPWR.n11 VPWR.t7 26.595
R75 VPWR.n5 VPWR.t4 26.595
R76 VPWR.n0 VPWR.t2 26.595
R77 VPWR.n0 VPWR.t1 26.595
R78 VPWR.n2 VPWR.n1 17.195
R79 VPWR.n18 VPWR.n17 9.089
R80 VPWR.n7 VPWR.n6 7.152
R81 VPWR.n4 VPWR.n3 4.65
R82 VPWR.n8 VPWR.n7 4.65
R83 VPWR.n10 VPWR.n9 4.65
R84 VPWR.n14 VPWR.n13 4.65
R85 VPWR.n16 VPWR.n15 4.65
R86 VPWR.n13 VPWR.n12 2.258
R87 VPWR.n19 VPWR.n18 2.132
R88 VPWR.n4 VPWR.n2 0.248
R89 VPWR.n19 VPWR.n16 0.191
R90 VPWR VPWR.n19 0.186
R91 VPWR.n8 VPWR.n4 0.119
R92 VPWR.n10 VPWR.n8 0.119
R93 VPWR.n14 VPWR.n10 0.119
R94 VPWR.n16 VPWR.n14 0.119
R95 Y.n9 Y.n4 138.276
R96 Y.n7 Y.n5 138.276
R97 Y.n2 Y.n1 132.322
R98 Y.n7 Y.n6 108.604
R99 Y.n9 Y.n8 108.133
R100 Y.n2 Y.n0 92.5
R101 Y.n9 Y.n7 29.672
R102 Y.n8 Y.t7 26.595
R103 Y.n8 Y.t8 26.595
R104 Y.n5 Y.t2 26.595
R105 Y.n5 Y.t1 26.595
R106 Y.n6 Y.t0 26.595
R107 Y.n6 Y.t3 26.595
R108 Y.n4 Y.t9 26.595
R109 Y.n4 Y.t11 26.595
R110 Y.n0 Y.t6 24.923
R111 Y.n0 Y.t5 24.923
R112 Y.n1 Y.t10 24.923
R113 Y.n1 Y.t4 24.923
R114 Y Y.n3 9.66
R115 Y.n3 Y 6.762
R116 Y Y.n9 4.081
R117 Y.n3 Y 1.659
R118 Y Y.n2 0.474
R119 VPB.t0 VPB.t8 556.386
R120 VPB.t5 VPB.t4 257.476
R121 VPB.t2 VPB.t3 248.598
R122 VPB.t1 VPB.t2 248.598
R123 VPB.t4 VPB.t1 248.598
R124 VPB.t6 VPB.t5 248.598
R125 VPB.t7 VPB.t6 248.598
R126 VPB.t8 VPB.t7 248.598
R127 VPB VPB.t0 189.408
R128 a_27_47.n0 a_27_47.t5 221.719
R129 a_27_47.n1 a_27_47.t6 221.719
R130 a_27_47.n3 a_27_47.t7 221.719
R131 a_27_47.n6 a_27_47.t9 221.719
R132 a_27_47.t1 a_27_47.n8 163.548
R133 a_27_47.n0 a_27_47.t4 149.419
R134 a_27_47.n1 a_27_47.t3 149.419
R135 a_27_47.n3 a_27_47.t8 149.419
R136 a_27_47.n6 a_27_47.t2 149.419
R137 a_27_47.n8 a_27_47.t0 122.808
R138 a_27_47.n7 a_27_47.n6 118.844
R139 a_27_47.n5 a_27_47.n2 102.88
R140 a_27_47.n5 a_27_47.n4 76
R141 a_27_47.n1 a_27_47.n0 74.977
R142 a_27_47.n2 a_27_47.n1 37.488
R143 a_27_47.n4 a_27_47.n3 37.488
R144 a_27_47.n8 a_27_47.n7 30.4
R145 a_27_47.n7 a_27_47.n5 28.8
R146 A_N.n0 A_N.t0 234.572
R147 A_N.n0 A_N.t1 162.272
R148 A_N A_N.n0 84
C0 VPWR Y 1.33fF
C1 VPWR VGND 0.11fF
C2 Y B 0.24fF
C3 VPWR VPB 0.11fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__nand3_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__nand3_1 Y A C B VGND VPWR VNB VPB
X0 VPWR.t0 B.t0 Y.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 Y.t1 A.t0 VPWR.t1 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 a_193_47.t1 B.t1 a_109_47.t0 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 Y.t2 A.t1 a_193_47.t0 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 Y.t3 C.t0 VPWR.t2 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 a_109_47.t1 C.t1 VGND.t0 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
R0 B.n0 B.t0 241.534
R1 B.n0 B.t1 169.234
R2 B B.n0 77.877
R3  B 11.605
R4 Y.n1 Y.t1 177.147
R5 Y Y.t2 123.196
R6 Y.n1 Y.n0 107.635
R7 Y Y.n1 67.484
R8 Y.n0 Y.t0 26.595
R9 Y.n0 Y.t3 26.595
R10 VPWR.n1 VPWR.n0 175.651
R11 VPWR.n1 VPWR.t2 156.096
R12 VPWR.n0 VPWR.t1 38.415
R13 VPWR.n0 VPWR.t0 26.595
R14 VPWR VPWR.n1 0.115
R15 VPB.t0 VPB.t1 284.112
R16 VPB.t2 VPB.t0 248.598
R17 VPB VPB.t2 189.408
R18 A.n0 A.t0 232.213
R19 A.n0 A.t1 159.913
R20 A A.n0 78.27
R21 a_109_47.t0 a_109_47.t1 49.846
R22 a_193_47.t0 a_193_47.t1 60.923
R23 VNB VNB.t2 6053.91
R24 VNB.t1 VNB.t0 2320.88
R25 VNB.t2 VNB.t1 2030.77
R26 C.n0 C.t0 230.361
R27 C.n0 C.t1 158.061
R28 C C.n0 79.2
R29  C 19.781
R30 VGND VGND.t0 186.361
C0 B Y 0.30fF
C1 Y VGND 0.25fF
C2 A Y 0.12fF
C3 VPWR Y 0.56fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__nand3_2.ext - technology: sky130A

.subckt sky130_fd_sc_hd__nand3_2 A Y B C VGND VPWR VNB VPB
X0 VGND.t1 C.t0 a_277_47.t2 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 VPWR.t3 B.t0 Y.t3 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 a_277_47.t1 C.t1 VGND.t0 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 Y.t2 B.t1 VPWR.t2 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 VPWR.t4 A.t0 Y.t4 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 a_27_47.t1 A.t1 Y.t5 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 a_27_47.t3 B.t2 a_277_47.t0 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 VPWR.t1 C.t2 Y.t1 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 Y.t0 C.t3 VPWR.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 a_277_47.t3 B.t3 a_27_47.t2 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 Y.t6 A.t2 VPWR.t5 VPB.t5 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 Y.t7 A.t3 a_27_47.t0 VNB.t5 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
R0 C.n1 C.t2 237.931
R1 C.n2 C.t3 218.506
R2 C.n1 C.t0 166.508
R3 C.n2 C.t1 146.206
R4 C.n1 C.n0 76
R5 C.n4 C.n3 76
R6 C.n3 C.n1 42.382
R7 C C.n4 18.56
R8 C.n0 C 16
R9 C.n3 C.n2 14.958
R10 C.n0 C 13.12
R11 C.n4 C 10.88
R12 a_277_47.n1 a_277_47.n0 249.474
R13 a_277_47.n0 a_277_47.t2 24.923
R14 a_277_47.n0 a_277_47.t1 24.923
R15 a_277_47.t0 a_277_47.n1 24.923
R16 a_277_47.n1 a_277_47.t3 24.923
R17 VGND.n0 VGND.t0 193.592
R18 VGND.n0 VGND.t1 96.127
R19 VGND VGND.n0 0.7
R20 VNB VNB.t5 6053.91
R21 VNB.t0 VNB.t1 4545.05
R22 VNB.t1 VNB.t2 2030.77
R23 VNB.t3 VNB.t0 2030.77
R24 VNB.t4 VNB.t3 2030.77
R25 VNB.t5 VNB.t4 2030.77
R26 B.n0 B.t0 218.506
R27 B.n1 B.t1 218.506
R28 B.n0 B.t2 146.206
R29 B.n1 B.t3 146.206
R30 B.n4 B.n0 90.958
R31 B.n3 B.n2 76
R32 B.n2 B.n0 64.82
R33 B.n4 B 18.56
R34 B.n3 B 17.28
R35 B B.n3 12.16
R36 B B.n4 10.88
R37 B.n2 B.n1 4.986
R38 Y.n2 Y.n0 168.531
R39 Y.n4 Y.n3 108.604
R40 Y.n2 Y.n1 108.604
R41 Y Y.n5 94.245
R42 Y.n4 Y.n2 29.672
R43 Y.n3 Y.t4 26.595
R44 Y.n3 Y.t6 26.595
R45 Y.n0 Y.t1 26.595
R46 Y.n0 Y.t0 26.595
R47 Y.n1 Y.t3 26.595
R48 Y.n1 Y.t2 26.595
R49 Y.n5 Y.t5 24.923
R50 Y.n5 Y.t7 24.923
R51 Y Y.n4 4.266
R52 VPWR.n6 VPWR.n5 174.594
R53 VPWR.n0 VPWR.t3 172.846
R54 VPWR.n0 VPWR.t0 172.846
R55 VPWR.n2 VPWR.t1 152.947
R56 VPWR.n11 VPWR.t5 152.162
R57 VPWR.n5 VPWR.t2 26.595
R58 VPWR.n5 VPWR.t4 26.595
R59 VPWR.n1 VPWR.n0 8.593
R60 VPWR.n4 VPWR.n3 4.65
R61 VPWR.n8 VPWR.n7 4.65
R62 VPWR.n10 VPWR.n9 4.65
R63 VPWR.n12 VPWR.n11 4.65
R64 VPWR.n7 VPWR.n6 3.764
R65 VPWR.n2 VPWR.n1 2.105
R66 VPWR.n4 VPWR.n2 0.238
R67 VPWR.n8 VPWR.n4 0.119
R68 VPWR.n10 VPWR.n8 0.119
R69 VPWR.n12 VPWR.n10 0.119
R70 VPWR VPWR.n12 0.02
R71 VPB.t3 VPB.t0 556.386
R72 VPB.t0 VPB.t1 248.598
R73 VPB.t2 VPB.t3 248.598
R74 VPB.t4 VPB.t2 248.598
R75 VPB.t5 VPB.t4 248.598
R76 VPB VPB.t5 189.408
R77 A.n0 A.t0 212.079
R78 A.n1 A.t2 212.079
R79 A.n0 A.t1 139.779
R80 A.n1 A.t3 139.779
R81 A A.n1 112.547
R82 A.n1 A.n0 61.345
R83 a_27_47.n0 a_27_47.t3 238.823
R84 a_27_47.n0 a_27_47.t0 180.795
R85 a_27_47.n1 a_27_47.n0 92.5
R86 a_27_47.n1 a_27_47.t2 24.923
R87 a_27_47.t1 a_27_47.n1 24.923
C0 B Y 0.31fF
C1 C Y 0.11fF
C2 VPWR Y 1.16fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__nand3_4.ext - technology: sky130A

.subckt sky130_fd_sc_hd__nand3_4 Y A B C VGND VPWR VNB VPB
X0 a_27_47.t3 B.t0 a_445_47.t3 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 a_27_47.t2 B.t1 a_445_47.t2 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 Y.t3 B.t2 VPWR.t3 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 VPWR.t8 C.t0 Y.t12 VPB.t8 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 Y.t4 A.t0 a_445_47.t4 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 Y.t13 C.t1 VPWR.t9 VPB.t9 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 Y.t5 A.t1 a_445_47.t5 VNB.t5 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 VPWR.t10 C.t2 Y.t14 VPB.t10 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 a_27_47.t4 C.t3 VGND.t3 VNB.t8 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 a_27_47.t5 C.t4 VGND.t2 VNB.t9 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 a_445_47.t6 A.t2 Y.t6 VNB.t6 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 VPWR.t2 B.t3 Y.t2 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 a_445_47.t7 A.t3 Y.t7 VNB.t7 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 VGND.t1 C.t5 a_27_47.t6 VNB.t10 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14 a_445_47.t1 B.t4 a_27_47.t1 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X15 Y.t1 B.t5 VPWR.t1 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16 VPWR.t4 A.t4 Y.t8 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17 a_445_47.t0 B.t6 a_27_47.t0 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X18 VPWR.t0 B.t7 Y.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X19 Y.t9 A.t5 VPWR.t5 VPB.t5 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X20 VPWR.t6 A.t6 Y.t10 VPB.t6 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X21 Y.t15 C.t6 VPWR.t11 VPB.t11 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X22 Y.t11 A.t7 VPWR.t7 VPB.t7 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X23 VGND.t0 C.t7 a_27_47.t7 VNB.t11 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
R0 B.n1 B.t3 221.719
R1 B.n0 B.t5 221.719
R2 B.n6 B.t7 221.719
R3 B.n7 B.t2 221.719
R4 B.n1 B.t1 149.419
R5 B.n0 B.t6 149.419
R6 B.n6 B.t0 149.419
R7 B.n7 B.t4 149.419
R8 B.n3 B.n2 76
R9 B.n5 B.n4 76
R10 B.n9 B.n8 76
R11 B.n2 B.n1 37.488
R12 B.n2 B.n0 37.488
R13 B.n5 B.n0 37.488
R14 B.n6 B.n5 37.488
R15 B.n8 B.n6 37.488
R16 B.n8 B.n7 37.488
R17 B B.n9 23.68
R18 B.n4 B 21.12
R19 B B.n3 18.56
R20 B.n3 B 10.88
R21 B.n4 B 8.32
R22 B.n9 B 5.76
R23 a_445_47.n1 a_445_47.t6 210.358
R24 a_445_47.n2 a_445_47.t5 166.346
R25 a_445_47.n4 a_445_47.n3 139.247
R26 a_445_47.n1 a_445_47.n0 92.5
R27 a_445_47.n5 a_445_47.n4 92.5
R28 a_445_47.n4 a_445_47.n2 52.313
R29 a_445_47.n2 a_445_47.n1 46.747
R30 a_445_47.n3 a_445_47.t3 24.923
R31 a_445_47.n3 a_445_47.t1 24.923
R32 a_445_47.n0 a_445_47.t4 24.923
R33 a_445_47.n0 a_445_47.t7 24.923
R34 a_445_47.n5 a_445_47.t2 24.923
R35 a_445_47.t0 a_445_47.n5 24.923
R36 a_27_47.n4 a_27_47.t2 230.872
R37 a_27_47.n2 a_27_47.t7 130.175
R38 a_27_47.n3 a_27_47.n0 92.5
R39 a_27_47.n5 a_27_47.n4 92.5
R40 a_27_47.n4 a_27_47.n3 55.296
R41 a_27_47.n2 a_27_47.n1 52.431
R42 a_27_47.n3 a_27_47.n2 46.848
R43 a_27_47.n0 a_27_47.t1 24.923
R44 a_27_47.n0 a_27_47.t5 24.923
R45 a_27_47.n1 a_27_47.t6 24.923
R46 a_27_47.n1 a_27_47.t4 24.923
R47 a_27_47.n5 a_27_47.t0 24.923
R48 a_27_47.t3 a_27_47.n5 24.923
R49 VNB VNB.t11 6053.91
R50 VNB.t2 VNB.t5 4545.05
R51 VNB.t4 VNB.t6 2030.77
R52 VNB.t7 VNB.t4 2030.77
R53 VNB.t5 VNB.t7 2030.77
R54 VNB.t0 VNB.t2 2030.77
R55 VNB.t3 VNB.t0 2030.77
R56 VNB.t1 VNB.t3 2030.77
R57 VNB.t9 VNB.t1 2030.77
R58 VNB.t10 VNB.t9 2030.77
R59 VNB.t8 VNB.t10 2030.77
R60 VNB.t11 VNB.t8 2030.77
R61 VPWR.n0 VPWR.t4 198.311
R62 VPWR.n25 VPWR.n24 174.594
R63 VPWR.n19 VPWR.n18 174.594
R64 VPWR.n13 VPWR.n12 174.594
R65 VPWR.n2 VPWR.n1 174.594
R66 VPWR.n7 VPWR.t2 172.846
R67 VPWR.n7 VPWR.t7 172.846
R68 VPWR.n30 VPWR.t11 152.162
R69 VPWR.n24 VPWR.t9 26.595
R70 VPWR.n24 VPWR.t10 26.595
R71 VPWR.n18 VPWR.t3 26.595
R72 VPWR.n18 VPWR.t8 26.595
R73 VPWR.n12 VPWR.t1 26.595
R74 VPWR.n12 VPWR.t0 26.595
R75 VPWR.n1 VPWR.t5 26.595
R76 VPWR.n1 VPWR.t6 26.595
R77 VPWR.n14 VPWR.n13 15.811
R78 VPWR.n3 VPWR.n2 11.294
R79 VPWR.n20 VPWR.n19 9.788
R80 VPWR.n8 VPWR.n7 8.593
R81 VPWR.n4 VPWR.n3 4.65
R82 VPWR.n6 VPWR.n5 4.65
R83 VPWR.n9 VPWR.n8 4.65
R84 VPWR.n11 VPWR.n10 4.65
R85 VPWR.n15 VPWR.n14 4.65
R86 VPWR.n17 VPWR.n16 4.65
R87 VPWR.n21 VPWR.n20 4.65
R88 VPWR.n23 VPWR.n22 4.65
R89 VPWR.n27 VPWR.n26 4.65
R90 VPWR.n29 VPWR.n28 4.65
R91 VPWR.n31 VPWR.n30 4.65
R92 VPWR.n26 VPWR.n25 3.764
R93 VPWR.n4 VPWR.n0 0.552
R94 VPWR.n6 VPWR.n4 0.119
R95 VPWR.n9 VPWR.n6 0.119
R96 VPWR.n11 VPWR.n9 0.119
R97 VPWR.n15 VPWR.n11 0.119
R98 VPWR.n17 VPWR.n15 0.119
R99 VPWR.n21 VPWR.n17 0.119
R100 VPWR.n23 VPWR.n21 0.119
R101 VPWR.n27 VPWR.n23 0.119
R102 VPWR.n29 VPWR.n27 0.119
R103 VPWR.n31 VPWR.n29 0.119
R104 VPWR VPWR.n31 0.02
R105 Y.n5 Y.n3 138.276
R106 Y.n2 Y.n1 135.508
R107 Y.n5 Y.n4 108.604
R108 Y.n7 Y.n6 108.604
R109 Y.n9 Y.n8 108.604
R110 Y.n11 Y.n10 108.604
R111 Y.n13 Y.n12 108.604
R112 Y.n2 Y.n0 92.5
R113 Y.n11 Y.n9 59.927
R114 Y Y.n13 38.702
R115 Y Y.n2 37.12
R116 Y.n7 Y.n5 29.672
R117 Y.n9 Y.n7 29.672
R118 Y.n13 Y.n11 29.672
R119 Y.n3 Y.t14 26.595
R120 Y.n3 Y.t15 26.595
R121 Y.n4 Y.t12 26.595
R122 Y.n4 Y.t13 26.595
R123 Y.n6 Y.t0 26.595
R124 Y.n6 Y.t3 26.595
R125 Y.n8 Y.t2 26.595
R126 Y.n8 Y.t1 26.595
R127 Y.n10 Y.t10 26.595
R128 Y.n10 Y.t11 26.595
R129 Y.n12 Y.t8 26.595
R130 Y.n12 Y.t9 26.595
R131 Y.n0 Y.t6 24.923
R132 Y.n0 Y.t4 24.923
R133 Y.n1 Y.t7 24.923
R134 Y.n1 Y.t5 24.923
R135 Y.n14 Y 11.13
R136 Y Y.n14 7.791
R137 Y.n14 Y 5.888
R138 VPB.t2 VPB.t7 556.386
R139 VPB.t5 VPB.t4 248.598
R140 VPB.t6 VPB.t5 248.598
R141 VPB.t7 VPB.t6 248.598
R142 VPB.t1 VPB.t2 248.598
R143 VPB.t0 VPB.t1 248.598
R144 VPB.t3 VPB.t0 248.598
R145 VPB.t8 VPB.t3 248.598
R146 VPB.t9 VPB.t8 248.598
R147 VPB.t10 VPB.t9 248.598
R148 VPB.t11 VPB.t10 248.598
R149 VPB VPB.t11 189.408
R150 C.n9 C.t6 234.572
R151 C.n2 C.t0 221.719
R152 C.n4 C.t1 221.719
R153 C.n0 C.t2 221.719
R154 C.n9 C.t7 162.272
R155 C.n2 C.t4 149.419
R156 C.n4 C.t5 149.419
R157 C.n0 C.t3 149.419
R158 C.n6 C.n5 76
R159 C.n8 C.n7 76
R160 C.n10 C.n9 76
R161 C.n3 C.n2 37.488
R162 C.n4 C.n3 37.488
R163 C.n5 C.n4 37.488
R164 C.n5 C.n0 37.488
R165 C.n8 C.n0 37.488
R166 C.n6 C.n1 26.88
R167 C.n7 C 24.96
R168 C.n9 C.n8 24.1
R169 C.n10 C 21.44
R170 C C.n10 8
R171 C.n7 C 4.48
R172 C C.n6 1.92
R173 C.n1 C 0.64
R174 A.n1 A.t4 221.719
R175 A.n3 A.t5 221.719
R176 A.n0 A.t6 221.719
R177 A.n8 A.t7 221.719
R178 A.n1 A.t2 149.419
R179 A.n3 A.t0 149.419
R180 A.n0 A.t3 149.419
R181 A.n8 A.t1 149.419
R182 A.n9 A.n8 118.844
R183 A.n2 A 86.88
R184 A.n5 A.n4 76
R185 A.n7 A.n6 76
R186 A.n7 A.n0 38.381
R187 A.n2 A.n1 37.488
R188 A.n3 A.n2 37.488
R189 A.n4 A.n3 37.488
R190 A.n4 A.n0 37.488
R191 A.n8 A.n7 36.596
R192 A A.n9 16.64
R193 A.n5 A 16
R194 A.n6 A 15.68
R195 A.n6 A 13.76
R196 A A.n5 13.44
R197 A.n9 A 12.8
R198 VGND.n2 VGND.n0 124.436
R199 VGND.n2 VGND.n1 120.435
R200 VGND.n0 VGND.t2 24.923
R201 VGND.n0 VGND.t1 24.923
R202 VGND.n1 VGND.t3 24.923
R203 VGND.n1 VGND.t0 24.923
R204 VGND VGND.n2 0.249
C0 VPWR Y 2.16fF
C1 C Y 0.23fF
C2 VPWR VGND 0.14fF
C3 B Y 0.42fF
C4 VPB VPWR 0.14fF
C5 A Y 0.68fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__nand3b_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__nand3b_1 B C A_N Y VGND VPWR VNB VPB
X0 Y.t0 a_53_93.t2 VPWR.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_232_47.t0 C.t0 VGND.t0 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 VPWR.t1 B.t0 Y.t2 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 VPWR.t3 A_N.t0 a_53_93.t0 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 VGND.t1 A_N.t1 a_53_93.t1 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 a_316_47.t1 B.t1 a_232_47.t1 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 Y.t1 a_53_93.t3 a_316_47.t0 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 Y.t3 C.t1 VPWR.t2 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
R0 a_53_93.t0 a_53_93.n1 429.74
R1 a_53_93.n0 a_53_93.t2 236.179
R2 a_53_93.n1 a_53_93.n0 227.241
R3 a_53_93.n0 a_53_93.t3 163.879
R4 a_53_93.n1 a_53_93.t1 131.071
R5 VPWR.n2 VPWR.n0 171.325
R6 VPWR.n2 VPWR.n1 130.646
R7 VPWR.n1 VPWR.t3 95.417
R8 VPWR.n0 VPWR.t1 38.415
R9 VPWR.n0 VPWR.t0 37.43
R10 VPWR.n1 VPWR.t2 26.336
R11 VPWR VPWR.n2 0.248
R12 Y.n4 Y.n3 292.5
R13 Y Y.t1 179.582
R14 Y.n2 Y.n0 154.693
R15 Y.n5 Y.n4 146.679
R16 Y.n4 Y.t0 26.595
R17 Y.n0 Y.t2 26.595
R18 Y.n0 Y.t3 26.595
R19 Y.n5 Y 5.948
R20 Y.n3 Y 2.82
R21 Y.n1 Y 2.206
R22 Y.n2 Y.n1 1.844
R23 Y.n3 Y.n2 1.627
R24 Y Y.n5 1.415
R25 Y.n1 Y 1.084
R26 VPB.t1 VPB.t0 316.666
R27 VPB.t3 VPB.t2 287.071
R28 VPB VPB.t3 269.314
R29 VPB.t2 VPB.t1 248.598
R30 C.n0 C.t1 236.179
R31 C.n0 C.t0 163.879
R32 C C.n0 78.607
R33 VGND VGND.n0 113.875
R34 VGND.n0 VGND.t1 58.571
R35 VGND.n0 VGND.t0 24
R36 a_232_47.t0 a_232_47.t1 49.846
R37 VNB VNB.t3 6706.66
R38 VNB.t2 VNB.t0 2586.81
R39 VNB.t3 VNB.t1 2345.05
R40 VNB.t1 VNB.t2 2030.77
R41 B.n0 B.t0 236.179
R42 B.n0 B.t1 163.879
R43 B B.n0 78.521
R44 A_N.n0 A_N.t0 142.993
R45 A_N.n0 A_N.t1 126.926
R46 A_N A_N.n0 79.684
R47 a_316_47.t0 a_316_47.t1 71.076
C0 C B 0.11fF
C1 Y VGND 0.11fF
C2 VPWR Y 0.57fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__nand3b_2.ext - technology: sky130A

.subckt sky130_fd_sc_hd__nand3b_2 Y C A_N B VGND VPWR VNB VPB
X0 a_408_47.t1 B.t0 a_218_47.t1 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 a_408_47.t2 a_27_47.t2 Y.t5 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 Y.t4 a_27_47.t3 a_408_47.t3 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 VPWR.t2 A_N.t0 a_27_47.t0 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 VGND.t2 C.t0 a_218_47.t2 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 VPWR.t1 B.t1 Y.t1 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 a_218_47.t3 C.t1 VGND.t1 VNB.t5 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 Y.t0 B.t2 VPWR.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 VPWR.t3 C.t2 Y.t2 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 VPWR.t6 a_27_47.t4 Y.t7 VPB.t6 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 a_218_47.t0 B.t3 a_408_47.t0 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 Y.t3 C.t3 VPWR.t4 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 Y.t6 a_27_47.t5 VPWR.t5 VPB.t5 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13 VGND.t0 A_N.t1 a_27_47.t1 VNB.t6 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
R0 B.n4 B.t2 268.133
R1 B.n3 B.t1 221.719
R2 B.n1 B.t0 206.544
R3 B.n2 B.t3 149.419
R4 B.n1 B.n0 76
R5 B.n5 B.n4 76
R6 B.n0  29.12
R7 B.n4 B.n3 28.562
R8 B.n5  21.44
R9 B.n2 B.n1 17.851
R10 B.n3 B.n2 17.851
R11 B B.n5 2.56
R12 B.n0  1.6
R13 a_218_47.n1 a_218_47.n0 214.145
R14 a_218_47.n0 a_218_47.t2 24.923
R15 a_218_47.n0 a_218_47.t3 24.923
R16 a_218_47.n1 a_218_47.t1 24.923
R17 a_218_47.t0 a_218_47.n1 24.923
R18 a_408_47.n0 a_408_47.t2 226.776
R19 a_408_47.n0 a_408_47.t0 226.776
R20 a_408_47.n1 a_408_47.n0 50.6
R21 a_408_47.n1 a_408_47.t3 24.923
R22 a_408_47.t1 a_408_47.n1 24.923
R23 VNB VNB.t6 6438.23
R24 VNB.t4 VNB.t0 4545.05
R25 VNB.t6 VNB.t5 2593.81
R26 VNB.t3 VNB.t2 2030.77
R27 VNB.t1 VNB.t3 2030.77
R28 VNB.t0 VNB.t1 2030.77
R29 VNB.t5 VNB.t4 2030.77
R30 a_27_47.t0 a_27_47.n3 399.103
R31 a_27_47.n3 a_27_47.n2 327.151
R32 a_27_47.n0 a_27_47.t4 221.719
R33 a_27_47.n1 a_27_47.t5 221.719
R34 a_27_47.n3 a_27_47.t1 199.953
R35 a_27_47.n0 a_27_47.t2 149.419
R36 a_27_47.n1 a_27_47.t3 149.419
R37 a_27_47.n2 a_27_47.n1 48.2
R38 a_27_47.n2 a_27_47.n0 26.777
R39 Y.n3 Y.n1 183.219
R40 Y.n4 Y.n0 153.805
R41 Y.n3 Y.n2 153.547
R42 Y Y.n5 130.188
R43 Y.n4 Y.n3 79.801
R44 Y Y.n4 47.36
R45 Y.n0 Y.t7 26.595
R46 Y.n0 Y.t6 26.595
R47 Y.n2 Y.t1 26.595
R48 Y.n2 Y.t0 26.595
R49 Y.n1 Y.t2 26.595
R50 Y.n1 Y.t3 26.595
R51 Y.n5 Y.t5 24.923
R52 Y.n5 Y.t4 24.923
R53 A_N.n0 A_N.t0 329.006
R54 A_N.n0 A_N.t1 200.473
R55 A_N A_N.n0 78.011
R56 VPWR.n1 VPWR.t6 582.327
R57 VPWR.n0 VPWR.t5 580.936
R58 VPWR.n2 VPWR.t1 580.936
R59 VPWR.n7 VPWR.n6 314.711
R60 VPWR.n13 VPWR.n12 164.157
R61 VPWR.n12 VPWR.t2 101.464
R62 VPWR.n12 VPWR.t4 39.853
R63 VPWR.n6 VPWR.t0 26.595
R64 VPWR.n6 VPWR.t3 26.595
R65 VPWR.n3 VPWR.n2 4.65
R66 VPWR.n5 VPWR.n4 4.65
R67 VPWR.n9 VPWR.n8 4.65
R68 VPWR.n11 VPWR.n10 4.65
R69 VPWR.n14 VPWR.n13 4.031
R70 VPWR.n1 VPWR.n0 3.944
R71 VPWR.n8 VPWR.n7 2.635
R72 VPWR.n3 VPWR.n1 0.223
R73 VPWR.n14 VPWR.n11 0.135
R74 VPWR VPWR.n14 0.124
R75 VPWR.n5 VPWR.n3 0.119
R76 VPWR.n9 VPWR.n5 0.119
R77 VPWR.n11 VPWR.n9 0.119
R78 VPB.t1 VPB.t5 556.386
R79 VPB.t2 VPB.t4 322.585
R80 VPB.t5 VPB.t6 248.598
R81 VPB.t0 VPB.t1 248.598
R82 VPB.t3 VPB.t0 248.598
R83 VPB.t4 VPB.t3 248.598
R84 VPB VPB.t2 189.408
R85 C.n0 C.t2 221.719
R86 C.n1 C.t3 221.719
R87 C.n0 C.t0 149.419
R88 C.n1 C.t1 149.419
R89 C.n3 C.n2 76
R90 C.n2 C.n0 37.488
R91 C.n2 C.n1 37.488
R92  C.n3 19.52
R93 C.n3 C 9.92
R94 VGND.n1 VGND.t2 198.672
R95 VGND.n1 VGND.n0 69.837
R96 VGND.n0 VGND.t0 61.212
R97 VGND.n0 VGND.t1 35.029
R98 VGND VGND.n1 0.212
C0 VPWR Y 0.72fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__nand3b_4.ext - technology: sky130A

.subckt sky130_fd_sc_hd__nand3b_4 A_N Y B C VGND VPWR VNB VPB
X0 VGND.t4 C.t0 a_633_47.t3 VNB.t8 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 Y.t11 B.t0 VPWR.t7 VPB.t7 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 Y.t0 a_27_47.t2 a_215_47.t7 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 Y.t1 a_27_47.t3 a_215_47.t6 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 a_633_47.t5 B.t1 a_215_47.t3 VNB.t10 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 VPWR.t6 B.t2 Y.t10 VPB.t6 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 Y.t15 C.t1 VPWR.t12 VPB.t12 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 a_633_47.t6 B.t3 a_215_47.t2 VNB.t11 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 VPWR.t11 C.t2 Y.t14 VPB.t11 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 a_215_47.t5 a_27_47.t4 Y.t2 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 Y.t13 C.t3 VPWR.t10 VPB.t10 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 a_215_47.t1 B.t4 a_633_47.t7 VNB.t12 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 a_215_47.t0 B.t5 a_633_47.t4 VNB.t9 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 Y.t9 B.t6 VPWR.t5 VPB.t5 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14 VPWR.t0 a_27_47.t5 Y.t3 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 Y.t4 a_27_47.t6 VPWR.t1 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16 a_633_47.t2 C.t4 VGND.t3 VNB.t7 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X17 a_633_47.t1 C.t5 VGND.t2 VNB.t6 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X18 VPWR.t2 a_27_47.t7 Y.t5 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X19 VPWR.t9 C.t6 Y.t12 VPB.t9 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X20 a_215_47.t4 a_27_47.t8 Y.t6 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X21 Y.t7 a_27_47.t9 VPWR.t3 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X22 VPWR.t8 A_N.t0 a_27_47.t0 VPB.t8 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X23 VGND.t1 C.t7 a_633_47.t0 VNB.t5 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X24 VPWR.t4 B.t7 Y.t8 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X25 VGND.t0 A_N.t1 a_27_47.t1 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
R0 C.n0 C.t6 221.719
R1 C.n1 C.t1 221.719
R2 C.n7 C.t2 221.719
R3 C.n3 C.t3 221.719
R4 C.n0 C.t0 149.419
R5 C.n1 C.t5 149.419
R6 C.n7 C.t7 149.419
R7 C.n3 C.t4 149.419
R8 C.n4 C.n3 118.844
R9 C C.n2 86.56
R10 C.n9 C.n8 76
R11 C.n6 C.n5 76
R12 C.n2 C.n0 38.381
R13 C.n8 C.n7 37.488
R14 C.n7 C.n6 37.488
R15 C.n6 C.n3 37.488
R16 C.n2 C.n1 36.596
R17 C.n4 C 16.64
R18 C C.n9 16
R19 C.n5 C 16
R20 C.n9 C 13.44
R21 C.n5 C 13.44
R22 C C.n4 12.8
R23 a_633_47.n2 a_633_47.n1 132.322
R24 a_633_47.n2 a_633_47.n0 92.5
R25 a_633_47.n4 a_633_47.n3 87.175
R26 a_633_47.n4 a_633_47.n2 68.827
R27 a_633_47.n5 a_633_47.n4 52.817
R28 a_633_47.n3 a_633_47.t3 24.923
R29 a_633_47.n3 a_633_47.t1 24.923
R30 a_633_47.n1 a_633_47.t7 24.923
R31 a_633_47.n1 a_633_47.t5 24.923
R32 a_633_47.n0 a_633_47.t4 24.923
R33 a_633_47.n0 a_633_47.t6 24.923
R34 a_633_47.t0 a_633_47.n5 24.923
R35 a_633_47.n5 a_633_47.t2 24.923
R36 VGND.n7 VGND.t3 195.032
R37 VGND.n26 VGND.t0 195.032
R38 VGND.n2 VGND.n1 114.711
R39 VGND.n0 VGND.t4 106.913
R40 VGND.n1 VGND.t2 24.923
R41 VGND.n1 VGND.t1 24.923
R42 VGND.n3 VGND.n2 12.8
R43 VGND.n8 VGND.n7 6.4
R44 VGND.n4 VGND.n3 4.65
R45 VGND.n6 VGND.n5 4.65
R46 VGND.n9 VGND.n8 4.65
R47 VGND.n11 VGND.n10 4.65
R48 VGND.n13 VGND.n12 4.65
R49 VGND.n15 VGND.n14 4.65
R50 VGND.n17 VGND.n16 4.65
R51 VGND.n19 VGND.n18 4.65
R52 VGND.n21 VGND.n20 4.65
R53 VGND.n23 VGND.n22 4.65
R54 VGND.n25 VGND.n24 4.65
R55 VGND.n27 VGND.n26 4.05
R56 VGND.n4 VGND.n0 0.505
R57 VGND.n27 VGND.n25 0.134
R58 VGND VGND.n27 0.124
R59 VGND.n6 VGND.n4 0.119
R60 VGND.n9 VGND.n6 0.119
R61 VGND.n11 VGND.n9 0.119
R62 VGND.n13 VGND.n11 0.119
R63 VGND.n15 VGND.n13 0.119
R64 VGND.n17 VGND.n15 0.119
R65 VGND.n19 VGND.n17 0.119
R66 VGND.n21 VGND.n19 0.119
R67 VGND.n23 VGND.n21 0.119
R68 VGND.n25 VGND.n23 0.119
R69 VNB VNB.t4 6053.91
R70 VNB.t9 VNB.t7 4545.05
R71 VNB.t4 VNB.t0 4545.05
R72 VNB.t6 VNB.t8 2030.77
R73 VNB.t5 VNB.t6 2030.77
R74 VNB.t7 VNB.t5 2030.77
R75 VNB.t11 VNB.t9 2030.77
R76 VNB.t12 VNB.t11 2030.77
R77 VNB.t10 VNB.t12 2030.77
R78 VNB.t2 VNB.t10 2030.77
R79 VNB.t1 VNB.t2 2030.77
R80 VNB.t3 VNB.t1 2030.77
R81 VNB.t0 VNB.t3 2030.77
R82 B.n0 B.t7 221.719
R83 B.n3 B.t0 221.719
R84 B.n4 B.t2 221.719
R85 B.n5 B.t6 221.719
R86 B.n0 B.t5 149.419
R87 B.n3 B.t3 149.419
R88 B.n4 B.t4 149.419
R89 B.n5 B.t1 149.419
R90 B.n2 B.n1 76
R91 B.n7 B.n6 76
R92 B.n4 B.n3 74.977
R93 B.n6 B.n5 61.588
R94 B.n2 B.n0 41.951
R95 B.n3 B.n2 33.025
R96 B.n7 B 26.56
R97 B.n1 B 16.96
R98 B.n6 B.n4 13.388
R99 B.n1 B 12.48
R100 B B.n7 2.88
R101 VPWR.n19 VPWR.n18 314.711
R102 VPWR.n2 VPWR.n1 174.594
R103 VPWR.n25 VPWR.n24 174.594
R104 VPWR.n13 VPWR.n12 174.594
R105 VPWR.n7 VPWR.t4 172.846
R106 VPWR.n7 VPWR.t10 172.846
R107 VPWR.n0 VPWR.t9 164.78
R108 VPWR.n30 VPWR.t3 124.097
R109 VPWR.n30 VPWR.t8 124.096
R110 VPWR.n1 VPWR.t12 26.595
R111 VPWR.n1 VPWR.t11 26.595
R112 VPWR.n24 VPWR.t1 26.595
R113 VPWR.n24 VPWR.t2 26.595
R114 VPWR.n18 VPWR.t5 26.595
R115 VPWR.n18 VPWR.t0 26.595
R116 VPWR.n12 VPWR.t7 26.595
R117 VPWR.n12 VPWR.t6 26.595
R118 VPWR.n14 VPWR.n13 14.305
R119 VPWR.n3 VPWR.n2 12.8
R120 VPWR.n31 VPWR.n30 10.419
R121 VPWR.n8 VPWR.n7 8.593
R122 VPWR.n20 VPWR.n19 8.282
R123 VPWR.n4 VPWR.n3 4.65
R124 VPWR.n6 VPWR.n5 4.65
R125 VPWR.n9 VPWR.n8 4.65
R126 VPWR.n11 VPWR.n10 4.65
R127 VPWR.n15 VPWR.n14 4.65
R128 VPWR.n17 VPWR.n16 4.65
R129 VPWR.n21 VPWR.n20 4.65
R130 VPWR.n23 VPWR.n22 4.65
R131 VPWR.n27 VPWR.n26 4.65
R132 VPWR.n29 VPWR.n28 4.65
R133 VPWR.n26 VPWR.n25 2.258
R134 VPWR.n32 VPWR.n31 2.132
R135 VPWR.n4 VPWR.n0 0.505
R136 VPWR.n32 VPWR.n29 0.191
R137 VPWR VPWR.n32 0.186
R138 VPWR.n6 VPWR.n4 0.119
R139 VPWR.n9 VPWR.n6 0.119
R140 VPWR.n11 VPWR.n9 0.119
R141 VPWR.n15 VPWR.n11 0.119
R142 VPWR.n17 VPWR.n15 0.119
R143 VPWR.n21 VPWR.n17 0.119
R144 VPWR.n23 VPWR.n21 0.119
R145 VPWR.n27 VPWR.n23 0.119
R146 VPWR.n29 VPWR.n27 0.119
R147 Y.n9 Y.n8 142.047
R148 Y.n2 Y.n0 138.276
R149 Y.n13 Y.n12 132.322
R150 Y.n2 Y.n1 108.604
R151 Y.n4 Y.n3 108.604
R152 Y.n9 Y.n7 98.902
R153 Y.n6 Y.n5 98.902
R154 Y.n13 Y.n11 92.5
R155 Y.n4 Y.n2 59.927
R156 Y Y.n13 33.97
R157 Y.n6 Y.n4 33.443
R158 Y.n5 Y.t10 26.595
R159 Y.n5 Y.t9 26.595
R160 Y.n7 Y.t3 26.595
R161 Y.n7 Y.t4 26.595
R162 Y.n8 Y.t5 26.595
R163 Y.n8 Y.t7 26.595
R164 Y.n0 Y.t12 26.595
R165 Y.n0 Y.t15 26.595
R166 Y.n1 Y.t14 26.595
R167 Y.n1 Y.t13 26.595
R168 Y.n3 Y.t8 26.595
R169 Y.n3 Y.t11 26.595
R170 Y.n11 Y.t2 24.923
R171 Y.n11 Y.t1 24.923
R172 Y.n12 Y.t6 24.923
R173 Y.n12 Y.t0 24.923
R174 Y Y.n10 14.268
R175 Y Y.n9 10.742
R176 Y.n10 Y.n6 8.114
R177 Y.n10 Y 0.342
R178 VPB.t4 VPB.t10 556.386
R179 VPB.t8 VPB.t3 556.386
R180 VPB.t12 VPB.t9 248.598
R181 VPB.t11 VPB.t12 248.598
R182 VPB.t10 VPB.t11 248.598
R183 VPB.t7 VPB.t4 248.598
R184 VPB.t6 VPB.t7 248.598
R185 VPB.t5 VPB.t6 248.598
R186 VPB.t0 VPB.t5 248.598
R187 VPB.t1 VPB.t0 248.598
R188 VPB.t2 VPB.t1 248.598
R189 VPB.t3 VPB.t2 248.598
R190 VPB VPB.t8 189.408
R191 a_27_47.n0 a_27_47.t5 221.719
R192 a_27_47.n2 a_27_47.t6 221.719
R193 a_27_47.n5 a_27_47.t7 221.719
R194 a_27_47.n8 a_27_47.t9 221.719
R195 a_27_47.t0 a_27_47.n10 182.097
R196 a_27_47.n0 a_27_47.t4 149.419
R197 a_27_47.n2 a_27_47.t3 149.419
R198 a_27_47.n5 a_27_47.t8 149.419
R199 a_27_47.n8 a_27_47.t2 149.419
R200 a_27_47.n9 a_27_47.n8 118.844
R201 a_27_47.n4 a_27_47.n1 102.88
R202 a_27_47.n10 a_27_47.t1 91.728
R203 a_27_47.n7 a_27_47.n6 76
R204 a_27_47.n4 a_27_47.n3 76
R205 a_27_47.n10 a_27_47.n9 55.073
R206 a_27_47.n1 a_27_47.n0 37.488
R207 a_27_47.n3 a_27_47.n2 37.488
R208 a_27_47.n6 a_27_47.n5 37.488
R209 a_27_47.n7 a_27_47.n4 26.88
R210 a_27_47.n9 a_27_47.n7 22.125
R211 a_215_47.n1 a_215_47.t0 226.776
R212 a_215_47.n3 a_215_47.t7 226.776
R213 a_215_47.n1 a_215_47.n0 92.5
R214 a_215_47.n3 a_215_47.n2 92.5
R215 a_215_47.n5 a_215_47.n4 92.5
R216 a_215_47.n4 a_215_47.n1 51.2
R217 a_215_47.n4 a_215_47.n3 51.2
R218 a_215_47.n2 a_215_47.t6 24.923
R219 a_215_47.n2 a_215_47.t4 24.923
R220 a_215_47.n0 a_215_47.t2 24.923
R221 a_215_47.n0 a_215_47.t1 24.923
R222 a_215_47.t3 a_215_47.n5 24.923
R223 a_215_47.n5 a_215_47.t5 24.923
R224 A_N.n0 A_N.t0 237.653
R225 A_N.n0 A_N.t1 165.353
R226 A_N A_N.n0 78.011
C0 B Y 0.37fF
C1 VPB VPWR 0.17fF
C2 C Y 0.45fF
C3 VPWR Y 2.04fF
C4 VGND VPWR 0.19fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__nand4_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__nand4_1 C B Y D A VPWR VGND VNB VPB
X0 Y.t1 B.t0 VPWR.t1 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 VPWR.t3 A.t0 Y.t4 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 VPWR.t2 C.t0 Y.t2 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 a_193_47.t0 C.t1 a_109_47.t0 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 Y.t3 A.t1 a_277_47.t0 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 a_277_47.t1 B.t1 a_193_47.t1 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 Y.t0 D.t0 VPWR.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 a_109_47.t1 D.t1 VGND.t0 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
R0 B.n0 B.t0 241.534
R1 B.n0 B.t1 169.234
R2 B B.n0 108.054
R3 VPWR.n2 VPWR.t3 198.089
R4 VPWR.n1 VPWR.n0 174.594
R5 VPWR.n5 VPWR.t0 151.631
R6 VPWR.n0 VPWR.t1 26.595
R7 VPWR.n0 VPWR.t2 26.595
R8 VPWR.n2 VPWR.n1 7.83
R9 VPWR.n4 VPWR.n3 4.65
R10 VPWR.n6 VPWR.n5 4.65
R11 VPWR.n4 VPWR.n2 0.206
R12 VPWR.n6 VPWR.n4 0.119
R13 VPWR VPWR.n6 0.02
R14 Y.n2 Y.n1 160.716
R15 Y.n2 Y.n0 104.452
R16 Y.n3 Y.t3 86.714
R17 Y.n3 Y.n2 62.494
R18 Y.n0 Y.t4 32.505
R19 Y.n0 Y.t1 32.505
R20 Y.n1 Y.t2 26.595
R21 Y.n1 Y.t0 26.595
R22 Y Y.n3 4.042
R23 VPB.t1 VPB.t3 284.112
R24 VPB.t2 VPB.t1 248.598
R25 VPB.t0 VPB.t2 248.598
R26 VPB VPB.t0 189.408
R27 A.n0 A.t0 228.647
R28 A.n0 A.t1 156.347
R29 A.n1 A.n0 76
R30  A.n1 15.2
R31 A.n1 A 2.933
R32 C.n0 C.t0 241.534
R33 C.n0 C.t1 169.234
R34 C.n1 C.n0 83.369
R35  C.n1 13.693
R36 C.n1 C 3.49
R37 a_109_47.t0 a_109_47.t1 49.846
R38 a_193_47.t0 a_193_47.t1 49.846
R39 VNB VNB.t1 6053.91
R40 VNB.t3 VNB.t2 2320.88
R41 VNB.t0 VNB.t3 2030.77
R42 VNB.t1 VNB.t0 2030.77
R43 a_277_47.t0 a_277_47.t1 60.923
R44 D.n0 D.t0 231.014
R45 D.n0 D.t1 158.714
R46 D D.n0 80.266
R47 VGND VGND.t0 107.16
C0 VPWR Y 0.62fF
C1 C Y 0.10fF
C2 C B 0.21fF
C3 B Y 0.23fF
C4 D C 0.11fF
C5 Y VGND 0.13fF
C6 A Y 0.15fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__nand4_2.ext - technology: sky130A

.subckt sky130_fd_sc_hd__nand4_2 B A Y D C VGND VPWR VNB VPB
X0 VPWR.t7 C.t0 Y.t9 VPB.t7 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_471_47.t2 B.t0 a_277_47.t1 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 Y.t8 C.t1 VPWR.t6 VPB.t6 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 VPWR.t0 D.t0 Y.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 VPWR.t4 A.t0 Y.t5 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 a_27_47.t1 D.t1 VGND.t1 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 a_27_47.t3 C.t2 a_277_47.t3 VNB.t7 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 Y.t6 A.t1 VPWR.t5 VPB.t5 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 a_277_47.t0 B.t1 a_471_47.t1 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 VPWR.t2 B.t2 Y.t3 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 Y.t7 A.t2 a_471_47.t3 VNB.t5 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 a_277_47.t2 C.t3 a_27_47.t2 VNB.t6 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 Y.t4 B.t3 VPWR.t3 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13 a_471_47.t0 A.t3 Y.t2 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14 Y.t1 D.t2 VPWR.t1 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 VGND.t0 D.t3 a_27_47.t0 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
R0 C.n0 C.t0 221.719
R1 C.n1 C.t1 221.719
R2 C.n0 C.t2 149.419
R3 C.n1 C.t3 149.419
R4 C.n3 C.n2 76
R5 C.n2 C.n0 37.488
R6 C.n2 C.n1 37.488
R7 C C.n3 28.8
R8 C.n3 C 0.64
R9 Y.n3 Y.n1 138.276
R10 Y.n3 Y.n2 108.604
R11 Y.n5 Y.n4 108.604
R12 Y.n6 Y.n0 106.92
R13 Y Y.n7 106.646
R14 Y.n5 Y.n3 38.981
R15 Y.n6 Y 26.763
R16 Y.n1 Y.t0 26.595
R17 Y.n1 Y.t1 26.595
R18 Y.n2 Y.t9 26.595
R19 Y.n2 Y.t8 26.595
R20 Y.n4 Y.t3 26.595
R21 Y.n4 Y.t4 26.595
R22 Y.n0 Y.t5 26.595
R23 Y.n0 Y.t6 26.595
R24 Y.n7 Y.t2 24.923
R25 Y.n7 Y.t7 24.923
R26 Y Y.n5 13.09
R27 Y.n5 Y 4.266
R28 Y Y.n6 2.536
R29 VPWR.n13 VPWR.n12 174.594
R30 VPWR.n0 VPWR.t4 165.401
R31 VPWR.n8 VPWR.n7 164.214
R32 VPWR.n2 VPWR.n1 164.214
R33 VPWR.n18 VPWR.t1 152.162
R34 VPWR.n1 VPWR.t2 69.935
R35 VPWR.n1 VPWR.t5 62.055
R36 VPWR.n7 VPWR.t3 42.355
R37 VPWR.n7 VPWR.t7 42.355
R38 VPWR.n12 VPWR.t6 26.595
R39 VPWR.n12 VPWR.t0 26.595
R40 VPWR.n4 VPWR.n3 4.65
R41 VPWR.n6 VPWR.n5 4.65
R42 VPWR.n9 VPWR.n8 4.65
R43 VPWR.n11 VPWR.n10 4.65
R44 VPWR.n15 VPWR.n14 4.65
R45 VPWR.n17 VPWR.n16 4.65
R46 VPWR.n19 VPWR.n18 4.65
R47 VPWR.n14 VPWR.n13 3.764
R48 VPWR.n3 VPWR.n2 0.376
R49 VPWR.n4 VPWR.n0 0.235
R50 VPWR.n6 VPWR.n4 0.119
R51 VPWR.n9 VPWR.n6 0.119
R52 VPWR.n11 VPWR.n9 0.119
R53 VPWR.n15 VPWR.n11 0.119
R54 VPWR.n17 VPWR.n15 0.119
R55 VPWR.n19 VPWR.n17 0.119
R56 VPWR VPWR.n19 0.02
R57 VPB.t2 VPB.t5 485.358
R58 VPB.t7 VPB.t3 343.302
R59 VPB.t5 VPB.t4 248.598
R60 VPB.t3 VPB.t2 248.598
R61 VPB.t6 VPB.t7 248.598
R62 VPB.t0 VPB.t6 248.598
R63 VPB.t1 VPB.t0 248.598
R64 VPB VPB.t1 189.408
R65 B.n4 B.t3 237.785
R66 B.n0 B.t2 221.719
R67 B.n1 B.t0 192.263
R68 B.n3 B.t1 149.419
R69 B B.n4 79.2
R70 B.n2 B.n1 76
R71 B.n4 B.n3 55.34
R72 B.n1 B.n0 28.562
R73 B B.n2 28.16
R74 B.n2 B 1.28
R75 a_277_47.n1 a_277_47.n0 251.37
R76 a_277_47.n0 a_277_47.t3 24.923
R77 a_277_47.n0 a_277_47.t2 24.923
R78 a_277_47.n1 a_277_47.t1 24.923
R79 a_277_47.t0 a_277_47.n1 24.923
R80 a_471_47.n0 a_471_47.t1 222.061
R81 a_471_47.n0 a_471_47.t0 135.814
R82 a_471_47.n1 a_471_47.n0 50.6
R83 a_471_47.n1 a_471_47.t3 24.923
R84 a_471_47.t2 a_471_47.n1 24.923
R85 VNB VNB.t1 6053.91
R86 VNB.t7 VNB.t3 4738.46
R87 VNB.t5 VNB.t2 2030.77
R88 VNB.t4 VNB.t5 2030.77
R89 VNB.t3 VNB.t4 2030.77
R90 VNB.t6 VNB.t7 2030.77
R91 VNB.t0 VNB.t6 2030.77
R92 VNB.t1 VNB.t0 2030.77
R93 D.n2 D.t2 234.572
R94 D.n0 D.t0 221.719
R95 D.n2 D.t3 162.272
R96 D.n0 D.t1 149.419
R97 D.n1 D 80.48
R98 D.n3 D.n2 76
R99 D.n1 D.n0 37.488
R100 D.n2 D.n1 24.1
R101 D.n3 D 21.44
R102 D D.n3 8
R103 A.n0 A.t1 221.719
R104 A.n1 A.t0 218.506
R105 A.n0 A.t2 149.419
R106 A.n1 A.t3 146.206
R107 A A.n1 137.967
R108 A.n1 A.n0 74.053
R109 VGND VGND.n0 119.177
R110 VGND.n0 VGND.t1 24.923
R111 VGND.n0 VGND.t0 24.923
R112 a_27_47.n0 a_27_47.t3 225.861
R113 a_27_47.n0 a_27_47.t0 143.678
R114 a_27_47.n1 a_27_47.n0 42.273
R115 a_27_47.n1 a_27_47.t2 24.923
R116 a_27_47.t1 a_27_47.n1 24.923
C0 VPWR Y 1.36fF
C1 VGND VPWR 0.10fF
C2 C Y 0.17fF
C3 VPB VPWR 0.10fF
C4 B Y 0.24fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__nand4_4.ext - technology: sky130A

.subckt sky130_fd_sc_hd__nand4_4 A D C B Y VPWR VGND VNB VPB
X0 a_27_47.t7 C.t0 a_445_47.t3 VNB.t7 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 a_27_47.t6 C.t1 a_445_47.t2 VNB.t6 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 Y.t7 C.t2 VPWR.t7 VPB.t7 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 VPWR.t0 D.t0 Y.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 VPWR.t9 A.t0 Y.t9 VPB.t9 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 Y.t10 A.t1 VPWR.t10 VPB.t10 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 a_445_47.t4 B.t0 a_803_47.t3 VNB.t12 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 Y.t1 D.t1 VPWR.t1 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 a_445_47.t5 B.t1 a_803_47.t2 VNB.t13 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 VPWR.t2 D.t2 Y.t2 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 VPWR.t11 A.t2 Y.t11 VPB.t11 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 a_27_47.t0 D.t3 VGND.t3 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 a_27_47.t1 D.t4 VGND.t2 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 Y.t12 A.t3 a_803_47.t7 VNB.t8 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14 Y.t13 A.t4 a_803_47.t6 VNB.t9 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X15 a_803_47.t1 B.t2 a_445_47.t6 VNB.t14 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X16 VPWR.t6 C.t3 Y.t6 VPB.t6 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17 a_803_47.t0 B.t3 a_445_47.t7 VNB.t15 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X18 VGND.t1 D.t5 a_27_47.t2 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X19 a_445_47.t1 C.t4 a_27_47.t5 VNB.t5 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X20 Y.t5 C.t5 VPWR.t5 VPB.t5 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X21 a_803_47.t5 A.t5 Y.t14 VNB.t10 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X22 VPWR.t13 B.t4 Y.t17 VPB.t13 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X23 Y.t15 A.t6 VPWR.t12 VPB.t12 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X24 a_445_47.t0 C.t6 a_27_47.t4 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X25 a_803_47.t4 A.t7 Y.t16 VNB.t11 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X26 VPWR.t4 C.t7 Y.t4 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X27 Y.t18 B.t5 VPWR.t14 VPB.t14 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X28 VPWR.t15 B.t6 Y.t19 VPB.t15 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X29 Y.t3 D.t6 VPWR.t3 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X30 Y.t8 B.t7 VPWR.t8 VPB.t8 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X31 VGND.t0 D.t7 a_27_47.t3 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
R0 C.n0 C.t3 221.719
R1 C.n2 C.t5 221.719
R2 C.n6 C.t7 221.719
R3 C.n3 C.t2 221.719
R4 C.n0 C.t1 149.419
R5 C.n2 C.t6 149.419
R6 C.n6 C.t0 149.419
R7 C.n3 C.t4 149.419
R8 C.n9 C.n1 76
R9 C.n8 C.n7 76
R10 C.n5 C.n4 76
R11 C.n6 C.n5 38.381
R12 C.n1 C.n0 37.488
R13 C.n2 C.n1 37.488
R14 C.n7 C.n2 37.488
R15 C.n7 C.n6 37.488
R16 C.n5 C.n3 36.596
R17 C.n4 C 23.36
R18 C.n8 C 21.12
R19 C.n9 C 18.56
R20 C C.n9 10.88
R21 C C.n8 8.32
R22 C.n4 C 6.08
R23 a_445_47.n4 a_445_47.n3 135.508
R24 a_445_47.n2 a_445_47.n0 135.508
R25 a_445_47.n2 a_445_47.n1 92.5
R26 a_445_47.n5 a_445_47.n4 92.5
R27 a_445_47.n4 a_445_47.n2 69.632
R28 a_445_47.n3 a_445_47.t3 24.923
R29 a_445_47.n3 a_445_47.t1 24.923
R30 a_445_47.n1 a_445_47.t7 24.923
R31 a_445_47.n1 a_445_47.t5 24.923
R32 a_445_47.n0 a_445_47.t6 24.923
R33 a_445_47.n0 a_445_47.t4 24.923
R34 a_445_47.n5 a_445_47.t2 24.923
R35 a_445_47.t0 a_445_47.n5 24.923
R36 a_27_47.t6 a_27_47.n5 213.093
R37 a_27_47.n2 a_27_47.t3 163.859
R38 a_27_47.n2 a_27_47.n1 94.758
R39 a_27_47.n4 a_27_47.n3 92.5
R40 a_27_47.n5 a_27_47.n0 92.5
R41 a_27_47.n5 a_27_47.n4 57.288
R42 a_27_47.n4 a_27_47.n2 45.266
R43 a_27_47.n0 a_27_47.t4 24.923
R44 a_27_47.n0 a_27_47.t7 24.923
R45 a_27_47.n3 a_27_47.t5 24.923
R46 a_27_47.n3 a_27_47.t1 24.923
R47 a_27_47.n1 a_27_47.t2 24.923
R48 a_27_47.n1 a_27_47.t0 24.923
R49 VNB VNB.t3 6053.91
R50 VNB.t6 VNB.t13 4545.05
R51 VNB.t14 VNB.t8 2320.88
R52 VNB.t9 VNB.t11 2030.77
R53 VNB.t10 VNB.t9 2030.77
R54 VNB.t8 VNB.t10 2030.77
R55 VNB.t12 VNB.t14 2030.77
R56 VNB.t15 VNB.t12 2030.77
R57 VNB.t13 VNB.t15 2030.77
R58 VNB.t4 VNB.t6 2030.77
R59 VNB.t7 VNB.t4 2030.77
R60 VNB.t5 VNB.t7 2030.77
R61 VNB.t1 VNB.t5 2030.77
R62 VNB.t2 VNB.t1 2030.77
R63 VNB.t0 VNB.t2 2030.77
R64 VNB.t3 VNB.t0 2030.77
R65 VPWR.n37 VPWR.n36 174.594
R66 VPWR.n31 VPWR.n30 174.594
R67 VPWR.n25 VPWR.n24 174.594
R68 VPWR.n14 VPWR.n13 174.594
R69 VPWR.n8 VPWR.n7 174.594
R70 VPWR.n2 VPWR.n1 174.594
R71 VPWR.n0 VPWR.t9 155.133
R72 VPWR.n42 VPWR.t3 152.162
R73 VPWR.n19 VPWR.t8 64.531
R74 VPWR.n19 VPWR.t6 64.531
R75 VPWR.n20 VPWR.n19 62.752
R76 VPWR.n7 VPWR.t13 33.49
R77 VPWR.n7 VPWR.t12 31.52
R78 VPWR.n36 VPWR.t1 26.595
R79 VPWR.n36 VPWR.t2 26.595
R80 VPWR.n30 VPWR.t7 26.595
R81 VPWR.n30 VPWR.t0 26.595
R82 VPWR.n24 VPWR.t5 26.595
R83 VPWR.n24 VPWR.t4 26.595
R84 VPWR.n13 VPWR.t14 26.595
R85 VPWR.n13 VPWR.t15 26.595
R86 VPWR.n1 VPWR.t10 26.595
R87 VPWR.n1 VPWR.t11 26.595
R88 VPWR.n26 VPWR.n25 15.811
R89 VPWR.n15 VPWR.n14 11.294
R90 VPWR.n32 VPWR.n31 9.788
R91 VPWR.n9 VPWR.n8 7.905
R92 VPWR.n4 VPWR.n3 4.65
R93 VPWR.n6 VPWR.n5 4.65
R94 VPWR.n10 VPWR.n9 4.65
R95 VPWR.n12 VPWR.n11 4.65
R96 VPWR.n16 VPWR.n15 4.65
R97 VPWR.n18 VPWR.n17 4.65
R98 VPWR.n21 VPWR.n20 4.65
R99 VPWR.n23 VPWR.n22 4.65
R100 VPWR.n27 VPWR.n26 4.65
R101 VPWR.n29 VPWR.n28 4.65
R102 VPWR.n33 VPWR.n32 4.65
R103 VPWR.n35 VPWR.n34 4.65
R104 VPWR.n39 VPWR.n38 4.65
R105 VPWR.n41 VPWR.n40 4.65
R106 VPWR.n43 VPWR.n42 4.65
R107 VPWR.n38 VPWR.n37 3.764
R108 VPWR.n3 VPWR.n2 3.764
R109 VPWR.n4 VPWR.n0 0.746
R110 VPWR.n6 VPWR.n4 0.119
R111 VPWR.n10 VPWR.n6 0.119
R112 VPWR.n12 VPWR.n10 0.119
R113 VPWR.n16 VPWR.n12 0.119
R114 VPWR.n18 VPWR.n16 0.119
R115 VPWR.n21 VPWR.n18 0.119
R116 VPWR.n23 VPWR.n21 0.119
R117 VPWR.n27 VPWR.n23 0.119
R118 VPWR.n29 VPWR.n27 0.119
R119 VPWR.n33 VPWR.n29 0.119
R120 VPWR.n35 VPWR.n33 0.119
R121 VPWR.n39 VPWR.n35 0.119
R122 VPWR.n41 VPWR.n39 0.119
R123 VPWR.n43 VPWR.n41 0.119
R124 VPWR VPWR.n43 0.02
R125 Y.n2 Y.n0 147.876
R126 Y.n5 Y.n3 138.276
R127 Y.n17 Y.n15 135.508
R128 Y.n5 Y.n4 108.604
R129 Y.n7 Y.n6 108.604
R130 Y.n9 Y.n8 108.604
R131 Y.n11 Y.n10 108.604
R132 Y.n13 Y.n12 108.604
R133 Y.n2 Y.n1 104.452
R134 Y.n17 Y.n16 92.5
R135 Y.n11 Y.n9 59.927
R136 Y.n14 Y.n13 36.945
R137 Y.n7 Y.n5 29.672
R138 Y.n9 Y.n7 29.672
R139 Y.n13 Y.n11 29.672
R140 Y.n1 Y.t11 26.595
R141 Y.n1 Y.t15 26.595
R142 Y.n3 Y.t2 26.595
R143 Y.n3 Y.t3 26.595
R144 Y.n4 Y.t0 26.595
R145 Y.n4 Y.t1 26.595
R146 Y.n6 Y.t4 26.595
R147 Y.n6 Y.t7 26.595
R148 Y.n8 Y.t6 26.595
R149 Y.n8 Y.t5 26.595
R150 Y.n10 Y.t19 26.595
R151 Y.n10 Y.t8 26.595
R152 Y.n12 Y.t17 26.595
R153 Y.n12 Y.t18 26.595
R154 Y.n0 Y.t9 26.595
R155 Y.n0 Y.t10 26.595
R156 Y.n15 Y.t16 24.923
R157 Y.n15 Y.t13 24.923
R158 Y.n16 Y.t14 24.923
R159 Y.n16 Y.t12 24.923
R160 Y Y.n14 24.177
R161 Y Y.n17 19.342
R162 Y.n14 Y.n2 5.818
R163 VPB.t6 VPB.t8 556.386
R164 VPB.t13 VPB.t12 284.112
R165 VPB.t10 VPB.t9 248.598
R166 VPB.t11 VPB.t10 248.598
R167 VPB.t12 VPB.t11 248.598
R168 VPB.t14 VPB.t13 248.598
R169 VPB.t15 VPB.t14 248.598
R170 VPB.t8 VPB.t15 248.598
R171 VPB.t5 VPB.t6 248.598
R172 VPB.t4 VPB.t5 248.598
R173 VPB.t7 VPB.t4 248.598
R174 VPB.t0 VPB.t7 248.598
R175 VPB.t1 VPB.t0 248.598
R176 VPB.t2 VPB.t1 248.598
R177 VPB.t3 VPB.t2 248.598
R178 VPB VPB.t3 189.408
R179 D.n3 D.t6 234.39
R180 D.n0 D.t0 221.719
R181 D.n1 D.t1 221.719
R182 D.n7 D.t2 221.719
R183 D.n3 D.t7 162.09
R184 D.n0 D.t4 149.419
R185 D.n1 D.t5 149.419
R186 D.n7 D.t3 149.419
R187 D.n10 D.n2 76
R188 D.n9 D.n8 76
R189 D.n6 D.n5 76
R190 D.n4 D.n3 76
R191 D.n2 D.n0 37.488
R192 D.n2 D.n1 37.488
R193 D.n8 D.n7 37.488
R194 D.n7 D.n6 37.488
R195 D.n10 D.n9 26.88
R196 D.n5 D 24.96
R197 D.n6 D.n3 24.1
R198 D D.n4 21.44
R199 D.n4 D 8
R200 D.n5 D 4.48
R201 D.n9 D 1.92
R202 D D.n10 0.64
R203 A.n0 A.t0 234.572
R204 A.n3 A.t1 221.719
R205 A.n5 A.t2 221.719
R206 A.n4 A.t6 221.719
R207 A.n0 A.t7 162.272
R208 A.n3 A.t4 149.419
R209 A.n5 A.t5 149.419
R210 A.n4 A.t3 149.419
R211 A A.n0 78.88
R212 A.n2 A.n1 76
R213 A.n7 A.n6 76
R214 A.n5 A.n4 74.977
R215 A.n6 A.n3 53.555
R216 A.n2 A.n0 40.166
R217 A.n1 A 28.8
R218 A.n7 A 26.24
R219 A.n3 A.n2 21.422
R220 A.n6 A.n5 21.422
R221 A A.n7 3.2
R222 A.n1 A 0.64
R223 B.n0 B.t4 221.719
R224 B.n1 B.t5 221.719
R225 B.n7 B.t6 221.719
R226 B.n3 B.t7 221.719
R227 B.n0 B.t2 149.419
R228 B.n1 B.t0 149.419
R229 B.n7 B.t3 149.419
R230 B.n3 B.t1 149.419
R231 B.n4 B.n3 118.844
R232 B B.n2 86.88
R233 B.n9 B.n8 76
R234 B.n6 B.n5 76
R235 B.n2 B.n0 37.488
R236 B.n2 B.n1 37.488
R237 B.n8 B.n7 37.488
R238 B.n7 B.n6 37.488
R239 B.n6 B.n3 37.488
R240 B.n4 B 16.64
R241 B B.n9 16
R242 B.n5 B 16
R243 B.n9 B 13.44
R244 B.n5 B 13.44
R245 B B.n4 12.8
R246 a_803_47.n4 a_803_47.t2 213.093
R247 a_803_47.n1 a_803_47.t4 132.789
R248 a_803_47.n1 a_803_47.n0 92.5
R249 a_803_47.n5 a_803_47.n4 92.5
R250 a_803_47.n3 a_803_47.n2 50.599
R251 a_803_47.n4 a_803_47.n3 48.695
R252 a_803_47.n3 a_803_47.n1 48.139
R253 a_803_47.n2 a_803_47.t1 31.384
R254 a_803_47.n2 a_803_47.t7 29.538
R255 a_803_47.n0 a_803_47.t6 24.923
R256 a_803_47.n0 a_803_47.t5 24.923
R257 a_803_47.t3 a_803_47.n5 24.923
R258 a_803_47.n5 a_803_47.t0 24.923
R259 VGND.n2 VGND.n0 111.478
R260 VGND.n2 VGND.n1 111.325
R261 VGND.n0 VGND.t2 24.923
R262 VGND.n0 VGND.t1 24.923
R263 VGND.n1 VGND.t3 24.923
R264 VGND.n1 VGND.t0 24.923
R265 VGND VGND.n2 0.242
C0 Y B 0.47fF
C1 VPB VPWR 0.16fF
C2 Y A 0.36fF
C3 Y D 0.23fF
C4 Y VPWR 2.76fF
C5 Y C 0.42fF
C6 VGND VPWR 0.17fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__nand4b_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__nand4b_1 Y C D A_N B VGND VPWR VNB VPB
X0 Y.t4 B.t0 VPWR.t4 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_232_47.t0 D.t0 VGND.t1 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 VPWR.t1 C.t0 Y.t1 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 VPWR.t3 A_N.t0 a_41_93.t1 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 VPWR.t2 a_41_93.t2 Y.t3 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 a_316_47.t0 C.t1 a_232_47.t1 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 Y.t2 a_41_93.t3 a_423_47.t0 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 a_423_47.t1 B.t1 a_316_47.t1 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 Y.t0 D.t1 VPWR.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 VGND.t0 A_N.t1 a_41_93.t0 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
R0 B.n0 B.t0 241.534
R1 B.n0 B.t1 169.234
R2 B B.n0 78.707
R3  B 16.738
R4 VPWR.n0 VPWR.t2 206.637
R5 VPWR.n2 VPWR.n1 167.037
R6 VPWR.n8 VPWR.n7 126.43
R7 VPWR.n7 VPWR.t3 95.417
R8 VPWR.n1 VPWR.t1 38.415
R9 VPWR.n1 VPWR.t4 37.43
R10 VPWR.n7 VPWR.t0 26.336
R11 VPWR.n9 VPWR.n8 5.652
R12 VPWR.n4 VPWR.n3 4.65
R13 VPWR.n6 VPWR.n5 4.65
R14 VPWR.n3 VPWR.n2 1.505
R15 VPWR.n4 VPWR.n0 0.313
R16 VPWR.n9 VPWR.n6 0.132
R17 VPWR VPWR.n9 0.129
R18 VPWR.n6 VPWR.n4 0.119
R19 Y.n2 Y.n0 154.693
R20 Y.n2 Y.n1 107.441
R21 Y Y.n4 93.809
R22 Y.n3 Y.n2 87.473
R23 Y.n1 Y.t3 50.235
R24 Y.n4 Y.t2 37.846
R25 Y.n0 Y.t1 26.595
R26 Y.n0 Y.t0 26.595
R27 Y.n1 Y.t4 26.595
R28 Y Y.n3 8.581
R29 VPB.t4 VPB.t2 319.626
R30 VPB.t1 VPB.t4 316.666
R31 VPB.t3 VPB.t0 287.071
R32 VPB VPB.t3 269.314
R33 VPB.t0 VPB.t1 248.598
R34 D.n0 D.t1 236.179
R35 D.n0 D.t0 163.879
R36 D D.n0 78.607
R37 VGND VGND.n0 126.322
R38 VGND.n0 VGND.t0 65.714
R39 VGND.n0 VGND.t1 29.538
R40 a_232_47.t0 a_232_47.t1 49.846
R41 VNB VNB.t1 6440.72
R42 VNB.t4 VNB.t0 2610.99
R43 VNB.t1 VNB.t2 2610.99
R44 VNB.t3 VNB.t4 2586.81
R45 VNB.t2 VNB.t3 2030.77
R46 C.n0 C.t0 236.179
R47 C.n0 C.t1 163.879
R48 C C.n0 78.816
R49  C 17.408
R50 A_N.n0 A_N.t0 142.993
R51 A_N.n0 A_N.t1 126.926
R52 A_N A_N.n0 79.684
R53 a_41_93.n1 a_41_93.t1 427.719
R54 a_41_93.n1 a_41_93.n0 270.677
R55 a_41_93.n0 a_41_93.t2 236.179
R56 a_41_93.n0 a_41_93.t3 163.879
R57 a_41_93.t0 a_41_93.n1 132.5
R58 a_316_47.t0 a_316_47.t1 71.076
R59 a_423_47.t0 a_423_47.t1 72
C0 VPWR Y 0.66fF
C1 C B 0.14fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__nand4b_2.ext - technology: sky130A

.subckt sky130_fd_sc_hd__nand4b_2 D C B Y A_N VGND VPWR VNB VPB
X0 Y.t5 a_27_47.t2 a_215_47.t3 VNB.t6 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 a_465_47.t3 B.t0 a_215_47.t0 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 VGND.t1 D.t0 a_655_47.t2 VNB.t7 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 a_215_47.t1 B.t1 a_465_47.t2 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 VPWR.t6 A_N.t0 a_27_47.t0 VPB.t6 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 a_655_47.t3 D.t1 VGND.t0 VNB.t8 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 a_655_47.t0 C.t0 a_465_47.t0 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 VPWR.t5 B.t2 Y.t2 VPB.t5 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 Y.t3 B.t3 VPWR.t4 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 a_465_47.t1 C.t1 a_655_47.t1 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 VPWR.t8 a_27_47.t3 Y.t7 VPB.t8 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 VPWR.t1 C.t2 Y.t1 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 VPWR.t3 D.t2 Y.t8 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13 Y.t9 D.t3 VPWR.t2 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14 a_215_47.t2 a_27_47.t4 Y.t4 VNB.t5 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X15 Y.t6 a_27_47.t5 VPWR.t7 VPB.t7 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16 Y.t0 C.t3 VPWR.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17 VGND.t2 A_N.t1 a_27_47.t1 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
R0 a_27_47.t0 a_27_47.n2 438.894
R1 a_27_47.n0 a_27_47.t3 212.079
R2 a_27_47.n1 a_27_47.t5 212.079
R3 a_27_47.n2 a_27_47.t1 184.026
R4 a_27_47.n2 a_27_47.n1 151.916
R5 a_27_47.n0 a_27_47.t4 139.779
R6 a_27_47.n1 a_27_47.t2 139.779
R7 a_27_47.n1 a_27_47.n0 61.345
R8 a_215_47.n0 a_215_47.t1 212.568
R9 a_215_47.n0 a_215_47.t3 143.23
R10 a_215_47.n1 a_215_47.n0 92.5
R11 a_215_47.t0 a_215_47.n1 24.923
R12 a_215_47.n1 a_215_47.t2 24.923
R13 Y.n3 Y.n1 201.644
R14 Y.n7 Y.n6 108.604
R15 Y.n3 Y.n2 108.604
R16 Y.n5 Y.n4 108.604
R17 Y Y.n0 94.95
R18 Y.n5 Y.n3 57.018
R19 Y.n7 Y.n5 29.672
R20 Y.n6 Y.t7 26.595
R21 Y.n6 Y.t6 26.595
R22 Y.n1 Y.t8 26.595
R23 Y.n1 Y.t9 26.595
R24 Y.n2 Y.t1 26.595
R25 Y.n2 Y.t0 26.595
R26 Y.n4 Y.t2 26.595
R27 Y.n4 Y.t3 26.595
R28 Y.n0 Y.t4 24.923
R29 Y.n0 Y.t5 24.923
R30 Y Y.n7 4.266
R31 VNB VNB.t4 6438.23
R32 VNB.t4 VNB.t6 5321.88
R33 VNB.t3 VNB.t1 4545.05
R34 VNB.t0 VNB.t7 2465.93
R35 VNB.t7 VNB.t8 2030.77
R36 VNB.t1 VNB.t0 2030.77
R37 VNB.t2 VNB.t3 2030.77
R38 VNB.t5 VNB.t2 2030.77
R39 VNB.t6 VNB.t5 2030.77
R40 B.n1 B.t2 212.079
R41 B.n2 B.t3 212.079
R42 B.n1 B.t1 139.779
R43 B.n2 B.t0 139.779
R44 B.n1 B.n0 104.481
R45 B.n4 B.n3 76
R46 B.n3 B.n1 45.278
R47 B.n0 B 25.28
R48 B B.n4 22.4
R49 B.n3 B.n2 16.066
R50 B.n4 B 7.04
R51 B.n0 B 4.16
R52 a_465_47.n1 a_465_47.n0 267.895
R53 a_465_47.n0 a_465_47.t0 24.923
R54 a_465_47.n0 a_465_47.t1 24.923
R55 a_465_47.t2 a_465_47.n1 24.923
R56 a_465_47.n1 a_465_47.t3 24.923
R57 D.n2 D.t3 219.382
R58 D.n1 D.t2 212.079
R59 D.n2 D.t0 139.779
R60 D.n0 D.t1 139.779
R61 D.n0 D 120.507
R62 D.n4 D.n3 76
R63 D.n3 D.n2 35.784
R64 D.n4 D 26.56
R65 D.n3 D.n1 18.257
R66 D.n1 D.n0 7.303
R67 D D.n4 2.88
R68 a_655_47.n0 a_655_47.t1 207.875
R69 a_655_47.n0 a_655_47.t3 136.374
R70 a_655_47.n1 a_655_47.n0 48.532
R71 a_655_47.n1 a_655_47.t2 33.23
R72 a_655_47.t0 a_655_47.n1 33.23
R73 VGND.n1 VGND.t2 149.228
R74 VGND.n1 VGND.n0 123.498
R75 VGND.n0 VGND.t0 24.923
R76 VGND.n0 VGND.t1 24.923
R77 VGND VGND.n1 0.141
R78 A_N.n0 A_N.t0 323.548
R79 A_N.n0 A_N.t1 195.015
R80 A_N.n1 A_N.n0 76
R81 A_N.n1 A_N 15.2
R82 A_N A_N.n1 2.933
R83 VPWR.n21 VPWR.t6 355.821
R84 VPWR.n13 VPWR.n12 174.594
R85 VPWR.n1 VPWR.n0 169.026
R86 VPWR.n2 VPWR.t3 161.926
R87 VPWR.n18 VPWR.t7 131.272
R88 VPWR.n7 VPWR.t0 72.78
R89 VPWR.n8 VPWR.n7 67.176
R90 VPWR.n7 VPWR.t5 57.02
R91 VPWR.n0 VPWR.t2 37.43
R92 VPWR.n0 VPWR.t1 33.49
R93 VPWR.n12 VPWR.t4 26.595
R94 VPWR.n12 VPWR.t8 26.595
R95 VPWR.n20 VPWR.n19 4.65
R96 VPWR.n4 VPWR.n3 4.65
R97 VPWR.n6 VPWR.n5 4.65
R98 VPWR.n9 VPWR.n8 4.65
R99 VPWR.n11 VPWR.n10 4.65
R100 VPWR.n15 VPWR.n14 4.65
R101 VPWR.n17 VPWR.n16 4.65
R102 VPWR.n23 VPWR.n22 4.65
R103 VPWR.n2 VPWR.n1 4.417
R104 VPWR.n14 VPWR.n13 2.258
R105 VPWR.n19 VPWR.n18 0.565
R106 VPWR.n22 VPWR.n21 0.232
R107 VPWR.n4 VPWR.n2 0.229
R108 VPWR.n6 VPWR.n4 0.119
R109 VPWR.n9 VPWR.n6 0.119
R110 VPWR.n11 VPWR.n9 0.119
R111 VPWR.n15 VPWR.n11 0.119
R112 VPWR.n17 VPWR.n15 0.119
R113 VPWR.n20 VPWR.n17 0.119
R114 VPWR.n23 VPWR.n20 0.119
R115 VPWR.n24 VPWR.n23 0.119
R116 VPWR VPWR.n24 0.02
R117 VPB.t6 VPB.t7 556.386
R118 VPB.t5 VPB.t0 526.791
R119 VPB.t1 VPB.t2 301.869
R120 VPB.t2 VPB.t3 248.598
R121 VPB.t0 VPB.t1 248.598
R122 VPB.t4 VPB.t5 248.598
R123 VPB.t8 VPB.t4 248.598
R124 VPB.t7 VPB.t8 248.598
R125 VPB VPB.t6 189.408
R126 C.n3 C.t3 219.382
R127 C.n2 C.t2 212.079
R128 C.n1 C.t0 141.239
R129 C.n3 C.t1 139.779
R130 C.n1 C.n0 76
R131 C.n5 C.n4 76
R132 C.n4 C.n2 48.2
R133 C C.n5 18.56
R134 C.n0 C 16.64
R135 C.n0 C 12.8
R136 C.n5 C 10.88
R137 C.n2 C.n1 5.842
R138 C.n4 C.n3 5.842
C0 VPWR VPB 0.12fF
C1 VPWR Y 1.49fF
C2 B Y 0.31fF
C3 VPWR VGND 0.12fF
C4 C Y 0.29fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__nand4b_4.ext - technology: sky130A

.subckt sky130_fd_sc_hd__nand4b_4 D C B Y A_N VGND VPWR VNB VPB
X0 a_991_47.t7 C.t0 a_633_47.t7 VNB.t14 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 Y.t12 B.t0 VPWR.t10 VPB.t10 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 a_991_47.t2 D.t0 VGND.t3 VNB.t9 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 Y.t0 a_27_47.t2 a_215_47.t7 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 a_991_47.t3 D.t1 VGND.t2 VNB.t10 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 Y.t1 a_27_47.t3 a_215_47.t6 VNB.t5 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 a_633_47.t0 B.t1 a_215_47.t3 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 VPWR.t9 B.t2 Y.t11 VPB.t9 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 Y.t16 C.t1 VPWR.t14 VPB.t14 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 a_633_47.t1 B.t3 a_215_47.t2 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 VGND.t1 D.t2 a_991_47.t0 VNB.t7 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 VPWR.t13 C.t2 Y.t15 VPB.t13 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 VGND.t0 D.t3 a_991_47.t1 VNB.t8 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 a_215_47.t5 a_27_47.t4 Y.t2 VNB.t6 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14 Y.t14 C.t3 VPWR.t12 VPB.t12 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 a_215_47.t1 B.t4 a_633_47.t3 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X16 a_215_47.t0 B.t5 a_633_47.t2 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X17 VPWR.t4 D.t4 Y.t7 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X18 Y.t10 B.t6 VPWR.t8 VPB.t8 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X19 Y.t8 D.t5 VPWR.t5 VPB.t5 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X20 VPWR.t0 a_27_47.t5 Y.t3 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X21 VPWR.t2 D.t6 Y.t5 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X22 Y.t4 a_27_47.t6 VPWR.t1 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X23 a_633_47.t6 C.t4 a_991_47.t6 VNB.t13 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X24 a_633_47.t5 C.t5 a_991_47.t5 VNB.t12 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X25 VPWR.t15 a_27_47.t7 Y.t17 VPB.t15 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X26 Y.t6 D.t7 VPWR.t3 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X27 VPWR.t11 C.t6 Y.t13 VPB.t11 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X28 a_215_47.t4 a_27_47.t8 Y.t18 VNB.t16 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X29 Y.t19 a_27_47.t9 VPWR.t16 VPB.t16 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X30 VPWR.t6 A_N.t0 a_27_47.t0 VPB.t6 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X31 a_991_47.t4 C.t7 a_633_47.t4 VNB.t11 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X32 VPWR.t7 B.t7 Y.t9 VPB.t7 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X33 VGND.t4 A_N.t1 a_27_47.t1 VNB.t15 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
R0 C.n0 C.t6 221.719
R1 C.n1 C.t1 221.719
R2 C.n7 C.t2 221.719
R3 C.n3 C.t3 221.719
R4 C.n0 C.t0 149.419
R5 C.n1 C.t5 149.419
R6 C.n7 C.t7 149.419
R7 C.n3 C.t4 149.419
R8 C.n4 C.n3 130.448
R9 C C.n2 87.2
R10 C.n9 C.n8 76
R11 C.n6 C.n5 76
R12 C.n2 C.n1 38.381
R13 C.n8 C.n7 37.488
R14 C.n7 C.n6 37.488
R15 C.n6 C.n3 37.488
R16 C.n2 C.n0 36.596
R17 C C.n4 16.96
R18 C C.n9 16
R19 C.n5 C 16
R20 C.n9 C 13.44
R21 C.n5 C 13.44
R22 C.n4 C 12.48
R23 a_633_47.n5 a_633_47.n4 132.322
R24 a_633_47.n2 a_633_47.n0 132.322
R25 a_633_47.n2 a_633_47.n1 92.5
R26 a_633_47.n4 a_633_47.n3 92.5
R27 a_633_47.n4 a_633_47.n2 64.474
R28 a_633_47.n3 a_633_47.t2 24.923
R29 a_633_47.n3 a_633_47.t1 24.923
R30 a_633_47.n1 a_633_47.t4 24.923
R31 a_633_47.n1 a_633_47.t6 24.923
R32 a_633_47.n0 a_633_47.t7 24.923
R33 a_633_47.n0 a_633_47.t5 24.923
R34 a_633_47.n5 a_633_47.t3 24.923
R35 a_633_47.t0 a_633_47.n5 24.923
R36 a_991_47.t6 a_991_47.n5 226.776
R37 a_991_47.n1 a_991_47.t3 130.601
R38 a_991_47.n5 a_991_47.n4 92.5
R39 a_991_47.n5 a_991_47.n3 54.999
R40 a_991_47.n1 a_991_47.n0 53.206
R41 a_991_47.n3 a_991_47.n1 51.476
R42 a_991_47.n3 a_991_47.n2 42.273
R43 a_991_47.n4 a_991_47.t5 24.923
R44 a_991_47.n4 a_991_47.t4 24.923
R45 a_991_47.n2 a_991_47.t0 24.923
R46 a_991_47.n2 a_991_47.t7 24.923
R47 a_991_47.n0 a_991_47.t1 24.923
R48 a_991_47.n0 a_991_47.t2 24.923
R49 VNB VNB.t15 6053.91
R50 VNB.t2 VNB.t13 4545.05
R51 VNB.t15 VNB.t4 4545.05
R52 VNB.t8 VNB.t10 2030.77
R53 VNB.t9 VNB.t8 2030.77
R54 VNB.t7 VNB.t9 2030.77
R55 VNB.t14 VNB.t7 2030.77
R56 VNB.t12 VNB.t14 2030.77
R57 VNB.t11 VNB.t12 2030.77
R58 VNB.t13 VNB.t11 2030.77
R59 VNB.t1 VNB.t2 2030.77
R60 VNB.t3 VNB.t1 2030.77
R61 VNB.t0 VNB.t3 2030.77
R62 VNB.t6 VNB.t0 2030.77
R63 VNB.t5 VNB.t6 2030.77
R64 VNB.t16 VNB.t5 2030.77
R65 VNB.t4 VNB.t16 2030.77
R66 B.n1 B.t7 240.693
R67 B.n0 B.t0 221.719
R68 B.n6 B.t2 221.719
R69 B.n7 B.t6 221.719
R70 B.n1 B.t5 168.393
R71 B.n0 B.t3 149.419
R72 B.n6 B.t4 149.419
R73 B.n7 B.t1 149.419
R74 B.n1 B 83.36
R75 B.n3 B.n2 76
R76 B.n5 B.n4 76
R77 B.n9 B.n8 76
R78 B.n8 B.n6 69.622
R79 B.n5 B.n0 58.911
R80 B.n2 B.n1 44.629
R81 B.n3 B 18.24
R82 B.n9 B 17.28
R83 B.n2 B.n0 16.959
R84 B.n6 B.n5 16.066
R85 B.n4 B 16
R86 B.n4 B 13.44
R87 B B.n9 12.16
R88 B B.n3 11.2
R89 B.n8 B.n7 5.355
R90 VPWR.n14 VPWR.n13 174.594
R91 VPWR.n8 VPWR.n7 174.594
R92 VPWR.n2 VPWR.n1 174.594
R93 VPWR.n37 VPWR.n36 174.594
R94 VPWR.n31 VPWR.n30 174.594
R95 VPWR.n25 VPWR.n24 174.594
R96 VPWR.n42 VPWR.t6 172.345
R97 VPWR.n0 VPWR.t4 155.546
R98 VPWR.n42 VPWR.t16 125.929
R99 VPWR.n19 VPWR.t12 70.897
R100 VPWR.n19 VPWR.t7 70.896
R101 VPWR.n20 VPWR.n19 67.448
R102 VPWR.n13 VPWR.t14 26.595
R103 VPWR.n13 VPWR.t13 26.595
R104 VPWR.n7 VPWR.t3 26.595
R105 VPWR.n7 VPWR.t11 26.595
R106 VPWR.n1 VPWR.t5 26.595
R107 VPWR.n1 VPWR.t2 26.595
R108 VPWR.n36 VPWR.t1 26.595
R109 VPWR.n36 VPWR.t15 26.595
R110 VPWR.n30 VPWR.t8 26.595
R111 VPWR.n30 VPWR.t0 26.595
R112 VPWR.n24 VPWR.t10 26.595
R113 VPWR.n24 VPWR.t9 26.595
R114 VPWR.n26 VPWR.n25 14.305
R115 VPWR.n15 VPWR.n14 12.8
R116 VPWR.n43 VPWR.n42 9.089
R117 VPWR.n32 VPWR.n31 8.282
R118 VPWR.n9 VPWR.n8 6.776
R119 VPWR.n4 VPWR.n3 4.65
R120 VPWR.n6 VPWR.n5 4.65
R121 VPWR.n10 VPWR.n9 4.65
R122 VPWR.n12 VPWR.n11 4.65
R123 VPWR.n16 VPWR.n15 4.65
R124 VPWR.n18 VPWR.n17 4.65
R125 VPWR.n21 VPWR.n20 4.65
R126 VPWR.n23 VPWR.n22 4.65
R127 VPWR.n27 VPWR.n26 4.65
R128 VPWR.n29 VPWR.n28 4.65
R129 VPWR.n33 VPWR.n32 4.65
R130 VPWR.n35 VPWR.n34 4.65
R131 VPWR.n39 VPWR.n38 4.65
R132 VPWR.n41 VPWR.n40 4.65
R133 VPWR.n38 VPWR.n37 2.258
R134 VPWR.n44 VPWR.n43 2.132
R135 VPWR.n4 VPWR.n0 0.805
R136 VPWR.n3 VPWR.n2 0.752
R137 VPWR.n44 VPWR.n41 0.191
R138 VPWR VPWR.n44 0.186
R139 VPWR.n6 VPWR.n4 0.119
R140 VPWR.n10 VPWR.n6 0.119
R141 VPWR.n12 VPWR.n10 0.119
R142 VPWR.n16 VPWR.n12 0.119
R143 VPWR.n18 VPWR.n16 0.119
R144 VPWR.n21 VPWR.n18 0.119
R145 VPWR.n23 VPWR.n21 0.119
R146 VPWR.n27 VPWR.n23 0.119
R147 VPWR.n29 VPWR.n27 0.119
R148 VPWR.n33 VPWR.n29 0.119
R149 VPWR.n35 VPWR.n33 0.119
R150 VPWR.n39 VPWR.n35 0.119
R151 VPWR.n41 VPWR.n39 0.119
R152 Y.n16 Y.n15 147.876
R153 Y.n5 Y.n3 138.276
R154 Y.n2 Y.n1 132.322
R155 Y.n5 Y.n4 108.604
R156 Y.n7 Y.n6 108.604
R157 Y.n9 Y.n8 108.604
R158 Y.n11 Y.n10 108.604
R159 Y.n13 Y.n12 108.604
R160 Y.n16 Y.n14 104.452
R161 Y.n2 Y.n0 92.5
R162 Y.n11 Y.n9 59.927
R163 Y.n17 Y.n13 36.654
R164 Y.n7 Y.n5 29.672
R165 Y.n9 Y.n7 29.672
R166 Y.n13 Y.n11 29.672
R167 Y.n14 Y.t3 26.595
R168 Y.n14 Y.t4 26.595
R169 Y.n15 Y.t17 26.595
R170 Y.n15 Y.t19 26.595
R171 Y.n3 Y.t7 26.595
R172 Y.n3 Y.t8 26.595
R173 Y.n4 Y.t5 26.595
R174 Y.n4 Y.t6 26.595
R175 Y.n6 Y.t13 26.595
R176 Y.n6 Y.t16 26.595
R177 Y.n8 Y.t15 26.595
R178 Y.n8 Y.t14 26.595
R179 Y.n10 Y.t9 26.595
R180 Y.n10 Y.t12 26.595
R181 Y.n12 Y.t11 26.595
R182 Y.n12 Y.t10 26.595
R183 Y.n0 Y.t2 24.923
R184 Y.n0 Y.t1 24.923
R185 Y.n1 Y.t18 24.923
R186 Y.n1 Y.t0 24.923
R187 Y Y.n17 16.422
R188 Y.n18 Y 9.66
R189 Y Y.n18 6.762
R190 Y.n17 Y 2.036
R191 Y.n18 Y 1.659
R192 Y Y.n16 0.581
R193 Y Y.n2 0.474
R194 VPB.t7 VPB.t12 556.386
R195 VPB.t6 VPB.t16 556.386
R196 VPB.t5 VPB.t4 248.598
R197 VPB.t2 VPB.t5 248.598
R198 VPB.t3 VPB.t2 248.598
R199 VPB.t11 VPB.t3 248.598
R200 VPB.t14 VPB.t11 248.598
R201 VPB.t13 VPB.t14 248.598
R202 VPB.t12 VPB.t13 248.598
R203 VPB.t10 VPB.t7 248.598
R204 VPB.t9 VPB.t10 248.598
R205 VPB.t8 VPB.t9 248.598
R206 VPB.t0 VPB.t8 248.598
R207 VPB.t1 VPB.t0 248.598
R208 VPB.t15 VPB.t1 248.598
R209 VPB.t16 VPB.t15 248.598
R210 VPB VPB.t6 189.408
R211 D.n0 D.t5 221.719
R212 D.n6 D.t6 221.719
R213 D.n7 D.t7 221.719
R214 D.n1 D.t4 218.506
R215 D.n0 D.t3 149.419
R216 D.n6 D.t0 149.419
R217 D.n7 D.t2 149.419
R218 D.n1 D.t1 146.206
R219 D.n1 D 118.769
R220 D.n3 D.n2 76
R221 D.n5 D.n4 76
R222 D.n9 D.n8 76
R223 D.n2 D.n0 37.488
R224 D.n5 D.n0 37.488
R225 D.n6 D.n5 37.488
R226 D.n8 D.n6 37.488
R227 D.n8 D.n7 37.488
R228 D.n2 D.n1 36.565
R229 D.n4 D 26.24
R230 D.n3 D 25.92
R231 D.n9 D 23.68
R232 D D.n9 5.76
R233 D.n4 D 3.2
R234 D D.n3 0.64
R235 VGND.n32 VGND.t4 195.032
R236 VGND.n1 VGND.n0 119.57
R237 VGND.n3 VGND.n2 114.711
R238 VGND.n0 VGND.t2 24.923
R239 VGND.n0 VGND.t0 24.923
R240 VGND.n2 VGND.t3 24.923
R241 VGND.n2 VGND.t1 24.923
R242 VGND.n5 VGND.n4 4.65
R243 VGND.n7 VGND.n6 4.65
R244 VGND.n9 VGND.n8 4.65
R245 VGND.n11 VGND.n10 4.65
R246 VGND.n13 VGND.n12 4.65
R247 VGND.n15 VGND.n14 4.65
R248 VGND.n17 VGND.n16 4.65
R249 VGND.n19 VGND.n18 4.65
R250 VGND.n21 VGND.n20 4.65
R251 VGND.n23 VGND.n22 4.65
R252 VGND.n25 VGND.n24 4.65
R253 VGND.n27 VGND.n26 4.65
R254 VGND.n29 VGND.n28 4.65
R255 VGND.n31 VGND.n30 4.65
R256 VGND.n33 VGND.n32 4.05
R257 VGND.n4 VGND.n3 3.764
R258 VGND.n5 VGND.n1 0.817
R259 VGND.n33 VGND.n31 0.134
R260 VGND VGND.n33 0.124
R261 VGND.n7 VGND.n5 0.119
R262 VGND.n9 VGND.n7 0.119
R263 VGND.n11 VGND.n9 0.119
R264 VGND.n13 VGND.n11 0.119
R265 VGND.n15 VGND.n13 0.119
R266 VGND.n17 VGND.n15 0.119
R267 VGND.n19 VGND.n17 0.119
R268 VGND.n21 VGND.n19 0.119
R269 VGND.n23 VGND.n21 0.119
R270 VGND.n25 VGND.n23 0.119
R271 VGND.n27 VGND.n25 0.119
R272 VGND.n29 VGND.n27 0.119
R273 VGND.n31 VGND.n29 0.119
R274 a_27_47.n0 a_27_47.t5 221.719
R275 a_27_47.n1 a_27_47.t6 221.719
R276 a_27_47.n3 a_27_47.t7 221.719
R277 a_27_47.n6 a_27_47.t9 221.719
R278 a_27_47.t0 a_27_47.n8 168.033
R279 a_27_47.n0 a_27_47.t4 149.419
R280 a_27_47.n1 a_27_47.t3 149.419
R281 a_27_47.n3 a_27_47.t8 149.419
R282 a_27_47.n6 a_27_47.t2 149.419
R283 a_27_47.n8 a_27_47.t1 122.868
R284 a_27_47.n7 a_27_47.n6 118.844
R285 a_27_47.n5 a_27_47.n2 102.88
R286 a_27_47.n5 a_27_47.n4 76
R287 a_27_47.n1 a_27_47.n0 74.977
R288 a_27_47.n2 a_27_47.n1 37.488
R289 a_27_47.n4 a_27_47.n3 37.488
R290 a_27_47.n8 a_27_47.n7 29.76
R291 a_27_47.n7 a_27_47.n5 28.8
R292 a_215_47.n1 a_215_47.t0 226.776
R293 a_215_47.n3 a_215_47.t7 136.83
R294 a_215_47.n1 a_215_47.n0 92.5
R295 a_215_47.n3 a_215_47.n2 92.5
R296 a_215_47.n5 a_215_47.n4 92.5
R297 a_215_47.n4 a_215_47.n1 51.2
R298 a_215_47.n4 a_215_47.n3 51.2
R299 a_215_47.n2 a_215_47.t6 24.923
R300 a_215_47.n2 a_215_47.t4 24.923
R301 a_215_47.n0 a_215_47.t2 24.923
R302 a_215_47.n0 a_215_47.t1 24.923
R303 a_215_47.t3 a_215_47.n5 24.923
R304 a_215_47.n5 a_215_47.t5 24.923
R305 A_N.n0 A_N.t0 233.987
R306 A_N.n0 A_N.t1 161.687
R307 A_N A_N.n0 84
C0 B Y 0.47fF
C1 VPB VPWR 0.18fF
C2 VPWR Y 2.77fF
C3 C Y 0.46fF
C4 VPWR VGND 0.19fF
C5 D Y 0.22fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__nand4bb_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__nand4bb_1 C D A_N Y B_N VPWR VGND VNB VPB
X0 VGND.t0 B_N.t0 a_27_93.t1 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1 a_496_21.t1 A_N.t0 VPWR.t4 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 Y.t3 a_496_21.t2 a_426_47.t1 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 VPWR.t2 a_496_21.t3 Y.t2 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 a_426_47.t0 a_27_93.t2 a_326_47.t0 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 VPWR.t0 B_N.t1 a_27_93.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 a_496_21.t0 A_N.t1 VGND.t1 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7 Y.t1 a_27_93.t3 VPWR.t3 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 a_218_47.t1 D.t0 VGND.t2 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 a_326_47.t1 C.t0 a_218_47.t0 VNB.t5 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 Y.t4 D.t1 VPWR.t5 VPB.t5 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 VPWR.t1 C.t1 Y.t0 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
R0 B_N.n0 B_N.t1 329.006
R1 B_N.n0 B_N.t0 126.566
R2 B_N.n1 B_N.n0 76
R3  B_N.n1 10.422
R4 B_N.n1 B_N 2.011
R5 a_27_93.t0 a_27_93.n1 454.594
R6 a_27_93.n0 a_27_93.t3 241.534
R7 a_27_93.n1 a_27_93.n0 222.861
R8 a_27_93.n0 a_27_93.t2 169.234
R9 a_27_93.n1 a_27_93.t1 138.6
R10 VGND.n1 VGND.t1 148.74
R11 VGND.n1 VGND.n0 130.131
R12 VGND.n0 VGND.t0 67.142
R13 VGND.n0 VGND.t2 29.538
R14 VGND VGND.n1 0.149
R15 VNB VNB.t0 6078.09
R16 VNB.t1 VNB.t2 5321.88
R17 VNB.t0 VNB.t4 2635.16
R18 VNB.t4 VNB.t5 2610.99
R19 VNB.t3 VNB.t1 2417.58
R20 VNB.t5 VNB.t3 2417.58
R21 A_N.n0 A_N.t0 336.328
R22 A_N.n0 A_N.t1 204.581
R23 A_N.n1 A_N.n0 76
R24 A_N  17.408
R25 A_N.n1 A_N 14.848
R26 A_N A_N.n1 2.56
R27 VPWR.n0 VPWR.t2 561.48
R28 VPWR.n1 VPWR.t4 358.325
R29 VPWR.n13 VPWR.n12 164.235
R30 VPWR.n7 VPWR.n6 164.214
R31 VPWR.n12 VPWR.t0 105.289
R32 VPWR.n12 VPWR.t5 36.314
R33 VPWR.n6 VPWR.t3 34.475
R34 VPWR.n6 VPWR.t1 34.475
R35 VPWR.n1 VPWR.n0 6.097
R36 VPWR.n3 VPWR.n2 4.65
R37 VPWR.n5 VPWR.n4 4.65
R38 VPWR.n9 VPWR.n8 4.65
R39 VPWR.n11 VPWR.n10 4.65
R40 VPWR.n14 VPWR.n13 4.05
R41 VPWR.n8 VPWR.n7 2.258
R42 VPWR.n3 VPWR.n1 2.061
R43 VPWR.n14 VPWR.n11 0.134
R44 VPWR VPWR.n14 0.126
R45 VPWR.n5 VPWR.n3 0.119
R46 VPWR.n9 VPWR.n5 0.119
R47 VPWR.n11 VPWR.n9 0.119
R48 a_496_21.n1 a_496_21.t1 413.18
R49 a_496_21.t0 a_496_21.n1 233.054
R50 a_496_21.n0 a_496_21.t3 212.079
R51 a_496_21.n1 a_496_21.n0 209.989
R52 a_496_21.n0 a_496_21.t2 139.779
R53 VPB.t3 VPB.t4 556.386
R54 VPB.t0 VPB.t5 322.585
R55 VPB.t5 VPB.t1 319.626
R56 VPB.t2 VPB.t3 295.95
R57 VPB.t1 VPB.t2 295.95
R58 VPB VPB.t0 192.367
R59 a_426_47.t0 a_426_47.t1 64.615
R60 Y.n2 Y.n1 172.01
R61 Y.n2 Y.n0 104.452
R62 Y.n4 Y.t3 83.875
R63 Y.n1 Y.t0 38.415
R64 Y.n1 Y.t4 38.415
R65 Y.n0 Y.t2 34.475
R66 Y.n0 Y.t1 34.475
R67 Y.n3 Y 14.336
R68 Y Y.n2 10.917
R69 Y.n4 Y 4.643
R70 Y Y.n4 3.733
R71 Y.n3 Y 3.072
R72 Y Y.n3 1.505
R73 a_326_47.t0 a_326_47.t1 64.615
R74 D.n0 D.t1 236.179
R75 D.n0 D.t0 163.879
R76 D D.n0 79.328
R77 a_218_47.t0 a_218_47.t1 72
R78 C.n0 C.t1 239.503
R79 C.n0 C.t0 167.203
R80 C C.n0 79.2
R81  C 19.781
C0 VPWR Y 0.55fF
C1 Y VGND 0.15fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__nand4bb_2.ext - technology: sky130A

.subckt sky130_fd_sc_hd__nand4bb_2 D C B_N A_N Y VGND VPWR VNB VPB
X0 VPWR.t9 a_193_47.t2 Y.t9 VPB.t9 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 Y.t2 D.t0 VPWR.t4 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 VPWR.t6 C.t0 Y.t4 VPB.t6 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 VGND.t3 D.t1 a_781_47.t1 VNB.t7 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 Y.t8 a_193_47.t3 VPWR.t8 VPB.t8 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 Y.t5 C.t1 VPWR.t7 VPB.t7 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 a_591_47.t3 C.t2 a_781_47.t2 VNB.t9 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 a_781_47.t0 D.t2 VGND.t2 VNB.t6 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 a_781_47.t3 C.t3 a_591_47.t2 VNB.t8 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 VPWR.t0 B_N.t0 a_27_47.t1 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10 a_193_47.t0 A_N.t0 VGND.t1 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11 Y.t6 a_193_47.t4 a_341_47.t3 VNB.t5 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 a_591_47.t1 a_27_47.t2 a_341_47.t1 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 VPWR.t5 D.t3 Y.t3 VPB.t5 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14 a_341_47.t2 a_193_47.t5 Y.t7 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X15 a_341_47.t0 a_27_47.t3 a_591_47.t0 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X16 VPWR.t1 a_27_47.t4 Y.t0 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17 Y.t1 a_27_47.t5 VPWR.t2 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X18 a_193_47.t1 A_N.t1 VPWR.t3 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19 VGND.t0 B_N.t1 a_27_47.t0 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
R0 a_193_47.n2 a_193_47.t1 443.367
R1 a_193_47.n0 a_193_47.t2 221.719
R2 a_193_47.n1 a_193_47.t3 212.079
R3 a_193_47.t0 a_193_47.n2 190.209
R4 a_193_47.n2 a_193_47.n1 155.603
R5 a_193_47.n0 a_193_47.t5 149.419
R6 a_193_47.n1 a_193_47.t4 139.779
R7 a_193_47.n1 a_193_47.n0 72.542
R8 Y.n7 Y.n5 162.969
R9 Y.n2 Y.n0 138.276
R10 Y.n7 Y.n6 124.112
R11 Y.n2 Y.n1 108.604
R12 Y.n8 Y.n4 104.452
R13 Y.n3 Y.n2 51.781
R14 Y.n8 Y.n7 39.272
R15 Y.n4 Y.t0 26.595
R16 Y.n4 Y.t1 26.595
R17 Y.n5 Y.t9 26.595
R18 Y.n5 Y.t8 26.595
R19 Y.n0 Y.t3 26.595
R20 Y.n0 Y.t2 26.595
R21 Y.n1 Y.t4 26.595
R22 Y.n1 Y.t5 26.595
R23 Y.n6 Y.t7 24.923
R24 Y.n6 Y.t6 24.923
R25 Y Y.n8 16
R26 Y.n3 Y 14.268
R27 Y Y.n3 1.745
R28 VPWR.n23 VPWR.n22 312.98
R29 VPWR.n2 VPWR.n1 174.594
R30 VPWR.n13 VPWR.n12 169.933
R31 VPWR.n17 VPWR.t8 159.46
R32 VPWR.n0 VPWR.t5 154.101
R33 VPWR.n7 VPWR.t7 70.897
R34 VPWR.n7 VPWR.t1 70.896
R35 VPWR.n8 VPWR.n7 67.448
R36 VPWR.n22 VPWR.t3 63.321
R37 VPWR.n22 VPWR.t0 63.321
R38 VPWR.n1 VPWR.t4 26.595
R39 VPWR.n1 VPWR.t6 26.595
R40 VPWR.n12 VPWR.t2 26.595
R41 VPWR.n12 VPWR.t9 26.595
R42 VPWR.n18 VPWR.n17 16.564
R43 VPWR.n4 VPWR.n3 4.65
R44 VPWR.n6 VPWR.n5 4.65
R45 VPWR.n11 VPWR.n10 4.65
R46 VPWR.n14 VPWR.n13 4.65
R47 VPWR.n16 VPWR.n15 4.65
R48 VPWR.n19 VPWR.n18 4.65
R49 VPWR.n21 VPWR.n20 4.65
R50 VPWR.n24 VPWR.n23 3.974
R51 VPWR.n3 VPWR.n2 3.011
R52 VPWR.n9 VPWR.n8 2.296
R53 VPWR.n4 VPWR.n0 0.76
R54 VPWR.n9 VPWR.n6 0.178
R55 VPWR.n11 VPWR.n9 0.178
R56 VPWR.n24 VPWR.n21 0.136
R57 VPWR VPWR.n24 0.124
R58 VPWR.n6 VPWR.n4 0.119
R59 VPWR.n14 VPWR.n11 0.119
R60 VPWR.n16 VPWR.n14 0.119
R61 VPWR.n19 VPWR.n16 0.119
R62 VPWR.n21 VPWR.n19 0.119
R63 VPB.t3 VPB.t8 680.685
R64 VPB.t1 VPB.t7 556.386
R65 VPB.t4 VPB.t5 248.598
R66 VPB.t6 VPB.t4 248.598
R67 VPB.t7 VPB.t6 248.598
R68 VPB.t2 VPB.t1 248.598
R69 VPB.t9 VPB.t2 248.598
R70 VPB.t8 VPB.t9 248.598
R71 VPB.t0 VPB.t3 248.598
R72 VPB VPB.t0 192.367
R73 D.n0 D.t3 234.037
R74 D.n1 D.t0 221.719
R75 D.n0 D.t2 161.737
R76 D.n1 D.t1 149.419
R77 D D.n2 83.36
R78 D.n0 D 77.6
R79 D.n2 D.n0 56.233
R80 D.n2 D.n1 5.355
R81 C.n0 C.t0 221.719
R82 C.n1 C.t1 221.719
R83 C.n0 C.t3 149.419
R84 C.n1 C.t2 149.419
R85 C C.n2 85.28
R86 C.n2 C.n0 37.488
R87 C.n2 C.n1 37.488
R88 C C.n3 19.52
R89 C.n3 C 9.92
R90 a_781_47.n1 a_781_47.t2 217.855
R91 a_781_47.t0 a_781_47.n1 141.96
R92 a_781_47.n1 a_781_47.n0 42.273
R93 a_781_47.n0 a_781_47.t1 24.923
R94 a_781_47.n0 a_781_47.t3 24.923
R95 VGND.n2 VGND.n1 121.147
R96 VGND.n2 VGND.n0 115.457
R97 VGND.n0 VGND.t1 38.571
R98 VGND.n0 VGND.t0 38.571
R99 VGND.n1 VGND.t2 24.923
R100 VGND.n1 VGND.t3 24.923
R101 VGND VGND.n2 0.14
R102 VNB.t2 VNB.t5 6680.7
R103 VNB VNB.t0 6470.59
R104 VNB.t1 VNB.t9 4545.05
R105 VNB.t0 VNB.t2 2717.65
R106 VNB.t7 VNB.t6 2030.77
R107 VNB.t8 VNB.t7 2030.77
R108 VNB.t9 VNB.t8 2030.77
R109 VNB.t3 VNB.t1 2030.77
R110 VNB.t4 VNB.t3 2030.77
R111 VNB.t5 VNB.t4 2030.77
R112 a_591_47.n1 a_591_47.n0 254.632
R113 a_591_47.n0 a_591_47.t0 24.923
R114 a_591_47.n0 a_591_47.t1 24.923
R115 a_591_47.t2 a_591_47.n1 24.923
R116 a_591_47.n1 a_591_47.t3 24.923
R117 B_N.n0 B_N.t0 314.906
R118 B_N.n0 B_N.t1 234.573
R119 B_N.n1 B_N.n0 76
R120 B_N.n1 B_N 10.971
R121 B_N B_N.n1 6.791
R122 a_27_47.n3 a_27_47.t1 469.232
R123 a_27_47.t0 a_27_47.n3 230.617
R124 a_27_47.n1 a_27_47.t4 221.719
R125 a_27_47.n0 a_27_47.t5 221.719
R126 a_27_47.n1 a_27_47.t3 149.419
R127 a_27_47.n0 a_27_47.t2 149.419
R128 a_27_47.n2 a_27_47.n1 63.643
R129 a_27_47.n3 a_27_47.n2 16.177
R130 a_27_47.n2 a_27_47.n0 10.112
R131 A_N.n0 A_N.t1 295.948
R132 A_N.n0 A_N.t0 228.468
R133 A_N.n1 A_N.n0 76
R134 A_N.n1 A_N 8.685
R135 A_N A_N.n1 6.857
R136 a_341_47.n0 a_341_47.t0 213.093
R137 a_341_47.n0 a_341_47.t3 203.862
R138 a_341_47.n1 a_341_47.n0 92.5
R139 a_341_47.t1 a_341_47.n1 24.923
R140 a_341_47.n1 a_341_47.t2 24.923
C0 B_N A_N 0.14fF
C1 VPWR Y 1.44fF
C2 VPB VPWR 0.13fF
C3 C Y 0.27fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__nand4bb_4.ext - technology: sky130A

.subckt sky130_fd_sc_hd__nand4bb_4 B_N A_N C Y D VGND VPWR VNB VPB
X0 Y.t15 a_27_47.t2 a_432_47.t7 VNB.t17 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 Y.t19 a_27_47.t3 VPWR.t17 VPB.t17 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 Y.t14 a_27_47.t4 a_432_47.t6 VNB.t16 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 VPWR.t6 C.t0 Y.t5 VPB.t6 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 a_850_47.t3 a_193_47.t2 a_432_47.t0 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 VGND.t3 D.t0 a_1266_47.t3 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 VPWR.t16 a_27_47.t5 Y.t18 VPB.t16 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 Y.t6 C.t1 VPWR.t7 VPB.t7 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 Y.t17 a_27_47.t6 VPWR.t15 VPB.t15 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 VPWR.t1 D.t1 Y.t0 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 a_432_47.t5 a_27_47.t7 Y.t13 VNB.t15 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 a_432_47.t1 a_193_47.t3 a_850_47.t2 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 a_432_47.t4 a_27_47.t8 Y.t12 VNB.t14 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 a_432_47.t2 a_193_47.t4 a_850_47.t1 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14 Y.t9 D.t2 VPWR.t10 VPB.t10 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 VPWR.t2 a_193_47.t5 Y.t1 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16 a_193_47.t0 B_N.t0 VPWR.t13 VPB.t13 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17 Y.t2 a_193_47.t6 VPWR.t3 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X18 VPWR.t11 D.t3 Y.t10 VPB.t11 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X19 a_193_47.t1 B_N.t1 VGND.t4 VNB.t10 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X20 Y.t11 D.t4 VPWR.t12 VPB.t12 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X21 a_850_47.t5 C.t2 a_1266_47.t7 VNB.t5 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X22 a_850_47.t0 a_193_47.t7 a_432_47.t3 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X23 a_850_47.t7 C.t3 a_1266_47.t6 VNB.t6 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X24 VPWR.t8 C.t4 Y.t7 VPB.t8 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X25 VGND.t2 D.t5 a_1266_47.t2 VNB.t9 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X26 Y.t8 C.t5 VPWR.t9 VPB.t9 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X27 VPWR.t4 a_193_47.t8 Y.t3 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X28 a_1266_47.t5 C.t6 a_850_47.t6 VNB.t7 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X29 Y.t4 a_193_47.t9 VPWR.t5 VPB.t5 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X30 a_1266_47.t4 C.t7 a_850_47.t4 VNB.t8 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X31 a_1266_47.t1 D.t6 VGND.t1 VNB.t11 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X32 a_1266_47.t0 D.t7 VGND.t0 VNB.t12 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X33 VPWR.t0 A_N.t0 a_27_47.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X34 VPWR.t14 a_27_47.t9 Y.t16 VPB.t14 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X35 VGND.t5 A_N.t1 a_27_47.t1 VNB.t13 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
R0 a_27_47.t0 a_27_47.n5 610.57
R1 a_27_47.n5 a_27_47.n4 240.318
R2 a_27_47.n1 a_27_47.t9 221.719
R3 a_27_47.n2 a_27_47.t3 221.719
R4 a_27_47.n0 a_27_47.t5 221.719
R5 a_27_47.n4 a_27_47.t6 212.079
R6 a_27_47.n5 a_27_47.t1 208.625
R7 a_27_47.n1 a_27_47.t8 149.419
R8 a_27_47.n2 a_27_47.t4 149.419
R9 a_27_47.n0 a_27_47.t7 149.419
R10 a_27_47.n4 a_27_47.t2 139.779
R11 a_27_47.n2 a_27_47.n1 74.977
R12 a_27_47.n3 a_27_47.n2 64.442
R13 a_27_47.n4 a_27_47.n3 61.75
R14 a_27_47.n3 a_27_47.n0 5.332
R15 a_432_47.n3 a_432_47.t7 241.523
R16 a_432_47.n1 a_432_47.t1 213.093
R17 a_432_47.n1 a_432_47.n0 92.5
R18 a_432_47.n3 a_432_47.n2 92.5
R19 a_432_47.n5 a_432_47.n4 92.5
R20 a_432_47.n4 a_432_47.n1 46.747
R21 a_432_47.n4 a_432_47.n3 46.747
R22 a_432_47.n2 a_432_47.t6 24.923
R23 a_432_47.n2 a_432_47.t5 24.923
R24 a_432_47.n0 a_432_47.t3 24.923
R25 a_432_47.n0 a_432_47.t2 24.923
R26 a_432_47.t0 a_432_47.n5 24.923
R27 a_432_47.n5 a_432_47.t4 24.923
R28 Y.n16 Y.n15 208.262
R29 Y.n5 Y.n3 138.276
R30 Y.n2 Y.n1 135.508
R31 Y.n5 Y.n4 108.604
R32 Y.n7 Y.n6 108.604
R33 Y.n9 Y.n8 108.604
R34 Y.n11 Y.n10 108.604
R35 Y.n13 Y.n12 108.604
R36 Y.n16 Y.n14 104.452
R37 Y.n2 Y.n0 92.5
R38 Y.n11 Y.n9 78.545
R39 Y.n7 Y.n5 29.672
R40 Y.n9 Y.n7 29.672
R41 Y.n13 Y.n11 29.672
R42 Y.n18 Y.n17 29.351
R43 Y.n14 Y.t16 26.595
R44 Y.n14 Y.t19 26.595
R45 Y.n15 Y.t18 26.595
R46 Y.n15 Y.t17 26.595
R47 Y.n3 Y.t0 26.595
R48 Y.n3 Y.t9 26.595
R49 Y.n4 Y.t10 26.595
R50 Y.n4 Y.t11 26.595
R51 Y.n6 Y.t7 26.595
R52 Y.n6 Y.t8 26.595
R53 Y.n8 Y.t5 26.595
R54 Y.n8 Y.t6 26.595
R55 Y.n10 Y.t1 26.595
R56 Y.n10 Y.t2 26.595
R57 Y.n12 Y.t3 26.595
R58 Y.n12 Y.t4 26.595
R59 Y.n0 Y.t12 24.923
R60 Y.n0 Y.t14 24.923
R61 Y.n1 Y.t13 24.923
R62 Y.n1 Y.t15 24.923
R63 Y.n17 Y.n13 21.817
R64 Y Y.n16 16
R65 Y.n18 Y.n2 7.936
R66 Y.n17 Y 1.454
R67 Y Y.n18 0.662
R68 VNB.t10 VNB.t17 7760.44
R69 VNB.t2 VNB.t5 6092.31
R70 VNB VNB.t13 6078.09
R71 VNB.t0 VNB.t12 2030.77
R72 VNB.t11 VNB.t0 2030.77
R73 VNB.t9 VNB.t11 2030.77
R74 VNB.t8 VNB.t9 2030.77
R75 VNB.t6 VNB.t8 2030.77
R76 VNB.t7 VNB.t6 2030.77
R77 VNB.t5 VNB.t7 2030.77
R78 VNB.t4 VNB.t2 2030.77
R79 VNB.t3 VNB.t4 2030.77
R80 VNB.t1 VNB.t3 2030.77
R81 VNB.t14 VNB.t1 2030.77
R82 VNB.t16 VNB.t14 2030.77
R83 VNB.t15 VNB.t16 2030.77
R84 VNB.t17 VNB.t15 2030.77
R85 VNB.t13 VNB.t10 2030.77
R86 VPWR.n56 VPWR.n55 312.98
R87 VPWR.n14 VPWR.n13 174.594
R88 VPWR.n8 VPWR.n7 174.594
R89 VPWR.n2 VPWR.n1 174.594
R90 VPWR.n38 VPWR.n37 174.594
R91 VPWR.n32 VPWR.n31 174.594
R92 VPWR.n44 VPWR.n43 169.933
R93 VPWR.n48 VPWR.t15 159.46
R94 VPWR.n0 VPWR.t1 153.613
R95 VPWR.n26 VPWR.n25 146.25
R96 VPWR.n22 VPWR.n21 146.25
R97 VPWR.n20 VPWR.n19 146.25
R98 VPWR.n25 VPWR.t2 36.445
R99 VPWR.n19 VPWR.t7 32.505
R100 VPWR.n13 VPWR.t9 26.595
R101 VPWR.n13 VPWR.t6 26.595
R102 VPWR.n7 VPWR.t12 26.595
R103 VPWR.n7 VPWR.t8 26.595
R104 VPWR.n1 VPWR.t10 26.595
R105 VPWR.n1 VPWR.t11 26.595
R106 VPWR.n37 VPWR.t5 26.595
R107 VPWR.n37 VPWR.t14 26.595
R108 VPWR.n31 VPWR.t3 26.595
R109 VPWR.n31 VPWR.t4 26.595
R110 VPWR.n43 VPWR.t17 26.595
R111 VPWR.n43 VPWR.t16 26.595
R112 VPWR.n55 VPWR.t13 26.595
R113 VPWR.n55 VPWR.t0 26.595
R114 VPWR.n49 VPWR.n48 16.188
R115 VPWR.n15 VPWR.n14 14.682
R116 VPWR.n9 VPWR.n8 8.658
R117 VPWR.n4 VPWR.n3 4.65
R118 VPWR.n6 VPWR.n5 4.65
R119 VPWR.n10 VPWR.n9 4.65
R120 VPWR.n12 VPWR.n11 4.65
R121 VPWR.n16 VPWR.n15 4.65
R122 VPWR.n18 VPWR.n17 4.65
R123 VPWR.n24 VPWR.n23 4.65
R124 VPWR.n28 VPWR.n27 4.65
R125 VPWR.n30 VPWR.n29 4.65
R126 VPWR.n34 VPWR.n33 4.65
R127 VPWR.n36 VPWR.n35 4.65
R128 VPWR.n40 VPWR.n39 4.65
R129 VPWR.n42 VPWR.n41 4.65
R130 VPWR.n45 VPWR.n44 4.65
R131 VPWR.n47 VPWR.n46 4.65
R132 VPWR.n50 VPWR.n49 4.65
R133 VPWR.n52 VPWR.n51 4.65
R134 VPWR.n54 VPWR.n53 4.65
R135 VPWR.n39 VPWR.n38 4.141
R136 VPWR.n57 VPWR.n56 3.974
R137 VPWR.n23 VPWR.n20 3.232
R138 VPWR.n3 VPWR.n2 2.635
R139 VPWR.n23 VPWR.n22 2.243
R140 VPWR.n33 VPWR.n32 1.882
R141 VPWR.n4 VPWR.n0 0.767
R142 VPWR.n27 VPWR.n26 0.725
R143 VPWR.n57 VPWR.n54 0.136
R144 VPWR VPWR.n57 0.124
R145 VPWR.n6 VPWR.n4 0.119
R146 VPWR.n10 VPWR.n6 0.119
R147 VPWR.n12 VPWR.n10 0.119
R148 VPWR.n16 VPWR.n12 0.119
R149 VPWR.n18 VPWR.n16 0.119
R150 VPWR.n24 VPWR.n18 0.119
R151 VPWR.n28 VPWR.n24 0.119
R152 VPWR.n30 VPWR.n28 0.119
R153 VPWR.n34 VPWR.n30 0.119
R154 VPWR.n36 VPWR.n34 0.119
R155 VPWR.n40 VPWR.n36 0.119
R156 VPWR.n42 VPWR.n40 0.119
R157 VPWR.n45 VPWR.n42 0.119
R158 VPWR.n47 VPWR.n45 0.119
R159 VPWR.n50 VPWR.n47 0.119
R160 VPWR.n52 VPWR.n50 0.119
R161 VPWR.n54 VPWR.n52 0.119
R162 VPB.t13 VPB.t15 950
R163 VPB.t2 VPB.t7 745.794
R164 VPB.t10 VPB.t1 248.598
R165 VPB.t11 VPB.t10 248.598
R166 VPB.t12 VPB.t11 248.598
R167 VPB.t8 VPB.t12 248.598
R168 VPB.t9 VPB.t8 248.598
R169 VPB.t6 VPB.t9 248.598
R170 VPB.t7 VPB.t6 248.598
R171 VPB.t3 VPB.t2 248.598
R172 VPB.t4 VPB.t3 248.598
R173 VPB.t5 VPB.t4 248.598
R174 VPB.t14 VPB.t5 248.598
R175 VPB.t17 VPB.t14 248.598
R176 VPB.t16 VPB.t17 248.598
R177 VPB.t15 VPB.t16 248.598
R178 VPB.t0 VPB.t13 248.598
R179 VPB VPB.t0 192.367
R180 C.n0 C.t4 221.719
R181 C.n2 C.t5 221.719
R182 C.n7 C.t0 221.719
R183 C.n3 C.t1 221.719
R184 C.n0 C.t7 149.419
R185 C.n2 C.t3 149.419
R186 C.n7 C.t6 149.419
R187 C.n3 C.t2 149.419
R188 C.n4 C.n3 118.844
R189 C C.n1 91.68
R190 C.n9 C.n8 76
R191 C.n6 C.n5 76
R192 C.n1 C.n0 37.488
R193 C.n8 C.n2 37.488
R194 C.n8 C.n7 37.488
R195 C.n7 C.n6 37.488
R196 C.n6 C.n3 37.488
R197 C.n4 C 21.44
R198 C.n5 C 20.8
R199 C.n9 C 18.24
R200 C C.n9 11.2
R201 C.n5 C 8.64
R202 C C.n4 8
R203 a_193_47.t0 a_193_47.n13 518.213
R204 a_193_47.n0 a_193_47.t5 221.719
R205 a_193_47.n5 a_193_47.t6 221.719
R206 a_193_47.n7 a_193_47.t8 221.719
R207 a_193_47.n10 a_193_47.t9 221.719
R208 a_193_47.n13 a_193_47.t1 210.425
R209 a_193_47.n0 a_193_47.t3 149.419
R210 a_193_47.n5 a_193_47.t7 149.419
R211 a_193_47.n7 a_193_47.t4 149.419
R212 a_193_47.n10 a_193_47.t2 149.419
R213 a_193_47.n2 a_193_47.n1 103.2
R214 a_193_47.n6 a_193_47.n5 38.381
R215 a_193_47.n1 a_193_47.n0 37.488
R216 a_193_47.n7 a_193_47.n6 36.596
R217 a_193_47.n11 a_193_47.n10 35.703
R218 a_193_47.n13 a_193_47.n12 29.209
R219 a_193_47.n8 a_193_47.n7 24.1
R220 a_193_47.n3 a_193_47.n2 21.76
R221 a_193_47.n9 a_193_47.n8 12.496
R222 a_193_47.n12 a_193_47.n11 9.3
R223 a_193_47.n4 a_193_47.n3 4.48
R224 a_193_47.n11 a_193_47.n9 2.677
R225 a_193_47.n12 a_193_47.n4 0.96
R226 a_850_47.n2 a_850_47.n0 139.247
R227 a_850_47.n5 a_850_47.n4 135.508
R228 a_850_47.n4 a_850_47.n2 124.841
R229 a_850_47.n2 a_850_47.n1 92.5
R230 a_850_47.n4 a_850_47.n3 92.5
R231 a_850_47.n3 a_850_47.t2 24.923
R232 a_850_47.n3 a_850_47.t0 24.923
R233 a_850_47.n1 a_850_47.t6 24.923
R234 a_850_47.n1 a_850_47.t5 24.923
R235 a_850_47.n0 a_850_47.t4 24.923
R236 a_850_47.n0 a_850_47.t7 24.923
R237 a_850_47.n5 a_850_47.t1 24.923
R238 a_850_47.t3 a_850_47.n5 24.923
R239 D.n0 D.t1 233.866
R240 D.n3 D.t2 221.719
R241 D.n4 D.t3 221.719
R242 D.n7 D.t4 221.719
R243 D.n0 D.t7 161.566
R244 D.n3 D.t0 149.419
R245 D.n4 D.t6 149.419
R246 D.n7 D.t5 149.419
R247 D D.n0 78.88
R248 D.n2 D.n1 76
R249 D.n6 D.n5 76
R250 D.n9 D.n8 76
R251 D.n3 D.n2 37.488
R252 D.n5 D.n3 37.488
R253 D.n5 D.n4 37.488
R254 D.n8 D.n7 37.488
R255 D.n2 D.n0 24.1
R256 D.n1 D 24
R257 D.n6 D 21.44
R258 D D.n9 18.88
R259 D.n9 D 10.56
R260 D D.n6 8
R261 D.n1 D 5.44
R262 a_1266_47.n1 a_1266_47.t0 214.053
R263 a_1266_47.n4 a_1266_47.t7 209.99
R264 a_1266_47.n1 a_1266_47.n0 92.5
R265 a_1266_47.n3 a_1266_47.n2 92.5
R266 a_1266_47.n5 a_1266_47.n4 92.5
R267 a_1266_47.n3 a_1266_47.n1 43.008
R268 a_1266_47.n4 a_1266_47.n3 43.008
R269 a_1266_47.n2 a_1266_47.t2 24.923
R270 a_1266_47.n2 a_1266_47.t4 24.923
R271 a_1266_47.n0 a_1266_47.t3 24.923
R272 a_1266_47.n0 a_1266_47.t1 24.923
R273 a_1266_47.t6 a_1266_47.n5 24.923
R274 a_1266_47.n5 a_1266_47.t5 24.923
R275 VGND.n3 VGND.n0 111.524
R276 VGND.n2 VGND.n1 108.015
R277 VGND.n37 VGND.n36 107.239
R278 VGND.n0 VGND.t0 24.923
R279 VGND.n0 VGND.t3 24.923
R280 VGND.n1 VGND.t1 24.923
R281 VGND.n1 VGND.t2 24.923
R282 VGND.n36 VGND.t4 24.923
R283 VGND.n36 VGND.t5 24.923
R284 VGND.n5 VGND.n4 4.65
R285 VGND.n7 VGND.n6 4.65
R286 VGND.n9 VGND.n8 4.65
R287 VGND.n11 VGND.n10 4.65
R288 VGND.n13 VGND.n12 4.65
R289 VGND.n15 VGND.n14 4.65
R290 VGND.n17 VGND.n16 4.65
R291 VGND.n19 VGND.n18 4.65
R292 VGND.n21 VGND.n20 4.65
R293 VGND.n23 VGND.n22 4.65
R294 VGND.n25 VGND.n24 4.65
R295 VGND.n27 VGND.n26 4.65
R296 VGND.n29 VGND.n28 4.65
R297 VGND.n31 VGND.n30 4.65
R298 VGND.n33 VGND.n32 4.65
R299 VGND.n35 VGND.n34 4.65
R300 VGND.n38 VGND.n37 3.932
R301 VGND.n3 VGND.n2 3.659
R302 VGND.n5 VGND.n3 0.256
R303 VGND.n38 VGND.n35 0.137
R304 VGND VGND.n38 0.123
R305 VGND.n7 VGND.n5 0.119
R306 VGND.n9 VGND.n7 0.119
R307 VGND.n11 VGND.n9 0.119
R308 VGND.n13 VGND.n11 0.119
R309 VGND.n15 VGND.n13 0.119
R310 VGND.n17 VGND.n15 0.119
R311 VGND.n19 VGND.n17 0.119
R312 VGND.n21 VGND.n19 0.119
R313 VGND.n23 VGND.n21 0.119
R314 VGND.n25 VGND.n23 0.119
R315 VGND.n27 VGND.n25 0.119
R316 VGND.n29 VGND.n27 0.119
R317 VGND.n31 VGND.n29 0.119
R318 VGND.n33 VGND.n31 0.119
R319 VGND.n35 VGND.n33 0.119
R320 B_N.n0 B_N.t0 241.534
R321 B_N.n0 B_N.t1 169.234
R322 B_N.n1 B_N.n0 76
R323  B_N.n1 9.475
R324 B_N.n1 B_N 1.828
R325 A_N.n0 A_N.t0 230.154
R326 A_N.n0 A_N.t1 157.854
R327 A_N.n1 A_N.n0 76
R328  A_N.n1 15.86
R329 A_N.n1 A_N 3.06
C0 VPWR Y 2.76fF
C1 VPB VPWR 0.21fF
C2 VPWR VGND 0.18fF
C3 C Y 0.48fF
C4 A_N B_N 0.13fF
C5 D Y 0.22fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__nor2_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__nor2_1 B Y A VGND VPWR VNB VPB
X0 VPWR.t0 A.t0 a_109_297.t1 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 VGND.t0 A.t1 Y.t1 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 a_109_297.t0 B.t0 Y.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 Y.t2 B.t1 VGND.t1 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
R0 A.n0 A.t0 231.833
R1 A.n0 A.t1 157.068
R2 A A.n0 78.011
R3 a_109_297.t0 a_109_297.t1 41.37
R4 VPWR VPWR.t0 149.986
R5 VPB.t0 VPB.t1 213.084
R6 VPB VPB.t0 189.408
R7 Y.n1 Y.n0 133.958
R8 Y.n1 Y.t0 121.129
R9 Y.n0 Y.t1 24.923
R10 Y.n0 Y.t2 24.923
R11 Y Y.n1 7.467
R12 VGND.n0 VGND.t1 114.511
R13 VGND.n0 VGND.t0 111.917
R14 VGND VGND.n0 0.124
R15 VNB VNB.t1 6053.91
R16 VNB.t1 VNB.t0 2030.77
R17 B.n0 B.t0 230.361
R18 B.n0 B.t1 158.061
R19 B B.n0 82.4
C0 Y VPWR 0.14fF
C1 B Y 0.10fF
C2 Y VGND 0.27fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__nor2_2.ext - technology: sky130A

.subckt sky130_fd_sc_hd__nor2_2 B Y A VGND VPWR VNB VPB
X0 Y.t3 B.t0 a_27_297.t1 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 Y.t1 B.t1 VGND.t1 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 a_27_297.t0 A.t0 VPWR.t1 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 VGND.t3 A.t1 Y.t5 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 Y.t4 A.t2 VGND.t2 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 VGND.t0 B.t2 Y.t0 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 VPWR.t0 A.t3 a_27_297.t3 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 a_27_297.t2 B.t3 Y.t2 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
R0 B.n0 B.t3 212.079
R1 B.n1 B.t0 212.079
R2 B.n0 B.t2 139.779
R3 B.n1 B.t1 139.779
R4  B.n2 76.64
R5 B.n2 B.n0 30.672
R6 B.n2 B.n1 30.672
R7  B 29.44
R8 a_27_297.n0 a_27_297.t2 257.327
R9 a_27_297.n0 a_27_297.t3 202.763
R10 a_27_297.n1 a_27_297.n0 87.815
R11 a_27_297.n1 a_27_297.t1 26.595
R12 a_27_297.t0 a_27_297.n1 26.595
R13 Y.n4 Y.n3 146.345
R14 Y.n2 Y.n0 88.89
R15 Y.n4 Y.n2 77.859
R16 Y.n2 Y.n1 52.624
R17 Y.n3 Y.t2 26.595
R18 Y.n3 Y.t3 26.595
R19 Y.n1 Y.t0 24.923
R20 Y.n1 Y.t1 24.923
R21 Y.n0 Y.t5 24.923
R22 Y.n0 Y.t4 24.923
R23 Y Y.n4 3.203
R24 VPB.t2 VPB.t1 248.598
R25 VPB.t0 VPB.t2 248.598
R26 VPB.t3 VPB.t0 248.598
R27 VPB VPB.t3 201.246
R28 VGND.n2 VGND.t0 192.178
R29 VGND.n1 VGND.n0 115.464
R30 VGND.n5 VGND.t2 104.607
R31 VGND.n0 VGND.t1 24.923
R32 VGND.n0 VGND.t3 24.923
R33 VGND.n2 VGND.n1 6.315
R34 VGND.n6 VGND.n5 4.65
R35 VGND.n4 VGND.n3 4.65
R36 VGND.n4 VGND.n2 0.213
R37 VGND.n6 VGND.n4 0.119
R38 VGND VGND.n6 0.02
R39 VNB VNB.t2 6150.61
R40 VNB.t1 VNB.t0 2030.77
R41 VNB.t3 VNB.t1 2030.77
R42 VNB.t2 VNB.t3 2030.77
R43 A.n0 A.t0 212.079
R44 A.n1 A.t3 212.079
R45 A.n0 A.t1 139.779
R46 A.n1 A.t2 139.779
R47  A.n2 78.24
R48 A.n2 A.n0 38.706
R49  A 29.44
R50 A.n2 A.n1 22.639
R51 VPWR VPWR.n0 167.774
R52 VPWR.n0 VPWR.t1 26.595
R53 VPWR.n0 VPWR.t0 26.595
C0 Y VGND 0.48fF
C1 B Y 0.25fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__nor2_4.ext - technology: sky130A

.subckt sky130_fd_sc_hd__nor2_4 Y A B VGND VPWR VNB VPB
X0 VPWR.t3 A.t0 a_27_297.t3 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 Y.t3 A.t1 VGND.t3 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 a_27_297.t2 A.t2 VPWR.t2 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 VGND.t2 A.t3 Y.t2 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 a_27_297.t4 B.t0 Y.t4 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 Y.t1 A.t4 VGND.t1 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 VGND.t0 A.t5 Y.t0 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 VGND.t4 B.t1 Y.t5 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 VGND.t5 B.t2 Y.t6 VNB.t5 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 Y.t7 B.t3 a_27_297.t5 VPB.t5 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 VPWR.t1 A.t6 a_27_297.t1 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 Y.t8 B.t4 VGND.t6 VNB.t6 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 Y.t9 B.t5 VGND.t7 VNB.t7 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 a_27_297.t6 B.t6 Y.t10 VPB.t6 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14 Y.t11 B.t7 a_27_297.t7 VPB.t7 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 a_27_297.t0 A.t7 VPWR.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
R0 A.n0 A.t7 212.079
R1 A.n2 A.t0 212.079
R2 A.n7 A.t2 212.079
R3 A.n8 A.t6 212.079
R4 A.n0 A.t5 139.779
R5 A.n2 A.t1 139.779
R6 A.n7 A.t3 139.779
R7 A.n8 A.t4 139.779
R8 A.n6 A.n5 76
R9 A.n10 A.n9 76
R10 A.n6 A.n3 49.66
R11 A.n9 A.n7 45.278
R12 A.n2 A.n1 42.357
R13  A.n10 28.8
R14 A.n5 A.n4 21.76
R15 A.n5 A 21.12
R16 A.n1 A.n0 18.987
R17 A.n9 A.n8 16.066
R18 A.n3 A.n2 7.303
R19 A.n7 A.n6 4.381
R20 A.n10 A 0.64
R21 a_27_297.n1 a_27_297.t4 215.054
R22 a_27_297.n3 a_27_297.t1 181.277
R23 a_27_297.n1 a_27_297.n0 150.25
R24 a_27_297.n3 a_27_297.n2 109.334
R25 a_27_297.n5 a_27_297.n4 91.601
R26 a_27_297.n4 a_27_297.n3 57.04
R27 a_27_297.n4 a_27_297.n1 53.037
R28 a_27_297.n2 a_27_297.t3 26.595
R29 a_27_297.n2 a_27_297.t2 26.595
R30 a_27_297.n0 a_27_297.t5 26.595
R31 a_27_297.n0 a_27_297.t6 26.595
R32 a_27_297.n5 a_27_297.t7 26.595
R33 a_27_297.t0 a_27_297.n5 26.595
R34 VPWR.n2 VPWR.n0 173.48
R35 VPWR.n2 VPWR.n1 167.523
R36 VPWR.n0 VPWR.t0 26.595
R37 VPWR.n0 VPWR.t3 26.595
R38 VPWR.n1 VPWR.t2 26.595
R39 VPWR.n1 VPWR.t1 26.595
R40 VPWR VPWR.n2 0.244
R41 VPB.t5 VPB.t4 248.598
R42 VPB.t6 VPB.t5 248.598
R43 VPB.t7 VPB.t6 248.598
R44 VPB.t0 VPB.t7 248.598
R45 VPB.t3 VPB.t0 248.598
R46 VPB.t2 VPB.t3 248.598
R47 VPB.t1 VPB.t2 248.598
R48 VPB VPB.t1 201.246
R49 VGND.n2 VGND.t5 193.83
R50 VGND.n1 VGND.n0 115.464
R51 VGND.n6 VGND.n5 115.464
R52 VGND.n12 VGND.n11 115.464
R53 VGND.n17 VGND.t1 104.607
R54 VGND.n0 VGND.t7 24.923
R55 VGND.n0 VGND.t4 24.923
R56 VGND.n5 VGND.t6 24.923
R57 VGND.n5 VGND.t0 24.923
R58 VGND.n11 VGND.t3 24.923
R59 VGND.n11 VGND.t2 24.923
R60 VGND.n2 VGND.n1 18.218
R61 VGND.n7 VGND.n6 8.282
R62 VGND.n18 VGND.n17 4.65
R63 VGND.n4 VGND.n3 4.65
R64 VGND.n8 VGND.n7 4.65
R65 VGND.n10 VGND.n9 4.65
R66 VGND.n14 VGND.n13 4.65
R67 VGND.n16 VGND.n15 4.65
R68 VGND.n13 VGND.n12 2.258
R69 VGND.n4 VGND.n2 0.356
R70 VGND.n8 VGND.n4 0.119
R71 VGND.n10 VGND.n8 0.119
R72 VGND.n14 VGND.n10 0.119
R73 VGND.n16 VGND.n14 0.119
R74 VGND.n18 VGND.n16 0.119
R75 VGND VGND.n18 0.02
R76 Y.n2 Y.n1 186.028
R77 Y.n2 Y.n0 150.188
R78 Y.n5 Y.n3 88.89
R79 Y.n5 Y.n4 52.624
R80 Y.n7 Y.n6 52.624
R81 Y.n9 Y.n8 52.624
R82 Y Y.n9 39.36
R83 Y.n7 Y.n5 36.266
R84 Y.n9 Y.n7 36.266
R85 Y.n0 Y.t4 26.595
R86 Y.n0 Y.t7 26.595
R87 Y.n1 Y.t10 26.595
R88 Y.n1 Y.t11 26.595
R89 Y.n3 Y.t2 24.923
R90 Y.n3 Y.t1 24.923
R91 Y.n4 Y.t0 24.923
R92 Y.n4 Y.t3 24.923
R93 Y.n6 Y.t5 24.923
R94 Y.n6 Y.t8 24.923
R95 Y.n8 Y.t6 24.923
R96 Y.n8 Y.t9 24.923
R97 Y Y.n2 23.36
R98 VNB VNB.t1 6150.61
R99 VNB.t7 VNB.t5 2030.77
R100 VNB.t4 VNB.t7 2030.77
R101 VNB.t6 VNB.t4 2030.77
R102 VNB.t0 VNB.t6 2030.77
R103 VNB.t3 VNB.t0 2030.77
R104 VNB.t2 VNB.t3 2030.77
R105 VNB.t1 VNB.t2 2030.77
R106 B.n0 B.t0 212.079
R107 B.n2 B.t3 212.079
R108 B.n7 B.t6 212.079
R109 B.n5 B.t7 212.079
R110 B.n0 B.t2 139.779
R111 B.n2 B.t5 139.779
R112 B.n7 B.t1 139.779
R113 B.n5 B.t4 139.779
R114 B.n9 B.n6 97.76
R115 B.n4 B.n1 97.76
R116 B.n4 B.n3 76
R117 B.n9 B.n8 76
R118 B.n6 B.n5 18.257
R119 B B.n9 17.6
R120 B.n1 B.n0 16.796
R121 B.n8 B.n7 6.572
R122 B.n3 B.n2 5.112
R123 B B.n4 4.16
C0 A Y 0.24fF
C1 Y VGND 0.96fF
C2 B Y 0.50fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__nor2_8.ext - technology: sky130A

.subckt sky130_fd_sc_hd__nor2_8 Y A B VGND VPWR VNB VPB
X0 VPWR.t7 A.t0 a_27_297.t7 VPB.t7 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 Y.t15 B.t0 a_27_297.t8 VPB.t8 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 a_27_297.t9 B.t1 Y.t14 VPB.t9 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 Y.t7 A.t1 VGND.t7 VNB.t7 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 a_27_297.t6 A.t2 VPWR.t6 VPB.t6 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 Y.t23 B.t2 VGND.t15 VNB.t15 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 a_27_297.t10 B.t3 Y.t13 VPB.t10 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 Y.t12 B.t4 a_27_297.t11 VPB.t11 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 VGND.t6 A.t3 Y.t6 VNB.t6 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 a_27_297.t5 A.t4 VPWR.t5 VPB.t5 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 Y.t5 A.t5 VGND.t5 VNB.t5 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 VGND.t4 A.t6 Y.t4 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 VGND.t3 A.t7 Y.t3 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 VGND.t2 A.t8 Y.t2 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14 VPWR.t4 A.t9 a_27_297.t4 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 a_27_297.t12 B.t5 Y.t11 VPB.t12 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16 Y.t10 B.t6 a_27_297.t13 VPB.t13 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17 VPWR.t3 A.t10 a_27_297.t3 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X18 Y.t1 A.t11 VGND.t1 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X19 a_27_297.t14 B.t7 Y.t9 VPB.t14 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X20 Y.t0 A.t12 VGND.t0 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X21 Y.t22 B.t8 VGND.t14 VNB.t14 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X22 Y.t21 B.t9 VGND.t13 VNB.t13 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X23 Y.t20 B.t10 VGND.t12 VNB.t12 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X24 Y.t8 B.t11 a_27_297.t15 VPB.t15 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X25 a_27_297.t2 A.t13 VPWR.t2 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X26 VGND.t11 B.t12 Y.t19 VNB.t11 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X27 VPWR.t1 A.t14 a_27_297.t1 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X28 VGND.t10 B.t13 Y.t18 VNB.t10 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X29 VGND.t9 B.t14 Y.t17 VNB.t9 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X30 VGND.t8 B.t15 Y.t16 VNB.t8 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X31 a_27_297.t0 A.t15 VPWR.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
R0 A.n0 A.t4 212.079
R1 A.n2 A.t9 212.079
R2 A.n5 A.t13 212.079
R3 A.n10 A.t14 212.079
R4 A.n13 A.t15 212.079
R5 A.n16 A.t0 212.079
R6 A.n19 A.t2 212.079
R7 A.n22 A.t10 212.079
R8 A.n0 A.t8 139.779
R9 A.n2 A.t12 139.779
R10 A.n5 A.t7 139.779
R11 A.n10 A.t11 139.779
R12 A.n13 A.t6 139.779
R13 A.n16 A.t1 139.779
R14 A.n19 A.t3 139.779
R15 A.n22 A.t5 139.779
R16 A.n4 A.n1 97.76
R17 A A.n23 76.32
R18 A.n4 A.n3 76
R19 A.n7 A.n6 76
R20 A.n9 A.n8 76
R21 A.n12 A.n11 76
R22 A.n15 A.n14 76
R23 A.n18 A.n17 76
R24 A.n21 A.n20 76
R25 A.n11 A.n10 30.672
R26 A.n7 A.n4 21.76
R27 A.n9 A.n7 21.76
R28 A.n12 A.n9 21.76
R29 A.n15 A.n12 21.76
R30 A.n18 A.n15 21.76
R31 A.n21 A.n18 21.76
R32 A A.n21 21.44
R33 A.n14 A.n13 18.987
R34 A.n1 A.n0 16.066
R35 A.n23 A.n22 16.066
R36 A.n6 A.n5 7.303
R37 A.n17 A.n16 7.303
R38 A.n3 A.n2 4.381
R39 A.n20 A.n19 4.381
R40 a_27_297.n4 a_27_297.t12 225.591
R41 a_27_297.n1 a_27_297.t3 169.847
R42 a_27_297.n4 a_27_297.n3 154.573
R43 a_27_297.n6 a_27_297.n5 154.573
R44 a_27_297.n8 a_27_297.n7 154.573
R45 a_27_297.n13 a_27_297.n12 109.737
R46 a_27_297.n11 a_27_297.n10 109.736
R47 a_27_297.n1 a_27_297.n0 109.736
R48 a_27_297.n9 a_27_297.n2 90.234
R49 a_27_297.n9 a_27_297.n8 64.95
R50 a_27_297.n11 a_27_297.n9 55.464
R51 a_27_297.n6 a_27_297.n4 44.423
R52 a_27_297.n8 a_27_297.n6 44.423
R53 a_27_297.n12 a_27_297.n1 35.961
R54 a_27_297.n12 a_27_297.n11 35.961
R55 a_27_297.n2 a_27_297.t11 26.595
R56 a_27_297.n2 a_27_297.t5 26.595
R57 a_27_297.n3 a_27_297.t13 26.595
R58 a_27_297.n3 a_27_297.t14 26.595
R59 a_27_297.n5 a_27_297.t15 26.595
R60 a_27_297.n5 a_27_297.t9 26.595
R61 a_27_297.n7 a_27_297.t8 26.595
R62 a_27_297.n7 a_27_297.t10 26.595
R63 a_27_297.n10 a_27_297.t4 26.595
R64 a_27_297.n10 a_27_297.t2 26.595
R65 a_27_297.n0 a_27_297.t7 26.595
R66 a_27_297.n0 a_27_297.t6 26.595
R67 a_27_297.n13 a_27_297.t1 26.595
R68 a_27_297.t0 a_27_297.n13 26.595
R69 VPWR.n3 VPWR.n2 175.843
R70 VPWR.n12 VPWR.n11 169.933
R71 VPWR.n1 VPWR.n0 169.933
R72 VPWR.n7 VPWR.n6 169.933
R73 VPWR.n2 VPWR.t5 26.595
R74 VPWR.n2 VPWR.t4 26.595
R75 VPWR.n0 VPWR.t2 26.595
R76 VPWR.n0 VPWR.t1 26.595
R77 VPWR.n6 VPWR.t0 26.595
R78 VPWR.n6 VPWR.t7 26.595
R79 VPWR.n11 VPWR.t6 26.595
R80 VPWR.n11 VPWR.t3 26.595
R81 VPWR.n3 VPWR.n1 5.772
R82 VPWR.n5 VPWR.n4 4.65
R83 VPWR.n8 VPWR.n7 4.65
R84 VPWR.n10 VPWR.n9 4.65
R85 VPWR.n13 VPWR.n12 4.024
R86 VPWR.n5 VPWR.n3 0.379
R87 VPWR.n13 VPWR.n10 0.135
R88 VPWR VPWR.n13 0.125
R89 VPWR.n8 VPWR.n5 0.119
R90 VPWR.n10 VPWR.n8 0.119
R91 VPB.t13 VPB.t12 248.598
R92 VPB.t14 VPB.t13 248.598
R93 VPB.t15 VPB.t14 248.598
R94 VPB.t9 VPB.t15 248.598
R95 VPB.t8 VPB.t9 248.598
R96 VPB.t10 VPB.t8 248.598
R97 VPB.t11 VPB.t10 248.598
R98 VPB.t5 VPB.t11 248.598
R99 VPB.t4 VPB.t5 248.598
R100 VPB.t2 VPB.t4 248.598
R101 VPB.t1 VPB.t2 248.598
R102 VPB.t0 VPB.t1 248.598
R103 VPB.t7 VPB.t0 248.598
R104 VPB.t6 VPB.t7 248.598
R105 VPB.t3 VPB.t6 248.598
R106 VPB VPB.t3 204.205
R107 B.n0 B.t5 212.079
R108 B.n1 B.t6 212.079
R109 B.n2 B.t7 212.079
R110 B.n6 B.t11 212.079
R111 B.n9 B.t1 212.079
R112 B.n17 B.t0 212.079
R113 B.n14 B.t3 212.079
R114 B.n12 B.t4 212.079
R115 B.n0 B.t15 139.779
R116 B.n1 B.t2 139.779
R117 B.n2 B.t14 139.779
R118 B.n6 B.t9 139.779
R119 B.n9 B.t12 139.779
R120 B.n17 B.t10 139.779
R121 B.n14 B.t13 139.779
R122 B.n12 B.t8 139.779
R123 B.n16 B.n13 97.76
R124 B.n5 B.n4 76
R125 B.n8 B.n7 76
R126 B.n11 B.n10 76
R127 B.n19 B.n18 76
R128 B.n16 B.n15 76
R129 B.n1 B.n0 61.345
R130 B.n5 B.n3 55.015
R131 B.n7 B.n6 28.481
R132 B.n3 B.n2 26.386
R133 B.n3 B.n1 23.92
R134 B.n8 B.n5 21.76
R135 B.n11 B.n8 21.76
R136 B.n19 B.n16 21.76
R137 B.n13 B.n12 18.257
R138 B.n10 B.n9 16.796
R139 B B.n11 16
R140 B.n15 B.n14 6.572
R141 B B.n19 5.76
R142 B.n18 B.n17 5.112
R143 Y.n2 Y.n0 199.508
R144 Y.n2 Y.n1 155.085
R145 Y.n4 Y.n3 155.085
R146 Y.n6 Y.n5 155.085
R147 Y.n10 Y.n8 88.89
R148 Y.n10 Y.n9 52.624
R149 Y.n12 Y.n11 52.624
R150 Y.n14 Y.n13 52.624
R151 Y.n16 Y.n15 52.624
R152 Y.n18 Y.n17 52.624
R153 Y.n20 Y.n19 52.624
R154 Y.n21 Y.n7 49.285
R155 Y.n21 Y.n20 47.999
R156 Y.n4 Y.n2 44.423
R157 Y.n6 Y.n4 44.423
R158 Y Y.n21 41.388
R159 Y.n12 Y.n10 36.266
R160 Y.n14 Y.n12 36.266
R161 Y.n16 Y.n14 36.266
R162 Y.n18 Y.n16 36.266
R163 Y.n20 Y.n18 36.266
R164 Y.n0 Y.t13 26.595
R165 Y.n0 Y.t12 26.595
R166 Y.n1 Y.t14 26.595
R167 Y.n1 Y.t15 26.595
R168 Y.n3 Y.t9 26.595
R169 Y.n3 Y.t8 26.595
R170 Y.n5 Y.t11 26.595
R171 Y.n5 Y.t10 26.595
R172 Y.n7 Y.t16 24.923
R173 Y.n7 Y.t23 24.923
R174 Y.n8 Y.t6 24.923
R175 Y.n8 Y.t5 24.923
R176 Y.n9 Y.t4 24.923
R177 Y.n9 Y.t7 24.923
R178 Y.n11 Y.t3 24.923
R179 Y.n11 Y.t1 24.923
R180 Y.n13 Y.t2 24.923
R181 Y.n13 Y.t0 24.923
R182 Y.n15 Y.t18 24.923
R183 Y.n15 Y.t22 24.923
R184 Y.n17 Y.t19 24.923
R185 Y.n17 Y.t20 24.923
R186 Y.n19 Y.t17 24.923
R187 Y.n19 Y.t21 24.923
R188 Y Y.n6 2.301
R189 VGND.n2 VGND.t8 192.131
R190 VGND.n1 VGND.n0 115.464
R191 VGND.n6 VGND.n5 115.464
R192 VGND.n12 VGND.n11 115.464
R193 VGND.n18 VGND.n17 115.464
R194 VGND.n22 VGND.n21 115.464
R195 VGND.n28 VGND.n27 115.464
R196 VGND.n34 VGND.n33 115.464
R197 VGND.n39 VGND.t5 104.607
R198 VGND.n0 VGND.t15 24.923
R199 VGND.n0 VGND.t9 24.923
R200 VGND.n5 VGND.t13 24.923
R201 VGND.n5 VGND.t11 24.923
R202 VGND.n11 VGND.t12 24.923
R203 VGND.n11 VGND.t10 24.923
R204 VGND.n17 VGND.t14 24.923
R205 VGND.n17 VGND.t2 24.923
R206 VGND.n21 VGND.t0 24.923
R207 VGND.n21 VGND.t3 24.923
R208 VGND.n27 VGND.t1 24.923
R209 VGND.n27 VGND.t4 24.923
R210 VGND.n33 VGND.t7 24.923
R211 VGND.n33 VGND.t6 24.923
R212 VGND.n19 VGND.n18 14.305
R213 VGND.n23 VGND.n22 14.305
R214 VGND.n13 VGND.n12 8.282
R215 VGND.n29 VGND.n28 8.282
R216 VGND.n2 VGND.n1 7.817
R217 VGND.n40 VGND.n39 4.65
R218 VGND.n4 VGND.n3 4.65
R219 VGND.n8 VGND.n7 4.65
R220 VGND.n10 VGND.n9 4.65
R221 VGND.n14 VGND.n13 4.65
R222 VGND.n16 VGND.n15 4.65
R223 VGND.n20 VGND.n19 4.65
R224 VGND.n24 VGND.n23 4.65
R225 VGND.n26 VGND.n25 4.65
R226 VGND.n30 VGND.n29 4.65
R227 VGND.n32 VGND.n31 4.65
R228 VGND.n36 VGND.n35 4.65
R229 VGND.n38 VGND.n37 4.65
R230 VGND.n7 VGND.n6 2.258
R231 VGND.n35 VGND.n34 2.258
R232 VGND.n4 VGND.n2 0.218
R233 VGND.n8 VGND.n4 0.119
R234 VGND.n10 VGND.n8 0.119
R235 VGND.n14 VGND.n10 0.119
R236 VGND.n16 VGND.n14 0.119
R237 VGND.n20 VGND.n16 0.119
R238 VGND.n24 VGND.n20 0.119
R239 VGND.n26 VGND.n24 0.119
R240 VGND.n30 VGND.n26 0.119
R241 VGND.n32 VGND.n30 0.119
R242 VGND.n36 VGND.n32 0.119
R243 VGND.n38 VGND.n36 0.119
R244 VGND.n40 VGND.n38 0.119
R245 VGND VGND.n40 0.022
R246 VNB VNB.t5 6174.79
R247 VNB.t15 VNB.t8 2030.77
R248 VNB.t9 VNB.t15 2030.77
R249 VNB.t13 VNB.t9 2030.77
R250 VNB.t11 VNB.t13 2030.77
R251 VNB.t12 VNB.t11 2030.77
R252 VNB.t10 VNB.t12 2030.77
R253 VNB.t14 VNB.t10 2030.77
R254 VNB.t2 VNB.t14 2030.77
R255 VNB.t0 VNB.t2 2030.77
R256 VNB.t3 VNB.t0 2030.77
R257 VNB.t1 VNB.t3 2030.77
R258 VNB.t4 VNB.t1 2030.77
R259 VNB.t7 VNB.t4 2030.77
R260 VNB.t6 VNB.t7 2030.77
R261 VNB.t5 VNB.t6 2030.77
C0 VPWR VGND 0.16fF
C1 A Y 0.55fF
C2 VPB B 0.11fF
C3 Y VGND 1.82fF
C4 B Y 1.01fF
C5 VPB VPWR 0.14fF
C6 VPB A 0.10fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__nor2b_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__nor2b_1 B_N Y A VGND VPWR VNB VPB
X0 Y.t0 a_74_47.t2 a_265_297.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 VPWR.t1 B_N.t0 a_74_47.t1 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 a_265_297.t1 A.t0 VPWR.t0 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 Y.t2 A.t1 VGND.t1 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 VGND.t2 B_N.t1 a_74_47.t0 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 VGND.t0 a_74_47.t3 Y.t1 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
R0 a_74_47.n1 a_74_47.t1 362.467
R1 a_74_47.n0 a_74_47.t2 236.179
R2 a_74_47.t0 a_74_47.n1 210.277
R3 a_74_47.n1 a_74_47.n0 170.4
R4 a_74_47.n0 a_74_47.t3 163.879
R5 a_265_297.t0 a_265_297.t1 41.37
R6 Y.n1 Y.t0 173.353
R7 Y.n1 Y.n0 166.613
R8 Y.n0 Y.t1 24.923
R9 Y.n0 Y.t2 24.923
R10 Y Y.n1 1.434
R11 VPB VPB.t2 334.423
R12 VPB.t2 VPB.t1 319.626
R13 VPB.t1 VPB.t0 213.084
R14 B_N.n0 B_N.t1 176.733
R15 B_N B_N.n0 147.046
R16 B_N.n0 B_N.t0 119.623
R17  B_N 19.342
R18 VPWR VPWR.n0 169.473
R19 VPWR.n0 VPWR.t1 121.952
R20 VPWR.n0 VPWR.t0 25.61
R21 A.n0 A.t0 236.179
R22 A.n0 A.t1 163.879
R23 A A.n0 80.676
R24 VGND.n1 VGND.t0 187.535
R25 VGND.n1 VGND.n0 81.179
R26 VGND.n0 VGND.t2 57.772
R27 VGND.n0 VGND.t1 24.789
R28 VGND VGND.n1 0.295
R29 VNB VNB.t2 8355.68
R30 VNB.t2 VNB.t1 2303.7
R31 VNB.t1 VNB.t0 2030.77
C0 Y VGND 0.33fF
C1 VPWR Y 0.14fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__nor2b_2.ext - technology: sky130A

.subckt sky130_fd_sc_hd__nor2b_2 B_N A Y VGND VPWR VNB VPB
X0 Y.t1 a_251_21.t2 a_27_297.t1 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 Y.t3 a_251_21.t3 VGND.t1 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 a_27_297.t2 A.t0 VPWR.t1 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 VGND.t2 A.t1 Y.t4 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 Y.t5 A.t2 VGND.t3 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 VGND.t0 a_251_21.t4 Y.t2 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 VPWR.t0 A.t3 a_27_297.t3 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 VPWR.t2 B_N.t0 a_251_21.t0 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 VGND.t4 B_N.t1 a_251_21.t1 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9 a_27_297.t0 a_251_21.t5 Y.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
R0 a_251_21.t0 a_251_21.n2 433.143
R1 a_251_21.n1 a_251_21.t5 212.079
R2 a_251_21.n0 a_251_21.t2 212.079
R3 a_251_21.n2 a_251_21.t1 156.452
R4 a_251_21.n1 a_251_21.t4 139.779
R5 a_251_21.n0 a_251_21.t3 139.779
R6 a_251_21.n2 a_251_21.n1 131.533
R7 a_251_21.n1 a_251_21.n0 61.345
R8 a_27_297.t0 a_27_297.n1 200.245
R9 a_27_297.n1 a_27_297.t3 190.115
R10 a_27_297.n1 a_27_297.n0 90.234
R11 a_27_297.n0 a_27_297.t1 26.595
R12 a_27_297.n0 a_27_297.t2 26.595
R13 Y.n2 Y.n1 190.893
R14 Y Y.n4 93.857
R15 Y.n2 Y.n0 90.831
R16 Y.n1 Y.t0 26.595
R17 Y.n1 Y.t1 26.595
R18 Y.n4 Y.t2 24.923
R19 Y.n4 Y.t3 24.923
R20 Y.n0 Y.t4 24.923
R21 Y.n0 Y.t5 24.923
R22 Y Y.n3 11.83
R23 Y.n3 Y.n2 3.103
R24 VPB.t0 VPB.t4 556.386
R25 VPB.t1 VPB.t0 248.598
R26 VPB.t2 VPB.t1 248.598
R27 VPB.t3 VPB.t2 248.598
R28 VPB VPB.t3 201.246
R29 VGND.n1 VGND.t4 169.161
R30 VGND.n5 VGND.n4 115.464
R31 VGND.n0 VGND.t0 114.4
R32 VGND.n10 VGND.t3 104.882
R33 VGND.n4 VGND.t1 24.923
R34 VGND.n4 VGND.t2 24.923
R35 VGND.n1 VGND.n0 12.335
R36 VGND.n11 VGND.n10 4.65
R37 VGND.n3 VGND.n2 4.65
R38 VGND.n7 VGND.n6 4.65
R39 VGND.n9 VGND.n8 4.65
R40 VGND.n6 VGND.n5 2.258
R41 VGND.n3 VGND.n1 0.218
R42 VGND.n7 VGND.n3 0.119
R43 VGND.n9 VGND.n7 0.119
R44 VGND.n11 VGND.n9 0.119
R45 VGND VGND.n11 0.02
R46 VNB VNB.t3 6150.61
R47 VNB.t0 VNB.t4 5321.88
R48 VNB.t1 VNB.t0 2030.77
R49 VNB.t2 VNB.t1 2030.77
R50 VNB.t3 VNB.t2 2030.77
R51 A.n0 A.t0 212.079
R52 A.n1 A.t3 212.079
R53 A.n0 A.t1 139.779
R54 A.n1 A.t2 139.779
R55 A A.n2 77.6
R56 A.n2 A.n0 38.706
R57 A.n2 A.n1 22.639
R58 VPWR.n1 VPWR.t2 381.226
R59 VPWR.n1 VPWR.n0 173.445
R60 VPWR.n0 VPWR.t1 26.595
R61 VPWR.n0 VPWR.t0 26.595
R62 VPWR VPWR.n1 0.142
R63 B_N.n0 B_N.t0 333.171
R64 B_N.n0 B_N.t1 130.731
R65 B_N.n1 B_N.n0 84.838
R66  B_N.n1 16.372
R67 B_N.n1 B_N 3.869
C0 Y VGND 0.49fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__nor2b_4.ext - technology: sky130A

.subckt sky130_fd_sc_hd__nor2b_4 B_N Y A VGND VPWR VNB VPB
X0 VPWR.t3 A.t0 a_27_297.t7 VPB.t7 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 Y.t11 A.t1 VGND.t6 VNB.t7 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 a_27_297.t6 A.t2 VPWR.t2 VPB.t6 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 VGND.t5 A.t3 Y.t10 VNB.t6 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 a_27_297.t0 a_419_21.t2 Y.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 Y.t9 A.t4 VGND.t4 VNB.t5 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 VGND.t7 A.t5 Y.t8 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 VGND.t0 a_419_21.t3 Y.t1 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 VGND.t1 a_419_21.t4 Y.t2 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 Y.t3 a_419_21.t5 a_27_297.t1 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 VPWR.t1 A.t6 a_27_297.t5 VPB.t5 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 Y.t4 a_419_21.t6 VGND.t2 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 VGND.t8 B_N.t0 a_419_21.t0 VNB.t8 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 Y.t5 a_419_21.t7 VGND.t3 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14 VPWR.t4 B_N.t1 a_419_21.t1 VPB.t8 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 a_27_297.t2 a_419_21.t8 Y.t6 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16 Y.t7 a_419_21.t9 a_27_297.t3 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17 a_27_297.t4 A.t7 VPWR.t0 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
R0 A.n0 A.t7 212.079
R1 A.n2 A.t0 212.079
R2 A.n5 A.t2 212.079
R3 A.n8 A.t6 212.079
R4 A.n0 A.t5 139.779
R5 A.n2 A.t1 139.779
R6 A.n5 A.t3 139.779
R7 A.n8 A.t4 139.779
R8 A.n4 A.n1 97.76
R9 A A.n9 76.64
R10 A.n4 A.n3 76
R11 A.n7 A.n6 76
R12 A.n7 A.n4 21.76
R13 A A.n7 21.12
R14 A.n1 A.n0 18.987
R15 A.n9 A.n8 16.066
R16 A.n3 A.n2 7.303
R17 A.n6 A.n5 4.381
R18 a_27_297.n2 a_27_297.t5 181.085
R19 a_27_297.t0 a_27_297.n5 169.982
R20 a_27_297.n5 a_27_297.n4 150.25
R21 a_27_297.n2 a_27_297.n1 109.334
R22 a_27_297.n3 a_27_297.n0 91.601
R23 a_27_297.n3 a_27_297.n2 57.039
R24 a_27_297.n5 a_27_297.n3 53.035
R25 a_27_297.n0 a_27_297.t3 26.595
R26 a_27_297.n0 a_27_297.t4 26.595
R27 a_27_297.n1 a_27_297.t7 26.595
R28 a_27_297.n1 a_27_297.t6 26.595
R29 a_27_297.n4 a_27_297.t1 26.595
R30 a_27_297.n4 a_27_297.t2 26.595
R31 VPWR.n1 VPWR.n0 169.933
R32 VPWR.n6 VPWR.n5 164.214
R33 VPWR.n2 VPWR.t4 146.245
R34 VPWR.n0 VPWR.t0 26.595
R35 VPWR.n0 VPWR.t3 26.595
R36 VPWR.n5 VPWR.t2 26.595
R37 VPWR.n5 VPWR.t1 26.595
R38 VPWR.n4 VPWR.n3 4.65
R39 VPWR.n2 VPWR.n1 4.126
R40 VPWR.n7 VPWR.n6 3.966
R41 VPWR.n7 VPWR.n4 0.137
R42 VPWR.n4 VPWR.n2 0.134
R43 VPWR VPWR.n7 0.122
R44 VPB.t0 VPB.t8 574.143
R45 VPB.t1 VPB.t0 248.598
R46 VPB.t2 VPB.t1 248.598
R47 VPB.t3 VPB.t2 248.598
R48 VPB.t4 VPB.t3 248.598
R49 VPB.t7 VPB.t4 248.598
R50 VPB.t6 VPB.t7 248.598
R51 VPB.t5 VPB.t6 248.598
R52 VPB VPB.t5 201.246
R53 VGND.n5 VGND.n4 115.464
R54 VGND.n11 VGND.n10 115.464
R55 VGND.n17 VGND.n16 115.464
R56 VGND.n1 VGND.t8 109.099
R57 VGND.n0 VGND.t1 106.289
R58 VGND.n22 VGND.t4 104.219
R59 VGND.n4 VGND.t3 24.923
R60 VGND.n4 VGND.t0 24.923
R61 VGND.n10 VGND.t2 24.923
R62 VGND.n10 VGND.t7 24.923
R63 VGND.n16 VGND.t6 24.923
R64 VGND.n16 VGND.t5 24.923
R65 VGND.n6 VGND.n5 14.305
R66 VGND.n1 VGND.n0 8.896
R67 VGND.n12 VGND.n11 8.282
R68 VGND.n23 VGND.n22 4.65
R69 VGND.n3 VGND.n2 4.65
R70 VGND.n7 VGND.n6 4.65
R71 VGND.n9 VGND.n8 4.65
R72 VGND.n13 VGND.n12 4.65
R73 VGND.n15 VGND.n14 4.65
R74 VGND.n19 VGND.n18 4.65
R75 VGND.n21 VGND.n20 4.65
R76 VGND.n18 VGND.n17 2.258
R77 VGND.n3 VGND.n1 0.266
R78 VGND.n7 VGND.n3 0.119
R79 VGND.n9 VGND.n7 0.119
R80 VGND.n13 VGND.n9 0.119
R81 VGND.n15 VGND.n13 0.119
R82 VGND.n19 VGND.n15 0.119
R83 VGND.n21 VGND.n19 0.119
R84 VGND.n23 VGND.n21 0.119
R85 VGND VGND.n23 0.02
R86 Y Y.n0 163.414
R87 Y.n9 Y.n1 152.296
R88 Y.n8 Y.n2 94.934
R89 Y.n6 Y.n4 88.89
R90 Y.n6 Y.n5 52.624
R91 Y.n7 Y.n3 49.285
R92 Y.n7 Y.n6 47.999
R93 Y.n9 Y.n8 26.763
R94 Y.n0 Y.t0 26.595
R95 Y.n0 Y.t3 26.595
R96 Y.n1 Y.t6 26.595
R97 Y.n1 Y.t7 26.595
R98 Y.n3 Y.t1 24.923
R99 Y.n3 Y.t4 24.923
R100 Y.n4 Y.t10 24.923
R101 Y.n4 Y.t9 24.923
R102 Y.n5 Y.t8 24.923
R103 Y.n5 Y.t11 24.923
R104 Y.n2 Y.t2 24.923
R105 Y.n2 Y.t5 24.923
R106 Y Y.n9 12.16
R107 Y.n8 Y.n7 5.688
R108 VNB VNB.t5 6150.61
R109 VNB.t1 VNB.t8 4690.11
R110 VNB.t3 VNB.t1 2030.77
R111 VNB.t0 VNB.t3 2030.77
R112 VNB.t2 VNB.t0 2030.77
R113 VNB.t4 VNB.t2 2030.77
R114 VNB.t7 VNB.t4 2030.77
R115 VNB.t6 VNB.t7 2030.77
R116 VNB.t5 VNB.t6 2030.77
R117 a_419_21.n6 a_419_21.t2 212.079
R118 a_419_21.n0 a_419_21.t5 212.079
R119 a_419_21.n2 a_419_21.t8 212.079
R120 a_419_21.n1 a_419_21.t9 212.079
R121 a_419_21.t1 a_419_21.n8 154.904
R122 a_419_21.n6 a_419_21.t4 139.779
R123 a_419_21.n0 a_419_21.t7 139.779
R124 a_419_21.n2 a_419_21.t3 139.779
R125 a_419_21.n1 a_419_21.t6 139.779
R126 a_419_21.n8 a_419_21.t0 107.578
R127 a_419_21.n4 a_419_21.n3 97.76
R128 a_419_21.n7 a_419_21.n6 73.418
R129 a_419_21.n2 a_419_21.n1 61.345
R130 a_419_21.n3 a_419_21.n2 54.042
R131 a_419_21.n7 a_419_21.n4 29.163
R132 a_419_21.n6 a_419_21.n5 18.987
R133 a_419_21.n8 a_419_21.n7 15.119
R134 a_419_21.n3 a_419_21.n0 7.303
R135 B_N.n0 B_N.t1 229.752
R136 B_N.n0 B_N.t0 157.452
R137 B_N B_N.n0 83.314
C0 VPWR VGND 0.11fF
C1 B_N VPWR 0.11fF
C2 A Y 0.25fF
C3 Y VGND 0.92fF
C4 VPB VPWR 0.11fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__nor3_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__nor3_1 C Y A B VGND VPWR VNB VPB
X0 VPWR.t0 A.t0 a_193_297.t0 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_193_297.t1 B.t0 a_109_297.t1 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 Y.t3 B.t1 VGND.t2 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 VGND.t1 A.t1 Y.t2 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 a_109_297.t0 C.t0 Y.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 VGND.t0 C.t1 Y.t1 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
R0 A.n0 A.t0 229
R1 A.n0 A.t1 156.7
R2 A.n1 A.n0 76
R3  A 16.118
R4 A.n1  13.511
R5  A.n1 2.607
R6 a_193_297.t0 a_193_297.t1 53.19
R7 VPWR VPWR.t0 195.938
R8 VPB.t2 VPB.t1 248.598
R9 VPB.t0 VPB.t2 248.598
R10 VPB VPB.t0 189.408
R11 B.n0 B.t0 241.534
R12 B.n0 B.t1 169.234
R13 B B.n0 89.517
R14  B 18.519
R15 a_109_297.t0 a_109_297.t1 53.19
R16 VGND.n1 VGND.t1 189.916
R17 VGND.n1 VGND.n0 110.927
R18 VGND.n0 VGND.t2 24.923
R19 VGND.n0 VGND.t0 24.923
R20 VGND VGND.n1 0.253
R21 Y.n1 Y.t1 183.807
R22 Y.n2 Y.n1 169.378
R23 Y.n2 Y.t0 125.745
R24 Y.n1 Y.n0 100.405
R25 Y.n0 Y.t2 24.923
R26 Y.n0 Y.t3 24.923
R27 Y Y.n2 2.785
R28 VNB VNB.t0 6053.91
R29 VNB.t2 VNB.t1 2030.77
R30 VNB.t0 VNB.t2 2030.77
R31 C.n0 C.t0 231.014
R32 C.n0 C.t1 158.714
R33 C C.n0 80.266
C0 C B 0.11fF
C1 Y VGND 0.20fF
C2 A Y 0.14fF
C3 C Y 0.12fF
C4 Y VPWR 0.23fF
C5 B Y 0.32fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__nor3_2.ext - technology: sky130A

.subckt sky130_fd_sc_hd__nor3_2 C Y A B VGND VPWR VNB VPB
X0 Y.t7 C.t0 a_281_297.t3 VPB.t5 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_281_297.t0 B.t0 a_27_297.t2 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 Y.t0 B.t1 VGND.t2 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 a_27_297.t3 A.t0 VPWR.t1 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 VGND.t3 A.t1 Y.t3 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 Y.t2 A.t2 VGND.t0 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 VGND.t1 B.t2 Y.t1 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 VGND.t5 C.t1 Y.t5 VNB.t5 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 Y.t4 C.t2 VGND.t4 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 VPWR.t0 A.t3 a_27_297.t0 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 a_281_297.t2 C.t3 Y.t6 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 a_27_297.t1 B.t3 a_281_297.t1 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
R0 C.n0 C.t3 212.079
R1 C.n1 C.t0 212.079
R2 C.n0 C.t1 139.779
R3 C.n1 C.t2 139.779
R4 C.n3 C.n2 85.752
R5 C.n2 C.n0 48.2
R6 C.n2 C.n1 13.145
R7  C.n3 12.8
R8 C.n3 C 3.622
R9 a_281_297.n0 a_281_297.t2 225.591
R10 a_281_297.n1 a_281_297.n0 211.042
R11 a_281_297.n0 a_281_297.t3 182.726
R12 a_281_297.n1 a_281_297.t1 26.595
R13 a_281_297.t0 a_281_297.n1 26.595
R14 Y Y.n0 165.55
R15 Y.n3 Y.n1 88.89
R16 Y.n5 Y.n3 74.666
R17 Y.n3 Y.n2 52.624
R18 Y.n5 Y.n4 52.624
R19 Y.n0 Y.t6 26.595
R20 Y.n0 Y.t7 26.595
R21 Y.n1 Y.t3 24.923
R22 Y.n1 Y.t2 24.923
R23 Y.n2 Y.t1 24.923
R24 Y.n2 Y.t0 24.923
R25 Y.n4 Y.t5 24.923
R26 Y.n4 Y.t4 24.923
R27 Y Y.n5 21.085
R28 VPB.t1 VPB.t5 568.224
R29 VPB.t5 VPB.t4 248.598
R30 VPB.t0 VPB.t1 248.598
R31 VPB.t3 VPB.t0 248.598
R32 VPB.t2 VPB.t3 248.598
R33 VPB VPB.t2 201.246
R34 B.n0 B.t3 212.079
R35 B.n1 B.t0 212.079
R36 B.n0 B.t2 139.779
R37 B.n1 B.t1 139.779
R38 B B.n2 76.304
R39 B.n2 B.n0 32.863
R40 B.n2 B.n1 28.481
R41  B 28.038
R42 a_27_297.n0 a_27_297.t1 225.591
R43 a_27_297.n0 a_27_297.t0 181.527
R44 a_27_297.n1 a_27_297.n0 110.761
R45 a_27_297.t2 a_27_297.n1 26.595
R46 a_27_297.n1 a_27_297.t3 26.595
R47 VGND.n1 VGND.t5 192.17
R48 VGND.n2 VGND.t1 170.961
R49 VGND.n0 VGND.t4 170.961
R50 VGND.n8 VGND.n7 115.464
R51 VGND.n13 VGND.t0 105.27
R52 VGND.n7 VGND.t2 24.923
R53 VGND.n7 VGND.t3 24.923
R54 VGND.n14 VGND.n13 4.65
R55 VGND.n4 VGND.n3 4.65
R56 VGND.n6 VGND.n5 4.65
R57 VGND.n10 VGND.n9 4.65
R58 VGND.n12 VGND.n11 4.65
R59 VGND.n1 VGND.n0 4.613
R60 VGND.n9 VGND.n8 2.258
R61 VGND.n3 VGND.n2 2.2
R62 VGND.n4 VGND.n1 0.22
R63 VGND.n6 VGND.n4 0.119
R64 VGND.n10 VGND.n6 0.119
R65 VGND.n12 VGND.n10 0.119
R66 VGND.n14 VGND.n12 0.119
R67 VGND VGND.n14 0.02
R68 VNB VNB.t0 6150.61
R69 VNB.t1 VNB.t4 4641.76
R70 VNB.t4 VNB.t5 2030.77
R71 VNB.t2 VNB.t1 2030.77
R72 VNB.t3 VNB.t2 2030.77
R73 VNB.t0 VNB.t3 2030.77
R74 A.n0 A.t0 212.079
R75 A.n1 A.t3 212.079
R76 A.n0 A.t1 139.779
R77 A.n1 A.t2 139.779
R78 A A.n2 78.133
R79 A.n2 A.n0 38.706
R80  A 28.038
R81 A.n2 A.n1 22.639
R82 VPWR VPWR.n0 175.636
R83 VPWR.n0 VPWR.t1 26.595
R84 VPWR.n0 VPWR.t0 26.595
C0 B Y 0.23fF
C1 Y VGND 0.87fF
C2 C Y 0.21fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__nor3_4.ext - technology: sky130A

.subckt sky130_fd_sc_hd__nor3_4 A C B Y VGND VPWR VNB VPB
X0 VPWR.t3 A.t0 a_27_297.t7 VPB.t11 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_449_297.t7 C.t0 Y.t15 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 a_27_297.t0 B.t0 a_449_297.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 Y.t7 A.t1 VGND.t7 VNB.t7 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 a_27_297.t6 A.t2 VPWR.t2 VPB.t10 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 Y.t14 C.t1 a_449_297.t6 VPB.t5 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 a_449_297.t5 C.t2 Y.t13 VPB.t6 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 VGND.t6 A.t3 Y.t6 VNB.t6 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 Y.t12 C.t3 a_449_297.t4 VPB.t7 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 Y.t5 A.t4 VGND.t5 VNB.t5 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 VGND.t4 A.t5 Y.t4 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 VGND.t3 B.t1 Y.t0 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 VGND.t11 C.t4 Y.t11 VNB.t11 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 a_449_297.t1 B.t2 a_27_297.t1 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14 VPWR.t1 A.t6 a_27_297.t5 VPB.t9 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 Y.t1 B.t3 VGND.t2 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X16 Y.t2 B.t4 VGND.t1 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X17 Y.t10 C.t5 VGND.t10 VNB.t10 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X18 Y.t9 C.t6 VGND.t9 VNB.t9 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X19 a_27_297.t2 B.t5 a_449_297.t2 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X20 VGND.t0 B.t6 Y.t3 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X21 a_449_297.t3 B.t7 a_27_297.t3 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X22 VGND.t8 C.t7 Y.t8 VNB.t8 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X23 a_27_297.t4 A.t7 VPWR.t0 VPB.t8 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
R0 A.n0 A.t7 212.079
R1 A.n2 A.t0 212.079
R2 A.n5 A.t2 212.079
R3 A.n8 A.t6 212.079
R4 A.n0 A.t5 139.779
R5 A.n2 A.t1 139.779
R6 A.n5 A.t3 139.779
R7 A.n8 A.t4 139.779
R8 A.n4 A.n1 96.723
R9 A A.n9 77.828
R10 A.n4 A.n3 76
R11 A.n7 A.n6 76
R12 A.n1 A.n0 21.909
R13 A.n7 A.n4 20.723
R14 A A.n7 18.895
R15 A.n9 A.n8 13.145
R16 A.n3 A.n2 10.224
R17 A.n6 A.n5 1.46
R18 a_27_297.t0 a_27_297.n5 223.217
R19 a_27_297.n3 a_27_297.t5 181.527
R20 a_27_297.n5 a_27_297.n0 156.927
R21 a_27_297.n3 a_27_297.n2 110.76
R22 a_27_297.n4 a_27_297.n1 92.444
R23 a_27_297.n4 a_27_297.n3 61.667
R24 a_27_297.n5 a_27_297.n4 28.87
R25 a_27_297.n2 a_27_297.t7 26.595
R26 a_27_297.n2 a_27_297.t6 26.595
R27 a_27_297.n1 a_27_297.t3 26.595
R28 a_27_297.n1 a_27_297.t4 26.595
R29 a_27_297.n0 a_27_297.t1 26.595
R30 a_27_297.n0 a_27_297.t2 26.595
R31 VPWR.n2 VPWR.n0 175.6
R32 VPWR.n2 VPWR.n1 175.407
R33 VPWR.n0 VPWR.t0 26.595
R34 VPWR.n0 VPWR.t3 26.595
R35 VPWR.n1 VPWR.t2 26.595
R36 VPWR.n1 VPWR.t1 26.595
R37 VPWR VPWR.n2 0.225
R38 VPB.t4 VPB.t0 248.598
R39 VPB.t5 VPB.t4 248.598
R40 VPB.t6 VPB.t5 248.598
R41 VPB.t7 VPB.t6 248.598
R42 VPB.t1 VPB.t7 248.598
R43 VPB.t2 VPB.t1 248.598
R44 VPB.t3 VPB.t2 248.598
R45 VPB.t8 VPB.t3 248.598
R46 VPB.t11 VPB.t8 248.598
R47 VPB.t10 VPB.t11 248.598
R48 VPB.t9 VPB.t10 248.598
R49 VPB VPB.t9 201.246
R50 C.n0 C.t0 212.079
R51 C.n2 C.t1 212.079
R52 C.n4 C.t2 212.079
R53 C.n3 C.t3 212.079
R54 C.n0 C.t6 139.779
R55 C.n2 C.t7 139.779
R56 C.n4 C.t5 139.779
R57 C.n3 C.t4 139.779
R58 C C.n1 92
R59 C C.n5 81.76
R60 C.n4 C.n3 61.345
R61 C.n5 C.n4 51.121
R62 C.n1 C.n0 21.909
R63 C.n5 C.n2 10.224
R64 Y.n2 Y.n1 343.865
R65 Y.n2 Y.n0 292.5
R66 Y Y.n2 98.757
R67 Y.n5 Y.n3 88.89
R68 Y Y.n13 66.206
R69 Y.n5 Y.n4 52.624
R70 Y.n7 Y.n6 52.624
R71 Y.n9 Y.n8 52.624
R72 Y.n11 Y.n10 52.624
R73 Y.n13 Y.n12 52.624
R74 Y.n7 Y.n5 36.266
R75 Y.n9 Y.n7 36.266
R76 Y.n11 Y.n9 36.266
R77 Y.n13 Y.n11 36.266
R78 Y.n0 Y.t15 26.595
R79 Y.n0 Y.t14 26.595
R80 Y.n1 Y.t13 26.595
R81 Y.n1 Y.t12 26.595
R82 Y.n3 Y.t6 24.923
R83 Y.n3 Y.t5 24.923
R84 Y.n4 Y.t4 24.923
R85 Y.n4 Y.t7 24.923
R86 Y.n6 Y.t0 24.923
R87 Y.n6 Y.t1 24.923
R88 Y.n8 Y.t11 24.923
R89 Y.n8 Y.t2 24.923
R90 Y.n10 Y.t8 24.923
R91 Y.n10 Y.t10 24.923
R92 Y.n12 Y.t3 24.923
R93 Y.n12 Y.t9 24.923
R94 a_449_297.n3 a_449_297.n2 360.928
R95 a_449_297.n4 a_449_297.n0 346.619
R96 a_449_297.n5 a_449_297.n4 292.5
R97 a_449_297.n3 a_449_297.n1 90.234
R98 a_449_297.n4 a_449_297.n3 69.798
R99 a_449_297.n1 a_449_297.t4 26.595
R100 a_449_297.n1 a_449_297.t1 26.595
R101 a_449_297.n2 a_449_297.t2 26.595
R102 a_449_297.n2 a_449_297.t3 26.595
R103 a_449_297.n0 a_449_297.t0 26.595
R104 a_449_297.n0 a_449_297.t7 26.595
R105 a_449_297.t6 a_449_297.n5 26.595
R106 a_449_297.n5 a_449_297.t5 26.595
R107 B.n4 B.n0 276.29
R108 B.n0 B.t0 236.179
R109 B.n1 B.t2 212.079
R110 B.n2 B.t5 212.079
R111 B.n5 B.t7 212.079
R112 B.n0 B.t6 163.879
R113 B.n1 B.t4 139.779
R114 B.n2 B.t1 139.779
R115 B.n5 B.t3 139.779
R116 B B.n6 87.58
R117 B.n4 B.n3 76
R118 B.n3 B.n1 59.884
R119 B.n6 B.n5 13.145
R120 B B.n4 9.142
R121 B.n3 B.n2 1.46
R122 VGND.n0 VGND.t0 199.065
R123 VGND.n2 VGND.n1 115.464
R124 VGND.n8 VGND.n7 115.464
R125 VGND.n12 VGND.n11 115.464
R126 VGND.n18 VGND.n17 115.464
R127 VGND.n24 VGND.n23 115.464
R128 VGND.n29 VGND.t5 104.607
R129 VGND.n1 VGND.t9 24.923
R130 VGND.n1 VGND.t8 24.923
R131 VGND.n7 VGND.t10 24.923
R132 VGND.n7 VGND.t11 24.923
R133 VGND.n11 VGND.t1 24.923
R134 VGND.n11 VGND.t3 24.923
R135 VGND.n17 VGND.t2 24.923
R136 VGND.n17 VGND.t4 24.923
R137 VGND.n23 VGND.t7 24.923
R138 VGND.n23 VGND.t6 24.923
R139 VGND.n9 VGND.n8 14.305
R140 VGND.n13 VGND.n12 14.305
R141 VGND.n3 VGND.n2 8.282
R142 VGND.n19 VGND.n18 8.282
R143 VGND.n30 VGND.n29 4.65
R144 VGND.n4 VGND.n3 4.65
R145 VGND.n6 VGND.n5 4.65
R146 VGND.n10 VGND.n9 4.65
R147 VGND.n14 VGND.n13 4.65
R148 VGND.n16 VGND.n15 4.65
R149 VGND.n20 VGND.n19 4.65
R150 VGND.n22 VGND.n21 4.65
R151 VGND.n26 VGND.n25 4.65
R152 VGND.n28 VGND.n27 4.65
R153 VGND.n25 VGND.n24 2.258
R154 VGND.n4 VGND.n0 0.551
R155 VGND.n6 VGND.n4 0.119
R156 VGND.n10 VGND.n6 0.119
R157 VGND.n14 VGND.n10 0.119
R158 VGND.n16 VGND.n14 0.119
R159 VGND.n20 VGND.n16 0.119
R160 VGND.n22 VGND.n20 0.119
R161 VGND.n26 VGND.n22 0.119
R162 VGND.n28 VGND.n26 0.119
R163 VGND.n30 VGND.n28 0.119
R164 VGND VGND.n30 0.02
R165 VNB VNB.t5 6150.61
R166 VNB.t9 VNB.t0 2030.77
R167 VNB.t8 VNB.t9 2030.77
R168 VNB.t10 VNB.t8 2030.77
R169 VNB.t11 VNB.t10 2030.77
R170 VNB.t1 VNB.t11 2030.77
R171 VNB.t3 VNB.t1 2030.77
R172 VNB.t2 VNB.t3 2030.77
R173 VNB.t4 VNB.t2 2030.77
R174 VNB.t7 VNB.t4 2030.77
R175 VNB.t6 VNB.t7 2030.77
R176 VNB.t5 VNB.t6 2030.77
C0 B Y 0.81fF
C1 VPB VPWR 0.11fF
C2 Y VGND 1.44fF
C3 C Y 0.20fF
C4 B C 0.41fF
C5 A Y 0.25fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__nor3b_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__nor3b_1 C_N Y A B VGND VPWR VNB VPB
X0 VGND.t2 a_91_199.t2 Y.t1 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 Y.t0 B.t0 VGND.t0 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 VPWR.t1 A.t0 a_245_297.t1 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 a_91_199.t1 C_N.t0 VGND.t1 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 VGND.t3 A.t1 Y.t3 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 a_245_297.t0 B.t1 a_161_297.t1 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 a_91_199.t0 C_N.t1 VPWR.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7 a_161_297.t0 a_91_199.t3 Y.t2 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
R0 a_91_199.t0 a_91_199.n1 355.821
R1 a_91_199.n1 a_91_199.t1 252.293
R2 a_91_199.n1 a_91_199.n0 242.774
R3 a_91_199.n0 a_91_199.t3 234.801
R4 a_91_199.n0 a_91_199.t2 162.501
R5 Y.n2 Y.t2 247.323
R6 Y.n1 Y.n0 165.099
R7 Y.n1 Y.t1 85.942
R8  Y.n1 52.745
R9 Y.n0 Y.t3 24.923
R10 Y.n0 Y.t0 24.923
R11  Y.n2 7.584
R12 Y.n2 Y 1.863
R13 VGND.n2 VGND.n0 111.769
R14 VGND.n2 VGND.n1 68.164
R15 VGND.n1 VGND.t1 57.889
R16 VGND.n0 VGND.t0 24.923
R17 VGND.n0 VGND.t2 24.923
R18 VGND.n1 VGND.t3 24.672
R19 VGND VGND.n2 0.427
R20 VNB VNB.t2 7397.8
R21 VNB.t3 VNB.t1 2303.7
R22 VNB.t0 VNB.t3 2030.77
R23 VNB.t2 VNB.t0 2030.77
R24 B.n0 B.t1 241.534
R25 B.n0 B.t0 169.234
R26 B B.n0 77.754
R27 A.n0 A.t0 241.534
R28 A.n0 A.t1 169.234
R29 A A.n0 78.167
R30 a_245_297.t0 a_245_297.t1 53.19
R31 VPWR VPWR.n0 318.418
R32 VPWR.n0 VPWR.t0 96.154
R33 VPWR.n0 VPWR.t1 27.364
R34 VPB VPB.t1 346.261
R35 VPB.t3 VPB.t0 287.071
R36 VPB.t2 VPB.t3 248.598
R37 VPB.t1 VPB.t2 248.598
R38 C_N.n0 C_N.t1 201.368
R39 C_N.n0 C_N.t0 132.281
R40 C_N C_N.n0 78.58
R41 a_161_297.t0 a_161_297.t1 53.19
C0 A C_N 0.14fF
C1 Y VGND 0.35fF
C2 B A 0.16fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__nor3b_2.ext - technology: sky130A

.subckt sky130_fd_sc_hd__nor3b_2 C_N Y A B VGND VPWR VNB VPB
X0 a_281_297.t3 B.t0 a_27_297.t3 VPB.t6 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 Y.t7 B.t1 VGND.t6 VNB.t6 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 a_27_297.t1 A.t0 VPWR.t1 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 VGND.t2 a_531_21.t2 Y.t2 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 VPWR.t2 C_N.t0 a_531_21.t0 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 VGND.t0 A.t1 Y.t0 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 Y.t1 A.t2 VGND.t1 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 VGND.t5 B.t2 Y.t6 VNB.t5 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 VPWR.t0 A.t3 a_27_297.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 a_281_297.t0 a_531_21.t3 Y.t3 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 Y.t4 a_531_21.t4 a_281_297.t1 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 VGND.t3 C_N.t1 a_531_21.t1 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12 a_27_297.t2 B.t3 a_281_297.t2 VPB.t5 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13 Y.t5 a_531_21.t5 VGND.t4 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
R0 B.n0 B.t3 212.079
R1 B.n1 B.t0 212.079
R2 B.n0 B.t2 139.779
R3 B.n1 B.t1 139.779
R4 B B.n2 76.304
R5 B.n2 B.n0 32.863
R6 B.n2 B.n1 28.481
R7  B 28.038
R8 a_27_297.n1 a_27_297.t2 225.591
R9 a_27_297.t0 a_27_297.n1 179.122
R10 a_27_297.n1 a_27_297.n0 110.76
R11 a_27_297.n0 a_27_297.t3 26.595
R12 a_27_297.n0 a_27_297.t1 26.595
R13 a_281_297.n1 a_281_297.n0 208.03
R14 a_281_297.n0 a_281_297.t0 182.039
R15 a_281_297.n0 a_281_297.t1 136.406
R16 a_281_297.t2 a_281_297.n1 26.595
R17 a_281_297.n1 a_281_297.t3 26.595
R18 VPB.t1 VPB.t2 580.062
R19 VPB.t5 VPB.t3 580.062
R20 VPB.t3 VPB.t1 248.598
R21 VPB.t6 VPB.t5 248.598
R22 VPB.t4 VPB.t6 248.598
R23 VPB.t0 VPB.t4 248.598
R24 VPB VPB.t0 201.246
R25 VGND.n7 VGND.t5 170.961
R26 VGND.n4 VGND.t4 170.961
R27 VGND.n1 VGND.t3 164.283
R28 VGND.n13 VGND.n12 115.464
R29 VGND.n0 VGND.t2 112.018
R30 VGND.n18 VGND.t1 104.607
R31 VGND.n12 VGND.t6 24.923
R32 VGND.n12 VGND.t0 24.923
R33 VGND.n19 VGND.n18 4.65
R34 VGND.n3 VGND.n2 4.65
R35 VGND.n6 VGND.n5 4.65
R36 VGND.n9 VGND.n8 4.65
R37 VGND.n11 VGND.n10 4.65
R38 VGND.n15 VGND.n14 4.65
R39 VGND.n17 VGND.n16 4.65
R40 VGND.n1 VGND.n0 4.034
R41 VGND.n14 VGND.n13 2.258
R42 VGND.n8 VGND.n7 2.2
R43 VGND.n3 VGND.n1 0.21
R44 VGND.n5 VGND.n4 0.2
R45 VGND.n6 VGND.n3 0.119
R46 VGND.n9 VGND.n6 0.119
R47 VGND.n11 VGND.n9 0.119
R48 VGND.n15 VGND.n11 0.119
R49 VGND.n17 VGND.n15 0.119
R50 VGND.n19 VGND.n17 0.119
R51 VGND VGND.n19 0.02
R52 Y.n4 Y.n3 190.575
R53 Y Y.n6 93.857
R54 Y.n2 Y.n0 88.89
R55 Y.n4 Y.n2 76.088
R56 Y.n2 Y.n1 52.624
R57 Y.n3 Y.t3 26.595
R58 Y.n3 Y.t4 26.595
R59 Y.n6 Y.t2 24.923
R60 Y.n6 Y.t5 24.923
R61 Y.n0 Y.t0 24.923
R62 Y.n0 Y.t1 24.923
R63 Y.n1 Y.t6 24.923
R64 Y.n1 Y.t7 24.923
R65 Y Y.n5 11.83
R66 Y.n5 Y.n4 3.296
R67 VNB VNB.t1 6150.61
R68 VNB.t2 VNB.t3 5548
R69 VNB.t5 VNB.t4 4738.46
R70 VNB.t4 VNB.t2 2030.77
R71 VNB.t6 VNB.t5 2030.77
R72 VNB.t0 VNB.t6 2030.77
R73 VNB.t1 VNB.t0 2030.77
R74 A.n0 A.t0 212.079
R75 A.n1 A.t3 212.079
R76 A.n0 A.t1 139.779
R77 A.n1 A.t2 139.779
R78 A A.n2 78.133
R79 A.n2 A.n0 38.706
R80  A 28.038
R81 A.n2 A.n1 22.639
R82 VPWR.n1 VPWR.t2 412.683
R83 VPWR.n1 VPWR.n0 175.493
R84 VPWR.n0 VPWR.t1 26.595
R85 VPWR.n0 VPWR.t0 26.595
R86 VPWR VPWR.n1 0.142
R87 a_531_21.t0 a_531_21.n2 377.635
R88 a_531_21.n1 a_531_21.t3 212.079
R89 a_531_21.n0 a_531_21.t4 212.079
R90 a_531_21.n2 a_531_21.t1 152.704
R91 a_531_21.n1 a_531_21.t2 139.779
R92 a_531_21.n0 a_531_21.t5 139.779
R93 a_531_21.n2 a_531_21.n1 135.372
R94 a_531_21.n1 a_531_21.n0 61.345
R95 C_N.n0 C_N.t0 147.813
R96 C_N.n0 C_N.t1 131.746
R97 C_N C_N.n0 81.485
C0 A Y 0.10fF
C1 VPWR VGND 0.10fF
C2 B Y 0.38fF
C3 VPB VPWR 0.10fF
C4 Y VGND 0.84fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__nor3b_4.ext - technology: sky130A

.subckt sky130_fd_sc_hd__nor3b_4 A C_N B Y VGND VPWR VNB VPB
X0 Y.t3 B.t0 VGND.t4 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 VPWR.t4 A.t0 a_197_297.t7 VPB.t8 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 Y.t8 a_27_47.t2 VGND.t9 VNB.t9 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 VGND.t5 A.t1 Y.t4 VNB.t5 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 a_555_297.t7 a_27_47.t3 Y.t9 VPB.t9 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 a_197_297.t6 A.t2 VPWR.t3 VPB.t7 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 VGND.t10 a_27_47.t4 Y.t10 VNB.t10 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 a_197_297.t3 B.t1 a_555_297.t3 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 VGND.t11 a_27_47.t5 Y.t11 VNB.t11 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 VGND.t3 B.t2 Y.t2 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 Y.t5 A.t3 VGND.t6 VNB.t6 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 VGND.t0 C_N.t0 a_27_47.t0 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 Y.t6 A.t4 VGND.t7 VNB.t7 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 Y.t12 a_27_47.t6 a_555_297.t6 VPB.t10 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14 Y.t13 a_27_47.t7 a_555_297.t5 VPB.t11 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 VPWR.t0 C_N.t1 a_27_47.t1 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16 a_555_297.t4 a_27_47.t8 Y.t14 VPB.t12 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17 VGND.t8 A.t5 Y.t7 VNB.t8 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X18 a_555_297.t2 B.t3 a_197_297.t2 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X19 a_197_297.t1 B.t4 a_555_297.t1 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X20 VGND.t2 B.t5 Y.t1 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X21 a_555_297.t0 B.t6 a_197_297.t0 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X22 VPWR.t2 A.t6 a_197_297.t5 VPB.t6 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X23 a_197_297.t4 A.t7 VPWR.t1 VPB.t5 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X24 Y.t0 B.t7 VGND.t1 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X25 Y.t15 a_27_47.t9 VGND.t12 VNB.t12 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
R0 B.n0 B.t3 212.079
R1 B.n1 B.t4 212.079
R2 B.n2 B.t6 212.079
R3 B.n4 B.t1 212.079
R4 B.n0 B.t2 139.779
R5 B.n1 B.t0 139.779
R6 B.n2 B.t5 139.779
R7 B.n4 B.t7 139.779
R8 B B.n5 87.58
R9 B.n1 B.n0 61.345
R10 B B.n3 42.198
R11 B.n3 B.n1 31.824
R12 B.n3 B.n2 18.432
R13 B.n5 B.n4 13.145
R14 VGND.n0 VGND.t11 200.093
R15 VGND.n2 VGND.n1 115.464
R16 VGND.n8 VGND.n7 115.464
R17 VGND.n12 VGND.n11 115.464
R18 VGND.n28 VGND.n27 115.464
R19 VGND.n34 VGND.n33 115.464
R20 VGND.n18 VGND.n17 92.5
R21 VGND.n22 VGND.n21 92.5
R22 VGND.n17 VGND.t1 24.923
R23 VGND.n21 VGND.t8 24.923
R24 VGND.n1 VGND.t12 24.923
R25 VGND.n1 VGND.t10 24.923
R26 VGND.n7 VGND.t9 24.923
R27 VGND.n7 VGND.t3 24.923
R28 VGND.n11 VGND.t4 24.923
R29 VGND.n11 VGND.t2 24.923
R30 VGND.n27 VGND.t7 24.923
R31 VGND.n27 VGND.t5 24.923
R32 VGND.n33 VGND.t6 24.923
R33 VGND.n33 VGND.t0 24.923
R34 VGND.n9 VGND.n8 15.811
R35 VGND.n13 VGND.n12 12.8
R36 VGND.n3 VGND.n2 9.788
R37 VGND.n29 VGND.n28 5.27
R38 VGND.n35 VGND.n34 4.899
R39 VGND.n4 VGND.n3 4.65
R40 VGND.n6 VGND.n5 4.65
R41 VGND.n10 VGND.n9 4.65
R42 VGND.n14 VGND.n13 4.65
R43 VGND.n16 VGND.n15 4.65
R44 VGND.n20 VGND.n19 4.65
R45 VGND.n24 VGND.n23 4.65
R46 VGND.n26 VGND.n25 4.65
R47 VGND.n30 VGND.n29 4.65
R48 VGND.n32 VGND.n31 4.65
R49 VGND.n23 VGND.n22 3
R50 VGND.n19 VGND.n18 2.076
R51 VGND.n4 VGND.n0 0.534
R52 VGND.n35 VGND.n32 0.132
R53 VGND VGND.n35 0.127
R54 VGND.n6 VGND.n4 0.119
R55 VGND.n10 VGND.n6 0.119
R56 VGND.n14 VGND.n10 0.119
R57 VGND.n16 VGND.n14 0.119
R58 VGND.n20 VGND.n16 0.119
R59 VGND.n24 VGND.n20 0.119
R60 VGND.n26 VGND.n24 0.119
R61 VGND.n30 VGND.n26 0.119
R62 VGND.n32 VGND.n30 0.119
R63 Y.n2 Y.n0 198.996
R64 Y.n2 Y.n1 154.573
R65 Y.n5 Y.n3 88.89
R66 Y.n7 Y.n5 73.244
R67 Y.n14 Y.n13 56.805
R68 Y.n5 Y.n4 52.624
R69 Y.n7 Y.n6 52.624
R70 Y.n9 Y.n8 52.624
R71 Y.n11 Y.n10 52.624
R72 Y.n13 Y.n12 52.624
R73 Y.n9 Y.n7 36.266
R74 Y.n11 Y.n9 36.266
R75 Y.n13 Y.n11 36.266
R76 Y.n14 Y.n2 34.258
R77 Y.n0 Y.t14 26.595
R78 Y.n0 Y.t13 26.595
R79 Y.n1 Y.t9 26.595
R80 Y.n1 Y.t12 26.595
R81 Y.n3 Y.t4 24.923
R82 Y.n3 Y.t5 24.923
R83 Y.n4 Y.t7 24.923
R84 Y.n4 Y.t6 24.923
R85 Y.n6 Y.t1 24.923
R86 Y.n6 Y.t0 24.923
R87 Y.n8 Y.t2 24.923
R88 Y.n8 Y.t3 24.923
R89 Y.n10 Y.t10 24.923
R90 Y.n10 Y.t8 24.923
R91 Y.n12 Y.t11 24.923
R92 Y.n12 Y.t15 24.923
R93 Y Y.n14 13.19
R94 VNB VNB.t0 6150.61
R95 VNB.t8 VNB.t1 4545.05
R96 VNB.t12 VNB.t11 2030.77
R97 VNB.t10 VNB.t12 2030.77
R98 VNB.t9 VNB.t10 2030.77
R99 VNB.t3 VNB.t9 2030.77
R100 VNB.t4 VNB.t3 2030.77
R101 VNB.t2 VNB.t4 2030.77
R102 VNB.t1 VNB.t2 2030.77
R103 VNB.t7 VNB.t8 2030.77
R104 VNB.t5 VNB.t7 2030.77
R105 VNB.t6 VNB.t5 2030.77
R106 VNB.t0 VNB.t6 2030.77
R107 A.n0 A.t6 212.079
R108 A.n3 A.t7 212.079
R109 A.n7 A.t0 212.079
R110 A.n6 A.t2 212.079
R111 A.n0 A.t5 139.779
R112 A.n3 A.t4 139.779
R113 A.n7 A.t1 139.779
R114 A.n6 A.t3 139.779
R115 A A.n8 87.58
R116 A.n2 A.n1 76
R117 A.n5 A.n4 76
R118 A.n7 A.n6 61.345
R119 A.n3 A.n2 39.436
R120 A.n1 A 26.209
R121 A.n2 A.n0 21.909
R122 A.n5 A 18.895
R123 A.n4 A.n3 10.224
R124 A A.n5 9.142
R125 A.n1 A 1.828
R126 A.n8 A.n7 1.46
R127 a_197_297.n4 a_197_297.n0 346.619
R128 a_197_297.n5 a_197_297.n4 292.5
R129 a_197_297.n3 a_197_297.n1 198.996
R130 a_197_297.n3 a_197_297.n2 154.573
R131 a_197_297.n4 a_197_297.n3 88.424
R132 a_197_297.n1 a_197_297.t7 26.595
R133 a_197_297.n1 a_197_297.t6 26.595
R134 a_197_297.n2 a_197_297.t5 26.595
R135 a_197_297.n2 a_197_297.t4 26.595
R136 a_197_297.n0 a_197_297.t2 26.595
R137 a_197_297.n0 a_197_297.t1 26.595
R138 a_197_297.t0 a_197_297.n5 26.595
R139 a_197_297.n5 a_197_297.t3 26.595
R140 VPWR.n2 VPWR.t2 557.228
R141 VPWR.n1 VPWR.n0 314.004
R142 VPWR.n6 VPWR.n5 171.981
R143 VPWR.n0 VPWR.t1 26.595
R144 VPWR.n0 VPWR.t4 26.595
R145 VPWR.n5 VPWR.t3 26.595
R146 VPWR.n5 VPWR.t0 26.595
R147 VPWR.n4 VPWR.n3 4.65
R148 VPWR.n7 VPWR.n6 4.024
R149 VPWR.n2 VPWR.n1 3.945
R150 VPWR.n4 VPWR.n2 0.272
R151 VPWR.n7 VPWR.n4 0.135
R152 VPWR VPWR.n7 0.123
R153 VPB.t6 VPB.t4 556.386
R154 VPB.t10 VPB.t9 248.598
R155 VPB.t12 VPB.t10 248.598
R156 VPB.t11 VPB.t12 248.598
R157 VPB.t3 VPB.t11 248.598
R158 VPB.t2 VPB.t3 248.598
R159 VPB.t1 VPB.t2 248.598
R160 VPB.t4 VPB.t1 248.598
R161 VPB.t5 VPB.t6 248.598
R162 VPB.t8 VPB.t5 248.598
R163 VPB.t7 VPB.t8 248.598
R164 VPB.t0 VPB.t7 248.598
R165 VPB VPB.t0 201.246
R166 a_27_47.n11 a_27_47.n10 323.799
R167 a_27_47.n0 a_27_47.t3 212.079
R168 a_27_47.n2 a_27_47.t6 212.079
R169 a_27_47.n5 a_27_47.t8 212.079
R170 a_27_47.n8 a_27_47.t7 212.079
R171 a_27_47.t1 a_27_47.n11 157.607
R172 a_27_47.n11 a_27_47.t0 149.854
R173 a_27_47.n0 a_27_47.t5 139.779
R174 a_27_47.n2 a_27_47.t9 139.779
R175 a_27_47.n5 a_27_47.t4 139.779
R176 a_27_47.n8 a_27_47.t2 139.779
R177 a_27_47.n4 a_27_47.n1 96.723
R178 a_27_47.n10 a_27_47.n9 76
R179 a_27_47.n4 a_27_47.n3 76
R180 a_27_47.n7 a_27_47.n6 76
R181 a_27_47.n1 a_27_47.n0 21.909
R182 a_27_47.n7 a_27_47.n4 20.723
R183 a_27_47.n10 a_27_47.n7 20.723
R184 a_27_47.n9 a_27_47.n8 13.145
R185 a_27_47.n3 a_27_47.n2 10.224
R186 a_27_47.n6 a_27_47.n5 1.46
R187 a_555_297.t3 a_555_297.n5 585.292
R188 a_555_297.n5 a_555_297.n4 292.5
R189 a_555_297.n1 a_555_297.t7 225.591
R190 a_555_297.n1 a_555_297.n0 154.573
R191 a_555_297.n3 a_555_297.n2 154.573
R192 a_555_297.n5 a_555_297.n3 49.271
R193 a_555_297.n3 a_555_297.n1 44.423
R194 a_555_297.n4 a_555_297.t1 26.595
R195 a_555_297.n4 a_555_297.t0 26.595
R196 a_555_297.n0 a_555_297.t6 26.595
R197 a_555_297.n0 a_555_297.t4 26.595
R198 a_555_297.n2 a_555_297.t5 26.595
R199 a_555_297.n2 a_555_297.t2 26.595
R200 C_N.n0 C_N.t1 229.558
R201 C_N.n0 C_N.t0 157.258
R202 C_N C_N.n0 83.619
C0 VPWR VGND 0.15fF
C1 A Y 0.34fF
C2 VPB VPWR 0.13fF
C3 Y VGND 1.50fF
C4 B Y 0.26fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__nor4_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__nor4_1 D C Y A B VGND VPWR VNB VPB
X0 Y.t2 B.t0 VGND.t2 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 a_191_297.t0 C.t0 a_109_297.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 VPWR.t0 A.t0 a_297_297.t0 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 VGND.t1 C.t1 Y.t1 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 VGND.t3 A.t1 Y.t3 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 a_297_297.t1 B.t1 a_191_297.t1 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 a_109_297.t1 D.t0 Y.t4 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 Y.t0 D.t1 VGND.t0 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
R0 B.n0 B.t1 241.534
R1 B.n0 B.t0 169.234
R2 B B.n0 112.721
R3 VGND.n5 VGND.t0 190.161
R4 VGND.n2 VGND.t3 190.026
R5 VGND.n1 VGND.n0 107.627
R6 VGND.n0 VGND.t1 25.846
R7 VGND.n0 VGND.t2 24.923
R8 VGND.n6 VGND.n5 4.65
R9 VGND.n4 VGND.n3 4.65
R10 VGND.n2 VGND.n1 3.704
R11 VGND.n4 VGND.n2 0.269
R12 VGND.n6 VGND.n4 0.119
R13 VGND VGND.n6 0.022
R14 Y.n2 Y.n1 167.228
R15 Y.n3 Y.t4 121.171
R16 Y.n2 Y.n0 97.088
R17 Y.n3 Y.n2 85.382
R18 Y.n0 Y.t0 42.461
R19 Y.n1 Y.t3 24.923
R20 Y.n1 Y.t2 24.923
R21 Y.n0 Y.t1 24.923
R22 Y Y.n3 7.358
R23 VNB VNB.t0 6078.09
R24 VNB.t0 VNB.t1 2490.11
R25 VNB.t1 VNB.t2 2054.95
R26 VNB.t2 VNB.t3 2030.77
R27 C.n0 C.t0 241.534
R28 C.n0 C.t1 169.234
R29 C C.n0 91.063
R30 a_109_297.t0 a_109_297.t1 51.22
R31 a_191_297.t0 a_191_297.t1 74.86
R32 VPB.t0 VPB.t2 313.707
R33 VPB.t2 VPB.t1 248.598
R34 VPB.t3 VPB.t0 242.679
R35 VPB VPB.t3 192.367
R36 A.n0 A.t0 230.154
R37 A.n0 A.t1 157.854
R38 A A.n0 95.446
R39 a_297_297.t0 a_297_297.t1 53.19
R40 VPWR VPWR.t0 200.117
R41 D.n0 D.t0 230.154
R42 D.n0 D.t1 157.854
R43 D D.n0 78.816
C0 C B 0.20fF
C1 Y VGND 0.22fF
C2 B VPWR 0.11fF
C3 D Y 0.13fF
C4 C Y 0.19fF
C5 B A 0.12fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__nor4_2.ext - technology: sky130A

.subckt sky130_fd_sc_hd__nor4_2 C D Y A B VGND VPWR VNB VPB
X0 a_281_297.t1 B.t0 a_27_297.t2 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 Y.t7 B.t1 VGND.t5 VNB.t5 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 a_27_297.t3 A.t0 VPWR.t1 VPB.t7 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 a_475_297.t1 D.t0 Y.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 VGND.t6 C.t0 Y.t8 VNB.t6 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 Y.t1 D.t1 a_475_297.t0 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 VGND.t0 D.t2 Y.t2 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 VGND.t2 A.t1 Y.t4 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 Y.t5 A.t2 VGND.t3 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 VGND.t4 B.t2 Y.t6 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 Y.t3 D.t3 VGND.t1 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 VPWR.t0 A.t3 a_27_297.t0 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 a_475_297.t2 C.t1 a_281_297.t2 VPB.t5 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13 a_281_297.t3 C.t2 a_475_297.t3 VPB.t6 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14 a_27_297.t1 B.t3 a_281_297.t0 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 Y.t9 C.t3 VGND.t7 VNB.t7 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
R0 B.n0 B.t3 212.079
R1 B.n1 B.t0 212.079
R2 B.n0 B.t2 139.779
R3 B.n1 B.t1 139.779
R4 B B.n2 76.874
R5 B.n2 B.n0 32.863
R6 B.n2 B.n1 28.481
R7 a_27_297.n1 a_27_297.t1 225.591
R8 a_27_297.t0 a_27_297.n1 181.528
R9 a_27_297.n1 a_27_297.n0 110.76
R10 a_27_297.n0 a_27_297.t2 26.595
R11 a_27_297.n0 a_27_297.t3 26.595
R12 a_281_297.n1 a_281_297.n0 395.733
R13 a_281_297.n0 a_281_297.t2 26.595
R14 a_281_297.n0 a_281_297.t3 26.595
R15 a_281_297.n1 a_281_297.t0 26.595
R16 a_281_297.t1 a_281_297.n1 26.595
R17 VPB.t3 VPB.t6 580.062
R18 VPB.t1 VPB.t0 248.598
R19 VPB.t5 VPB.t1 248.598
R20 VPB.t6 VPB.t5 248.598
R21 VPB.t4 VPB.t3 248.598
R22 VPB.t7 VPB.t4 248.598
R23 VPB.t2 VPB.t7 248.598
R24 VPB VPB.t2 201.246
R25 VGND.n2 VGND.t0 192.017
R26 VGND.n8 VGND.t4 165.357
R27 VGND.n5 VGND.t7 165.357
R28 VGND.n1 VGND.n0 115.464
R29 VGND.n14 VGND.n13 115.464
R30 VGND.n19 VGND.t3 104.607
R31 VGND.n0 VGND.t1 24.923
R32 VGND.n0 VGND.t6 24.923
R33 VGND.n13 VGND.t5 24.923
R34 VGND.n13 VGND.t2 24.923
R35 VGND.n2 VGND.n1 10.817
R36 VGND.n20 VGND.n19 4.65
R37 VGND.n4 VGND.n3 4.65
R38 VGND.n7 VGND.n6 4.65
R39 VGND.n10 VGND.n9 4.65
R40 VGND.n12 VGND.n11 4.65
R41 VGND.n16 VGND.n15 4.65
R42 VGND.n18 VGND.n17 4.65
R43 VGND.n15 VGND.n14 2.258
R44 VGND.n9 VGND.n8 2.2
R45 VGND.n4 VGND.n2 0.228
R46 VGND.n6 VGND.n5 0.2
R47 VGND.n7 VGND.n4 0.119
R48 VGND.n10 VGND.n7 0.119
R49 VGND.n12 VGND.n10 0.119
R50 VGND.n16 VGND.n12 0.119
R51 VGND.n18 VGND.n16 0.119
R52 VGND.n20 VGND.n18 0.119
R53 VGND VGND.n20 0.02
R54 Y.n8 Y.n7 202.979
R55 Y.n2 Y.n0 88.89
R56 Y.n4 Y.n2 76.088
R57 Y.n2 Y.n1 52.624
R58 Y.n4 Y.n3 52.624
R59 Y.n6 Y.n5 52.624
R60 Y.n6 Y.n4 36.266
R61 Y.n7 Y.t0 26.595
R62 Y.n7 Y.t1 26.595
R63 Y.n0 Y.t4 24.923
R64 Y.n0 Y.t5 24.923
R65 Y.n1 Y.t6 24.923
R66 Y.n1 Y.t7 24.923
R67 Y.n3 Y.t8 24.923
R68 Y.n3 Y.t9 24.923
R69 Y.n5 Y.t2 24.923
R70 Y.n5 Y.t3 24.923
R71 Y.n8 Y.n6 16.711
R72 Y Y.n8 1.91
R73 VNB VNB.t3 6150.61
R74 VNB.t4 VNB.t7 4738.46
R75 VNB.t1 VNB.t0 2030.77
R76 VNB.t6 VNB.t1 2030.77
R77 VNB.t7 VNB.t6 2030.77
R78 VNB.t5 VNB.t4 2030.77
R79 VNB.t2 VNB.t5 2030.77
R80 VNB.t3 VNB.t2 2030.77
R81 A.n0 A.t0 212.079
R82 A.n1 A.t3 212.079
R83 A.n0 A.t1 139.779
R84 A.n1 A.t2 139.779
R85 A A.n2 76.92
R86 A.n2 A.n0 38.706
R87 A.n2 A.n1 22.639
R88 VPWR VPWR.n0 175.636
R89 VPWR.n0 VPWR.t1 26.595
R90 VPWR.n0 VPWR.t0 26.595
R91 D.n0 D.t0 212.079
R92 D.n1 D.t1 212.079
R93 D.n0 D.t2 139.779
R94 D.n1 D.t3 139.779
R95 D D.n2 98.552
R96 D.n2 D.n0 33.593
R97 D.n2 D.n1 27.751
R98 a_475_297.n1 a_475_297.t3 246.119
R99 a_475_297.t1 a_475_297.n1 246.117
R100 a_475_297.n1 a_475_297.n0 90.234
R101 a_475_297.n0 a_475_297.t0 26.595
R102 a_475_297.n0 a_475_297.t2 26.595
R103 C.n0 C.t1 212.079
R104 C.n1 C.t2 212.079
R105 C.n0 C.t0 139.779
R106 C.n1 C.t3 139.779
R107 C C.n2 104.647
R108 C.n2 C.n0 30.672
R109 C.n2 C.n1 30.672
C0 C Y 0.17fF
C1 Y VGND 1.09fF
C2 D Y 0.19fF
C3 B Y 0.17fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__nor4_4.ext - technology: sky130A

.subckt sky130_fd_sc_hd__nor4_4 A C Y D B VGND VPWR VNB VPB
X0 VPWR.t3 A.t0 a_27_297.t3 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_807_297.t7 D.t0 Y.t15 VPB.t12 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 VGND.t15 C.t0 Y.t9 VNB.t15 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 Y.t3 A.t1 VGND.t3 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 Y.t14 D.t1 a_807_297.t6 VPB.t13 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 a_27_297.t2 A.t2 VPWR.t2 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 Y.t11 C.t1 VGND.t14 VNB.t14 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 Y.t19 D.t2 VGND.t11 VNB.t11 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 Y.t10 C.t2 VGND.t13 VNB.t13 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 Y.t18 D.t3 VGND.t10 VNB.t10 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 VGND.t2 A.t3 Y.t2 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 a_27_297.t4 B.t0 a_449_297.t3 VPB.t6 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 Y.t1 A.t4 VGND.t1 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 VGND.t0 A.t5 Y.t0 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14 VGND.t4 B.t1 Y.t5 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X15 VGND.t5 B.t2 Y.t6 VNB.t5 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X16 a_449_297.t2 B.t3 a_27_297.t5 VPB.t7 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17 a_807_297.t2 C.t3 a_449_297.t7 VPB.t10 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X18 VGND.t9 D.t4 Y.t17 VNB.t9 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X19 VGND.t8 D.t5 Y.t16 VNB.t8 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X20 a_807_297.t3 C.t4 a_449_297.t6 VPB.t11 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X21 VPWR.t1 A.t6 a_27_297.t1 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X22 a_449_297.t5 C.t5 a_807_297.t0 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X23 Y.t7 B.t4 VGND.t6 VNB.t6 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X24 Y.t8 B.t5 VGND.t7 VNB.t7 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X25 a_449_297.t4 C.t6 a_807_297.t1 VPB.t5 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X26 a_27_297.t6 B.t6 a_449_297.t1 VPB.t8 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X27 a_807_297.t5 D.t6 Y.t13 VPB.t14 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X28 a_449_297.t0 B.t7 a_27_297.t7 VPB.t9 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X29 Y.t12 D.t7 a_807_297.t4 VPB.t15 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X30 a_27_297.t0 A.t7 VPWR.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X31 VGND.t12 C.t7 Y.t4 VNB.t12 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
R0 A.n0 A.t7 212.079
R1 A.n2 A.t0 212.079
R2 A.n7 A.t2 212.079
R3 A.n5 A.t6 212.079
R4 A.n0 A.t5 139.779
R5 A.n2 A.t1 139.779
R6 A.n7 A.t3 139.779
R7 A.n5 A.t4 139.779
R8 A.n9 A.n6 96.723
R9 A.n4 A.n1 96.723
R10 A.n4 A.n3 76
R11 A.n9 A.n8 76
R12 A.n1 A.n0 21.909
R13 A.n6 A.n5 13.145
R14 A A.n4 11.58
R15 A.n3 A.n2 10.224
R16 A A.n9 9.142
R17 A.n8 A.n7 1.46
R18 a_27_297.n1 a_27_297.t4 224.108
R19 a_27_297.n3 a_27_297.t1 179.121
R20 a_27_297.n1 a_27_297.n0 154.573
R21 a_27_297.n3 a_27_297.n2 110.76
R22 a_27_297.n5 a_27_297.n4 90.234
R23 a_27_297.n4 a_27_297.n1 64.951
R24 a_27_297.n4 a_27_297.n3 64.951
R25 a_27_297.n2 a_27_297.t3 26.595
R26 a_27_297.n2 a_27_297.t2 26.595
R27 a_27_297.n0 a_27_297.t5 26.595
R28 a_27_297.n0 a_27_297.t6 26.595
R29 a_27_297.n5 a_27_297.t7 26.595
R30 a_27_297.t0 a_27_297.n5 26.595
R31 VPWR.n2 VPWR.n0 175.6
R32 VPWR.n2 VPWR.n1 175.407
R33 VPWR.n0 VPWR.t0 26.595
R34 VPWR.n0 VPWR.t3 26.595
R35 VPWR.n1 VPWR.t2 26.595
R36 VPWR.n1 VPWR.t1 26.595
R37 VPWR VPWR.n2 0.225
R38 VPB.t6 VPB.t5 556.386
R39 VPB.t15 VPB.t14 248.598
R40 VPB.t12 VPB.t15 248.598
R41 VPB.t13 VPB.t12 248.598
R42 VPB.t10 VPB.t13 248.598
R43 VPB.t4 VPB.t10 248.598
R44 VPB.t11 VPB.t4 248.598
R45 VPB.t5 VPB.t11 248.598
R46 VPB.t7 VPB.t6 248.598
R47 VPB.t8 VPB.t7 248.598
R48 VPB.t9 VPB.t8 248.598
R49 VPB.t0 VPB.t9 248.598
R50 VPB.t3 VPB.t0 248.598
R51 VPB.t2 VPB.t3 248.598
R52 VPB.t1 VPB.t2 248.598
R53 VPB VPB.t1 201.246
R54 D.n0 D.t6 212.079
R55 D.n2 D.t7 212.079
R56 D.n6 D.t0 212.079
R57 D.n5 D.t1 212.079
R58 D.n0 D.t5 139.779
R59 D.n2 D.t3 139.779
R60 D.n6 D.t4 139.779
R61 D.n5 D.t2 139.779
R62 D.n4 D.n1 96.723
R63 D.n4 D.n3 76
R64 D D.n7 41.589
R65 D.n7 D.n5 30.363
R66 D.n1 D.n0 26.29
R67 D.n7 D.n6 19.893
R68 D.n3 D.n2 14.606
R69 D D.n4 12.19
R70 Y.n17 Y.n15 198.996
R71 Y.n17 Y.n16 154.573
R72 Y.n2 Y.n0 88.89
R73 Y.n8 Y.n6 73.244
R74 Y.n2 Y.n1 52.624
R75 Y.n4 Y.n3 52.624
R76 Y.n6 Y.n5 52.624
R77 Y.n8 Y.n7 52.624
R78 Y.n10 Y.n9 52.624
R79 Y.n12 Y.n11 52.624
R80 Y.n14 Y.n13 52.624
R81 Y.n18 Y.n17 52.44
R82 Y.n4 Y.n2 36.266
R83 Y.n6 Y.n4 36.266
R84 Y.n10 Y.n8 36.266
R85 Y.n12 Y.n10 36.266
R86 Y.n14 Y.n12 36.266
R87 Y.n15 Y.t15 26.595
R88 Y.n15 Y.t14 26.595
R89 Y.n16 Y.t13 26.595
R90 Y.n16 Y.t12 26.595
R91 Y.n0 Y.t2 24.923
R92 Y.n0 Y.t1 24.923
R93 Y.n1 Y.t0 24.923
R94 Y.n1 Y.t3 24.923
R95 Y.n3 Y.t5 24.923
R96 Y.n3 Y.t7 24.923
R97 Y.n5 Y.t6 24.923
R98 Y.n5 Y.t8 24.923
R99 Y.n7 Y.t9 24.923
R100 Y.n7 Y.t10 24.923
R101 Y.n9 Y.t4 24.923
R102 Y.n9 Y.t11 24.923
R103 Y.n11 Y.t17 24.923
R104 Y.n11 Y.t19 24.923
R105 Y.n13 Y.t16 24.923
R106 Y.n13 Y.t18 24.923
R107 Y.n18 Y.n14 14.222
R108 Y Y.n18 2.37
R109 a_807_297.n3 a_807_297.t5 225.591
R110 a_807_297.n1 a_807_297.t1 224.711
R111 a_807_297.n3 a_807_297.n2 154.573
R112 a_807_297.n1 a_807_297.n0 154.573
R113 a_807_297.n5 a_807_297.n4 154.572
R114 a_807_297.n4 a_807_297.n1 44.423
R115 a_807_297.n4 a_807_297.n3 44.423
R116 a_807_297.n2 a_807_297.t4 26.595
R117 a_807_297.n2 a_807_297.t7 26.595
R118 a_807_297.n0 a_807_297.t0 26.595
R119 a_807_297.n0 a_807_297.t3 26.595
R120 a_807_297.t6 a_807_297.n5 26.595
R121 a_807_297.n5 a_807_297.t2 26.595
R122 C.n0 C.t3 212.079
R123 C.n2 C.t5 212.079
R124 C.n5 C.t4 212.079
R125 C.n8 C.t6 212.079
R126 C.n0 C.t7 139.779
R127 C.n2 C.t1 139.779
R128 C.n5 C.t0 139.779
R129 C.n8 C.t2 139.779
R130 C.n4 C.n1 96.723
R131 C C.n9 93.676
R132 C.n4 C.n3 76
R133 C.n7 C.n6 76
R134 C.n1 C.n0 21.909
R135 C.n7 C.n4 20.723
R136 C.n9 C.n8 13.145
R137 C.n3 C.n2 10.224
R138 C C.n7 3.047
R139 C.n6 C.n5 1.46
R140 VGND.n0 VGND.t8 200.618
R141 VGND.n2 VGND.n1 115.464
R142 VGND.n8 VGND.n7 115.464
R143 VGND.n14 VGND.n13 115.464
R144 VGND.n28 VGND.n27 115.464
R145 VGND.n34 VGND.n33 115.464
R146 VGND.n40 VGND.n39 115.464
R147 VGND.n45 VGND.t1 104.607
R148 VGND.n20 VGND.n19 92.5
R149 VGND.n22 VGND.n21 92.5
R150 VGND.n19 VGND.t13 24.923
R151 VGND.n21 VGND.t5 24.923
R152 VGND.n1 VGND.t10 24.923
R153 VGND.n1 VGND.t9 24.923
R154 VGND.n7 VGND.t11 24.923
R155 VGND.n7 VGND.t12 24.923
R156 VGND.n13 VGND.t14 24.923
R157 VGND.n13 VGND.t15 24.923
R158 VGND.n27 VGND.t7 24.923
R159 VGND.n27 VGND.t4 24.923
R160 VGND.n33 VGND.t6 24.923
R161 VGND.n33 VGND.t0 24.923
R162 VGND.n39 VGND.t3 24.923
R163 VGND.n39 VGND.t2 24.923
R164 VGND.n29 VGND.n28 14.305
R165 VGND.n15 VGND.n14 12.8
R166 VGND.n35 VGND.n34 8.282
R167 VGND.n9 VGND.n8 6.776
R168 VGND.n23 VGND.n22 5.4
R169 VGND.n23 VGND.n20 5
R170 VGND.n46 VGND.n45 4.65
R171 VGND.n4 VGND.n3 4.65
R172 VGND.n6 VGND.n5 4.65
R173 VGND.n10 VGND.n9 4.65
R174 VGND.n12 VGND.n11 4.65
R175 VGND.n16 VGND.n15 4.65
R176 VGND.n18 VGND.n17 4.65
R177 VGND.n24 VGND.n23 4.65
R178 VGND.n26 VGND.n25 4.65
R179 VGND.n30 VGND.n29 4.65
R180 VGND.n32 VGND.n31 4.65
R181 VGND.n36 VGND.n35 4.65
R182 VGND.n38 VGND.n37 4.65
R183 VGND.n42 VGND.n41 4.65
R184 VGND.n44 VGND.n43 4.65
R185 VGND.n41 VGND.n40 2.258
R186 VGND.n4 VGND.n0 1.179
R187 VGND.n3 VGND.n2 0.752
R188 VGND.n6 VGND.n4 0.119
R189 VGND.n10 VGND.n6 0.119
R190 VGND.n12 VGND.n10 0.119
R191 VGND.n16 VGND.n12 0.119
R192 VGND.n18 VGND.n16 0.119
R193 VGND.n24 VGND.n18 0.119
R194 VGND.n26 VGND.n24 0.119
R195 VGND.n30 VGND.n26 0.119
R196 VGND.n32 VGND.n30 0.119
R197 VGND.n36 VGND.n32 0.119
R198 VGND.n38 VGND.n36 0.119
R199 VGND.n42 VGND.n38 0.119
R200 VGND.n44 VGND.n42 0.119
R201 VGND.n46 VGND.n44 0.119
R202 VGND VGND.n46 0.02
R203 VNB VNB.t1 6150.61
R204 VNB.t5 VNB.t13 4545.05
R205 VNB.t10 VNB.t8 2030.77
R206 VNB.t9 VNB.t10 2030.77
R207 VNB.t11 VNB.t9 2030.77
R208 VNB.t12 VNB.t11 2030.77
R209 VNB.t14 VNB.t12 2030.77
R210 VNB.t15 VNB.t14 2030.77
R211 VNB.t13 VNB.t15 2030.77
R212 VNB.t7 VNB.t5 2030.77
R213 VNB.t4 VNB.t7 2030.77
R214 VNB.t6 VNB.t4 2030.77
R215 VNB.t0 VNB.t6 2030.77
R216 VNB.t3 VNB.t0 2030.77
R217 VNB.t2 VNB.t3 2030.77
R218 VNB.t1 VNB.t2 2030.77
R219 B.n0 B.t0 212.079
R220 B.n3 B.t3 212.079
R221 B.n8 B.t6 212.079
R222 B.n6 B.t7 212.079
R223 B.n0 B.t2 139.779
R224 B.n3 B.t5 139.779
R225 B.n8 B.t1 139.779
R226 B.n6 B.t4 139.779
R227 B.n10 B.n7 96.723
R228 B.n2 B.n1 76
R229 B.n5 B.n4 76
R230 B.n10 B.n9 76
R231 B.n1 B.n0 21.909
R232 B.n5 B.n2 20.723
R233 B B.n10 18.895
R234 B.n7 B.n6 13.145
R235 B.n4 B.n3 10.224
R236 B.n2 B 5.485
R237 B B.n5 1.828
R238 B.n9 B.n8 1.46
R239 a_449_297.n3 a_449_297.n1 198.996
R240 a_449_297.n4 a_449_297.n0 198.996
R241 a_449_297.n3 a_449_297.n2 154.573
R242 a_449_297.n5 a_449_297.n4 154.572
R243 a_449_297.n4 a_449_297.n3 83.576
R244 a_449_297.n1 a_449_297.t7 26.595
R245 a_449_297.n1 a_449_297.t5 26.595
R246 a_449_297.n2 a_449_297.t6 26.595
R247 a_449_297.n2 a_449_297.t4 26.595
R248 a_449_297.n0 a_449_297.t1 26.595
R249 a_449_297.n0 a_449_297.t0 26.595
R250 a_449_297.t3 a_449_297.n5 26.595
R251 a_449_297.n5 a_449_297.t2 26.595
C0 B Y 0.41fF
C1 VPB VPWR 0.14fF
C2 VPWR VGND 0.16fF
C3 C Y 0.27fF
C4 Y VGND 1.92fF
C5 D Y 0.50fF
C6 A Y 0.25fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__nor4b_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__nor4b_1 C B A D_N Y VGND VPWR VNB VPB
X0 Y.t2 a_91_199.t2 VGND.t2 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 Y.t4 B.t0 VGND.t3 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 VGND.t0 C.t0 Y.t0 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 a_91_199.t1 D_N.t0 VGND.t4 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 VGND.t1 A.t0 Y.t1 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 VPWR.t0 A.t1 a_341_297.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 a_245_297.t0 C.t1 a_161_297.t1 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 a_341_297.t1 B.t1 a_245_297.t1 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 a_91_199.t0 D_N.t1 VPWR.t1 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9 a_161_297.t0 a_91_199.t3 Y.t3 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
R0 a_91_199.t0 a_91_199.n1 355.821
R1 a_91_199.n1 a_91_199.t1 245.66
R2 a_91_199.n1 a_91_199.n0 240.958
R3 a_91_199.n0 a_91_199.t3 234.801
R4 a_91_199.n0 a_91_199.t2 162.501
R5 VGND.n6 VGND.t2 192.177
R6 VGND.n1 VGND.n0 107.627
R7 VGND.n3 VGND.n2 68.636
R8 VGND.n2 VGND.t4 57.889
R9 VGND.n0 VGND.t3 30.461
R10 VGND.n0 VGND.t0 30.461
R11 VGND.n2 VGND.t1 24.672
R12 VGND.n3 VGND.n1 7.946
R13 VGND.n5 VGND.n4 4.65
R14 VGND.n8 VGND.n7 4.65
R15 VGND.n5 VGND.n3 0.461
R16 VGND.n7 VGND.n6 0.376
R17 VGND.n8 VGND.n5 0.119
R18 VGND.n9 VGND.n8 0.119
R19 VGND VGND.n9 0.022
R20 Y Y.t3 236.01
R21 Y.n2 Y.n0 158.627
R22 Y.n2 Y.n1 108.18
R23 Y Y.n2 89.846
R24 Y.n0 Y.t1 24.923
R25 Y.n0 Y.t4 24.923
R26 Y.n1 Y.t0 24.923
R27 Y.n1 Y.t2 24.923
R28 VNB VNB.t2 7832.97
R29 VNB.t0 VNB.t3 2320.88
R30 VNB.t1 VNB.t4 2303.7
R31 VNB.t3 VNB.t1 2030.77
R32 VNB.t2 VNB.t0 2030.77
R33 B.n0 B.t1 241.534
R34 B.n0 B.t0 169.234
R35 B B.n0 78.167
R36 C.n0 C.t1 241.534
R37 C.n0 C.t0 169.234
R38 C C.n0 77.754
R39 D_N.n0 D_N.t1 211.008
R40 D_N.n0 D_N.t0 132.281
R41 D_N D_N.n0 78.993
R42 A.n0 A.t1 241.534
R43 A.n0 A.t0 169.234
R44 A A.n0 78.58
R45 a_341_297.t0 a_341_297.t1 53.19
R46 VPWR VPWR.n0 317.031
R47 VPWR.n0 VPWR.t1 96.154
R48 VPWR.n0 VPWR.t0 27.964
R49 VPB VPB.t1 346.261
R50 VPB.t0 VPB.t2 287.071
R51 VPB.t3 VPB.t4 284.112
R52 VPB.t4 VPB.t0 248.598
R53 VPB.t1 VPB.t3 248.598
R54 a_161_297.t0 a_161_297.t1 53.19
R55 a_245_297.t0 a_245_297.t1 65.01
C0 A D_N 0.14fF
C1 C B 0.16fF
C2 Y VGND 0.43fF
C3 B A 0.16fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__nor4b_2.ext - technology: sky130A

.subckt sky130_fd_sc_hd__nor4b_2 D_N Y C A B VGND VPWR VNB VPB
X0 VPWR.t1 D_N.t0 a_694_21.t0 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1 a_27_297.t1 B.t0 a_277_297.t3 VPB.t7 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 a_474_297.t3 a_694_21.t2 Y.t5 VPB.t5 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 a_277_297.t2 B.t1 a_27_297.t0 VPB.t8 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 Y.t4 a_694_21.t3 a_474_297.t2 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 VGND.t3 C.t0 Y.t1 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 VGND.t4 D_N.t1 a_694_21.t1 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7 a_27_297.t2 A.t0 VPWR.t0 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 VGND.t7 A.t1 Y.t8 VNB.t7 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 VGND.t1 B.t2 Y.t3 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 Y.t0 C.t1 VGND.t2 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 a_474_297.t0 C.t2 a_277_297.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 Y.t2 B.t3 VGND.t0 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 Y.t7 a_694_21.t4 VGND.t6 VNB.t6 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14 a_277_297.t1 C.t3 a_474_297.t1 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 VGND.t5 a_694_21.t5 Y.t6 VNB.t5 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X16 VPWR.t2 A.t2 a_27_297.t3 VPB.t6 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17 Y.t9 A.t3 VGND.t8 VNB.t8 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
R0 D_N.n0 D_N.t0 334.186
R1 D_N.n0 D_N.t1 131.746
R2 D_N.n1 D_N.n0 89.104
R3  D_N.n1 13.568
R4 D_N.n1 D_N 3.84
R5 a_694_21.t0 a_694_21.n2 427.77
R6 a_694_21.n1 a_694_21.t2 212.079
R7 a_694_21.n0 a_694_21.t3 212.079
R8 a_694_21.n2 a_694_21.t1 156.157
R9 a_694_21.n2 a_694_21.n1 151.951
R10 a_694_21.n1 a_694_21.t5 139.779
R11 a_694_21.n0 a_694_21.t4 139.779
R12 a_694_21.n1 a_694_21.n0 61.345
R13 VPWR.n1 VPWR.t1 383.988
R14 VPWR.n1 VPWR.n0 180.409
R15 VPWR.n0 VPWR.t0 26.595
R16 VPWR.n0 VPWR.t2 26.595
R17 VPWR VPWR.n1 0.144
R18 VPB.t7 VPB.t1 577.102
R19 VPB.t5 VPB.t3 556.386
R20 VPB.t4 VPB.t5 248.598
R21 VPB.t0 VPB.t4 248.598
R22 VPB.t1 VPB.t0 248.598
R23 VPB.t8 VPB.t7 248.598
R24 VPB.t2 VPB.t8 248.598
R25 VPB.t6 VPB.t2 248.598
R26 VPB VPB.t6 192.367
R27 B.n0 B.t0 212.079
R28 B.n1 B.t1 212.079
R29 B.n0 B.t2 139.779
R30 B.n1 B.t3 139.779
R31 B.n3 B.n2 76
R32 B.n2 B.n1 40.166
R33  B.n3 23.466
R34 B.n2 B.n0 21.178
R35 B.n3 B 4.571
R36 a_277_297.n1 a_277_297.n0 404.495
R37 a_277_297.n0 a_277_297.t3 26.595
R38 a_277_297.n0 a_277_297.t2 26.595
R39 a_277_297.t0 a_277_297.n1 26.595
R40 a_277_297.n1 a_277_297.t1 26.595
R41 a_27_297.t1 a_27_297.n1 220.97
R42 a_27_297.n1 a_27_297.t3 175.728
R43 a_27_297.n1 a_27_297.n0 110.76
R44 a_27_297.n0 a_27_297.t0 26.595
R45 a_27_297.n0 a_27_297.t2 26.595
R46 Y.n1 Y.n0 155.668
R47 Y.n4 Y.n2 88.89
R48 Y.n6 Y.n4 75.733
R49 Y.n4 Y.n3 52.624
R50 Y.n6 Y.n5 52.624
R51 Y.n8 Y.n7 52.624
R52 Y.n8 Y.n6 36.266
R53 Y.n0 Y.t5 26.595
R54 Y.n0 Y.t4 26.595
R55 Y.n7 Y.t6 24.923
R56 Y.n7 Y.t7 24.923
R57 Y.n2 Y.t8 24.923
R58 Y.n2 Y.t9 24.923
R59 Y.n3 Y.t3 24.923
R60 Y.n3 Y.t2 24.923
R61 Y.n5 Y.t1 24.923
R62 Y.n5 Y.t0 24.923
R63  Y.n8 15.304
R64  Y 13.6
R65 Y Y.n1 0.4
R66 Y.n1 Y 0.316
R67 a_474_297.n0 a_474_297.t3 246.286
R68 a_474_297.n0 a_474_297.t1 240.549
R69 a_474_297.n1 a_474_297.n0 90.234
R70 a_474_297.t2 a_474_297.n1 26.595
R71 a_474_297.n1 a_474_297.t0 26.595
R72 C.n0 C.t2 212.079
R73 C.n1 C.t3 212.079
R74 C.n0 C.t0 139.779
R75 C.n1 C.t1 139.779
R76 C.n3 C.n2 76
R77 C.n2 C.n1 40.166
R78  C.n3 23.466
R79 C.n2 C.n0 21.178
R80 C.n3 C 4.571
R81 VGND.n13 VGND.t1 170.961
R82 VGND.n10 VGND.t2 170.961
R83 VGND.n1 VGND.t4 170.384
R84 VGND.n5 VGND.n4 115.464
R85 VGND.n19 VGND.n18 115.464
R86 VGND.n0 VGND.t5 114.83
R87 VGND.n24 VGND.t8 108.671
R88 VGND.n4 VGND.t6 24.923
R89 VGND.n4 VGND.t3 24.923
R90 VGND.n18 VGND.t0 24.923
R91 VGND.n18 VGND.t7 24.923
R92 VGND.n1 VGND.n0 9.615
R93 VGND.n6 VGND.n5 8.658
R94 VGND.n25 VGND.n24 4.65
R95 VGND.n3 VGND.n2 4.65
R96 VGND.n7 VGND.n6 4.65
R97 VGND.n9 VGND.n8 4.65
R98 VGND.n12 VGND.n11 4.65
R99 VGND.n15 VGND.n14 4.65
R100 VGND.n17 VGND.n16 4.65
R101 VGND.n21 VGND.n20 4.65
R102 VGND.n23 VGND.n22 4.65
R103 VGND.n20 VGND.n19 3.764
R104 VGND.n14 VGND.n13 2.6
R105 VGND.n11 VGND.n10 0.7
R106 VGND.n3 VGND.n1 0.302
R107 VGND.n7 VGND.n3 0.119
R108 VGND.n9 VGND.n7 0.119
R109 VGND.n12 VGND.n9 0.119
R110 VGND.n15 VGND.n12 0.119
R111 VGND.n17 VGND.n15 0.119
R112 VGND.n21 VGND.n17 0.119
R113 VGND.n23 VGND.n21 0.119
R114 VGND.n25 VGND.n23 0.119
R115 VGND VGND.n25 0.022
R116 VNB VNB.t8 6078.09
R117 VNB.t5 VNB.t4 5321.88
R118 VNB.t1 VNB.t2 4714.29
R119 VNB.t6 VNB.t5 2030.77
R120 VNB.t3 VNB.t6 2030.77
R121 VNB.t2 VNB.t3 2030.77
R122 VNB.t0 VNB.t1 2030.77
R123 VNB.t7 VNB.t0 2030.77
R124 VNB.t8 VNB.t7 2030.77
R125 A.n0 A.t0 212.079
R126 A.n1 A.t2 212.079
R127 A.n0 A.t1 139.779
R128 A.n1 A.t3 139.779
R129 A.n3 A.n2 76
R130 A.n2 A.n0 38.706
R131 A  28.038
R132  A.n3 25.904
R133 A.n2 A.n1 22.639
R134 A.n3 A 2.133
C0 VPWR VGND 0.12fF
C1 C Y 0.20fF
C2 Y VGND 1.06fF
C3 A Y 0.17fF
C4 B Y 0.29fF
C5 VPB VPWR 0.11fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__nor4b_4.ext - technology: sky130A

.subckt sky130_fd_sc_hd__nor4b_4 B A D_N C Y VGND VPWR VNB VPB
X0 VGND.t3 B.t0 Y.t3 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 VGND.t2 B.t1 Y.t2 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 VGND.t4 D_N.t0 a_1191_21.t0 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 a_803_297.t7 a_1191_21.t2 Y.t4 VPB.t12 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 a_445_297.t3 B.t2 a_27_297.t3 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 a_27_297.t5 A.t0 VPWR.t4 VPB.t14 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 Y.t5 a_1191_21.t3 a_803_297.t6 VPB.t11 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 a_803_297.t5 a_1191_21.t4 Y.t6 VPB.t10 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 Y.t12 C.t0 VGND.t9 VNB.t9 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 VPWR.t3 A.t1 a_27_297.t6 VPB.t15 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 Y.t7 a_1191_21.t5 a_803_297.t4 VPB.t9 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 Y.t13 C.t1 VGND.t10 VNB.t10 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 Y.t8 a_1191_21.t6 VGND.t5 VNB.t5 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 a_27_297.t7 A.t2 VPWR.t2 VPB.t16 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14 VPWR.t0 D_N.t1 a_1191_21.t1 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 VGND.t13 A.t3 Y.t16 VNB.t13 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X16 VGND.t14 A.t4 Y.t17 VNB.t14 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X17 VGND.t11 C.t2 Y.t14 VNB.t11 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X18 a_27_297.t2 B.t3 a_445_297.t2 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X19 VGND.t12 C.t3 Y.t15 VNB.t12 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X20 VGND.t6 a_1191_21.t7 Y.t9 VNB.t6 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X21 VGND.t7 a_1191_21.t8 Y.t10 VNB.t7 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X22 Y.t18 A.t5 VGND.t15 VNB.t15 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X23 Y.t1 B.t4 VGND.t1 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X24 a_445_297.t1 B.t5 a_27_297.t1 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X25 a_803_297.t0 C.t4 a_445_297.t4 VPB.t5 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X26 Y.t0 B.t6 VGND.t0 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X27 a_27_297.t0 B.t7 a_445_297.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X28 a_445_297.t5 C.t5 a_803_297.t1 VPB.t6 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X29 a_803_297.t2 C.t6 a_445_297.t6 VPB.t7 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X30 Y.t11 a_1191_21.t9 VGND.t8 VNB.t8 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X31 VPWR.t1 A.t6 a_27_297.t4 VPB.t13 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X32 a_445_297.t7 C.t7 a_803_297.t3 VPB.t8 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X33 Y.t19 A.t7 VGND.t16 VNB.t16 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
R0 B.n0 B.t3 212.079
R1 B.n2 B.t5 212.079
R2 B.n7 B.t7 212.079
R3 B.n5 B.t2 212.079
R4 B.n0 B.t1 139.779
R5 B.n2 B.t6 139.779
R6 B.n7 B.t0 139.779
R7 B.n5 B.t4 139.779
R8 B.n9 B.n6 96.723
R9 B.n4 B.n1 96.723
R10 B.n4 B.n3 76
R11 B.n9 B.n8 76
R12 B.n1 B.n0 21.909
R13 B B.n9 18.895
R14 B.n6 B.n5 13.145
R15 B.n3 B.n2 10.224
R16 B B.n4 1.828
R17 B.n8 B.n7 1.46
R18 Y.n16 Y.n0 191.467
R19 Y.n18 Y.n17 146.393
R20 Y.n15 Y.n1 97.068
R21 Y.n5 Y.n3 88.89
R22 Y.n11 Y.n9 73.244
R23 Y.n5 Y.n4 52.624
R24 Y.n7 Y.n6 52.624
R25 Y.n9 Y.n8 52.624
R26 Y.n11 Y.n10 52.624
R27 Y.n13 Y.n12 52.624
R28 Y.n14 Y.n2 49.285
R29 Y.n14 Y.n13 47.999
R30 Y.n7 Y.n5 36.266
R31 Y.n9 Y.n7 36.266
R32 Y.n13 Y.n11 36.266
R33 Y.n17 Y.t6 26.595
R34 Y.n17 Y.t7 26.595
R35 Y.n0 Y.t4 26.595
R36 Y.n0 Y.t5 26.595
R37 Y.n2 Y.t9 24.923
R38 Y.n2 Y.t8 24.923
R39 Y.n3 Y.t16 24.923
R40 Y.n3 Y.t19 24.923
R41 Y.n4 Y.t17 24.923
R42 Y.n4 Y.t18 24.923
R43 Y.n6 Y.t3 24.923
R44 Y.n6 Y.t1 24.923
R45 Y.n8 Y.t2 24.923
R46 Y.n8 Y.t0 24.923
R47 Y.n10 Y.t15 24.923
R48 Y.n10 Y.t13 24.923
R49 Y.n12 Y.t14 24.923
R50 Y.n12 Y.t12 24.923
R51 Y.n1 Y.t10 24.923
R52 Y.n1 Y.t11 24.923
R53 Y.n16 Y.n15 23.222
R54 Y.n18 Y.n16 6.992
R55 Y Y.n18 4.192
R56 Y.n15 Y.n14 3.555
R57 VGND.n0 VGND.t7 193.925
R58 VGND.n5 VGND.n4 115.464
R59 VGND.n11 VGND.n10 115.464
R60 VGND.n17 VGND.n16 115.464
R61 VGND.n31 VGND.n30 115.464
R62 VGND.n37 VGND.n36 115.464
R63 VGND.n43 VGND.n42 115.464
R64 VGND.n48 VGND.t16 114.4
R65 VGND.n1 VGND.t4 112.946
R66 VGND.n23 VGND.n22 92.5
R67 VGND.n25 VGND.n24 92.5
R68 VGND.n22 VGND.t10 24.923
R69 VGND.n24 VGND.t2 24.923
R70 VGND.n4 VGND.t8 24.923
R71 VGND.n4 VGND.t6 24.923
R72 VGND.n10 VGND.t5 24.923
R73 VGND.n10 VGND.t11 24.923
R74 VGND.n16 VGND.t9 24.923
R75 VGND.n16 VGND.t12 24.923
R76 VGND.n30 VGND.t0 24.923
R77 VGND.n30 VGND.t3 24.923
R78 VGND.n36 VGND.t1 24.923
R79 VGND.n36 VGND.t14 24.923
R80 VGND.n42 VGND.t15 24.923
R81 VGND.n42 VGND.t13 24.923
R82 VGND.n32 VGND.n31 15.811
R83 VGND.n18 VGND.n17 11.294
R84 VGND.n1 VGND.n0 10.842
R85 VGND.n38 VGND.n37 9.788
R86 VGND.n49 VGND.n48 6.908
R87 VGND.n26 VGND.n25 5.8
R88 VGND.n12 VGND.n11 5.27
R89 VGND.n3 VGND.n2 4.65
R90 VGND.n7 VGND.n6 4.65
R91 VGND.n9 VGND.n8 4.65
R92 VGND.n13 VGND.n12 4.65
R93 VGND.n15 VGND.n14 4.65
R94 VGND.n19 VGND.n18 4.65
R95 VGND.n21 VGND.n20 4.65
R96 VGND.n27 VGND.n26 4.65
R97 VGND.n29 VGND.n28 4.65
R98 VGND.n33 VGND.n32 4.65
R99 VGND.n35 VGND.n34 4.65
R100 VGND.n39 VGND.n38 4.65
R101 VGND.n41 VGND.n40 4.65
R102 VGND.n45 VGND.n44 4.65
R103 VGND.n47 VGND.n46 4.65
R104 VGND.n26 VGND.n23 4.6
R105 VGND.n44 VGND.n43 3.764
R106 VGND.n6 VGND.n5 0.752
R107 VGND.n3 VGND.n1 0.206
R108 VGND.n7 VGND.n3 0.119
R109 VGND.n9 VGND.n7 0.119
R110 VGND.n13 VGND.n9 0.119
R111 VGND.n15 VGND.n13 0.119
R112 VGND.n19 VGND.n15 0.119
R113 VGND.n21 VGND.n19 0.119
R114 VGND.n27 VGND.n21 0.119
R115 VGND.n29 VGND.n27 0.119
R116 VGND.n33 VGND.n29 0.119
R117 VGND.n35 VGND.n33 0.119
R118 VGND.n39 VGND.n35 0.119
R119 VGND.n41 VGND.n39 0.119
R120 VGND.n45 VGND.n41 0.119
R121 VGND.n47 VGND.n45 0.119
R122 VGND.n49 VGND.n47 0.119
R123 VGND VGND.n49 0.022
R124 VNB VNB.t16 6078.09
R125 VNB.t7 VNB.t4 4545.05
R126 VNB.t2 VNB.t10 4545.05
R127 VNB.t8 VNB.t7 2030.77
R128 VNB.t6 VNB.t8 2030.77
R129 VNB.t5 VNB.t6 2030.77
R130 VNB.t11 VNB.t5 2030.77
R131 VNB.t9 VNB.t11 2030.77
R132 VNB.t12 VNB.t9 2030.77
R133 VNB.t10 VNB.t12 2030.77
R134 VNB.t0 VNB.t2 2030.77
R135 VNB.t3 VNB.t0 2030.77
R136 VNB.t1 VNB.t3 2030.77
R137 VNB.t14 VNB.t1 2030.77
R138 VNB.t15 VNB.t14 2030.77
R139 VNB.t13 VNB.t15 2030.77
R140 VNB.t16 VNB.t13 2030.77
R141 D_N.n0 D_N.t1 231.716
R142 D_N.n0 D_N.t0 159.416
R143 D_N D_N.n0 76.833
R144 a_1191_21.n0 a_1191_21.t2 212.079
R145 a_1191_21.n1 a_1191_21.t3 212.079
R146 a_1191_21.n3 a_1191_21.t4 212.079
R147 a_1191_21.n2 a_1191_21.t5 212.079
R148 a_1191_21.t1 a_1191_21.n7 169.477
R149 a_1191_21.n0 a_1191_21.t8 139.779
R150 a_1191_21.n1 a_1191_21.t9 139.779
R151 a_1191_21.n3 a_1191_21.t7 139.779
R152 a_1191_21.n2 a_1191_21.t6 139.779
R153 a_1191_21.n7 a_1191_21.t0 123.36
R154 a_1191_21.n7 a_1191_21.n0 114.706
R155 a_1191_21.n6 a_1191_21.n4 96.723
R156 a_1191_21.n6 a_1191_21.n5 76
R157 a_1191_21.n3 a_1191_21.n2 61.345
R158 a_1191_21.n4 a_1191_21.n3 51.121
R159 a_1191_21.n7 a_1191_21.n6 25.295
R160 a_1191_21.n4 a_1191_21.n1 10.224
R161 a_803_297.n4 a_803_297.t7 225.591
R162 a_803_297.n1 a_803_297.t3 225.591
R163 a_803_297.n1 a_803_297.n0 154.573
R164 a_803_297.n5 a_803_297.n4 154.572
R165 a_803_297.n3 a_803_297.n2 110.761
R166 a_803_297.n3 a_803_297.n1 44.423
R167 a_803_297.n4 a_803_297.n3 44.423
R168 a_803_297.n0 a_803_297.t1 26.595
R169 a_803_297.n0 a_803_297.t2 26.595
R170 a_803_297.n2 a_803_297.t4 26.595
R171 a_803_297.n2 a_803_297.t0 26.595
R172 a_803_297.t6 a_803_297.n5 26.595
R173 a_803_297.n5 a_803_297.t5 26.595
R174 VPB.t12 VPB.t4 556.386
R175 VPB.t2 VPB.t8 556.386
R176 VPB.t11 VPB.t12 248.598
R177 VPB.t10 VPB.t11 248.598
R178 VPB.t9 VPB.t10 248.598
R179 VPB.t5 VPB.t9 248.598
R180 VPB.t6 VPB.t5 248.598
R181 VPB.t7 VPB.t6 248.598
R182 VPB.t8 VPB.t7 248.598
R183 VPB.t1 VPB.t2 248.598
R184 VPB.t0 VPB.t1 248.598
R185 VPB.t3 VPB.t0 248.598
R186 VPB.t14 VPB.t3 248.598
R187 VPB.t15 VPB.t14 248.598
R188 VPB.t16 VPB.t15 248.598
R189 VPB.t13 VPB.t16 248.598
R190 VPB VPB.t13 192.367
R191 a_27_297.n4 a_27_297.t2 225.591
R192 a_27_297.n2 a_27_297.t4 176.028
R193 a_27_297.n5 a_27_297.n4 154.572
R194 a_27_297.n2 a_27_297.n1 110.76
R195 a_27_297.n3 a_27_297.n0 90.234
R196 a_27_297.n3 a_27_297.n2 64.95
R197 a_27_297.n4 a_27_297.n3 64.95
R198 a_27_297.n0 a_27_297.t3 26.595
R199 a_27_297.n0 a_27_297.t5 26.595
R200 a_27_297.n1 a_27_297.t6 26.595
R201 a_27_297.n1 a_27_297.t7 26.595
R202 a_27_297.n5 a_27_297.t1 26.595
R203 a_27_297.t0 a_27_297.n5 26.595
R204 a_445_297.n5 a_445_297.n4 198.997
R205 a_445_297.n2 a_445_297.n0 198.996
R206 a_445_297.n2 a_445_297.n1 154.573
R207 a_445_297.n4 a_445_297.n3 154.573
R208 a_445_297.n4 a_445_297.n2 83.576
R209 a_445_297.n0 a_445_297.t4 26.595
R210 a_445_297.n0 a_445_297.t5 26.595
R211 a_445_297.n1 a_445_297.t6 26.595
R212 a_445_297.n1 a_445_297.t7 26.595
R213 a_445_297.n3 a_445_297.t2 26.595
R214 a_445_297.n3 a_445_297.t1 26.595
R215 a_445_297.n5 a_445_297.t0 26.595
R216 a_445_297.t3 a_445_297.n5 26.595
R217 A.n0 A.t0 212.079
R218 A.n2 A.t1 212.079
R219 A.n7 A.t2 212.079
R220 A.n5 A.t6 212.079
R221 A.n0 A.t4 139.779
R222 A.n2 A.t5 139.779
R223 A.n7 A.t3 139.779
R224 A.n5 A.t7 139.779
R225 A.n9 A.n6 96.723
R226 A.n4 A.n1 96.723
R227 A.n4 A.n3 76
R228 A.n9 A.n8 76
R229 A.n1 A.n0 21.909
R230 A.n6 A.n5 13.145
R231 A A.n4 11.58
R232 A.n3 A.n2 10.224
R233 A A.n9 9.142
R234 A.n8 A.n7 1.46
R235 VPWR.n6 VPWR.n5 176.855
R236 VPWR.n1 VPWR.n0 171.981
R237 VPWR.n2 VPWR.t0 162.553
R238 VPWR.n0 VPWR.t4 26.595
R239 VPWR.n0 VPWR.t3 26.595
R240 VPWR.n5 VPWR.t2 26.595
R241 VPWR.n5 VPWR.t1 26.595
R242 VPWR.n4 VPWR.n3 4.65
R243 VPWR.n2 VPWR.n1 4.107
R244 VPWR.n7 VPWR.n6 4.05
R245 VPWR.n4 VPWR.n2 0.135
R246 VPWR.n7 VPWR.n4 0.134
R247 VPWR VPWR.n7 0.126
R248 C.n0 C.t4 212.079
R249 C.n2 C.t5 212.079
R250 C.n5 C.t6 212.079
R251 C.n8 C.t7 212.079
R252 C.n0 C.t2 139.779
R253 C.n2 C.t0 139.779
R254 C.n5 C.t3 139.779
R255 C.n8 C.t1 139.779
R256 C.n4 C.n1 96.723
R257 C C.n9 94.895
R258 C.n4 C.n3 76
R259 C.n7 C.n6 76
R260 C.n1 C.n0 21.909
R261 C.n7 C.n4 20.723
R262 C.n9 C.n8 13.145
R263 C.n3 C.n2 10.224
R264 C C.n7 1.828
R265 C.n6 C.n5 1.46
C0 B Y 0.34fF
C1 VPWR VGND 0.18fF
C2 VPWR VPB 0.17fF
C3 C Y 0.33fF
C4 Y VGND 1.86fF
C5 A Y 0.25fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__nor4bb_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__nor4bb_1 A C_N D_N B Y VGND VPWR VNB VPB
X0 Y.t4 B.t0 VGND.t3 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 VGND.t2 a_27_410.t2 Y.t2 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 VGND.t4 C_N.t0 a_27_410.t0 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3 VGND.t1 A.t0 Y.t1 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 VPWR.t1 C_N.t1 a_27_410.t1 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 a_205_93.t1 D_N.t0 VGND.t5 VNB.t5 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 VPWR.t0 A.t1 a_573_297.t0 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 a_205_93.t0 D_N.t1 VPWR.t2 VPB.t5 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 a_477_297.t0 a_27_410.t3 a_393_297.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 a_573_297.t1 B.t1 a_477_297.t1 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 a_393_297.t1 a_205_93.t2 Y.t3 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 Y.t0 a_205_93.t3 VGND.t0 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
R0 B.n0 B.t1 241.534
R1 B.n0 B.t0 169.234
R2 B B.n0 87.054
R3 VGND.n5 VGND.t0 190.315
R4 VGND.n10 VGND.n9 135.794
R5 VGND.n2 VGND.t1 107.734
R6 VGND.n1 VGND.n0 107.627
R7 VGND.n9 VGND.t4 44.285
R8 VGND.n9 VGND.t5 38.571
R9 VGND.n0 VGND.t3 30.461
R10 VGND.n0 VGND.t2 30.461
R11 VGND.n11 VGND.n10 7.911
R12 VGND.n4 VGND.n3 4.65
R13 VGND.n6 VGND.n5 4.65
R14 VGND.n8 VGND.n7 4.65
R15 VGND.n2 VGND.n1 3.776
R16 VGND.n4 VGND.n2 0.258
R17 VGND.n11 VGND.n8 0.132
R18 VGND VGND.n11 0.127
R19 VGND.n6 VGND.n4 0.119
R20 VGND.n8 VGND.n6 0.119
R21 Y.n1 Y.t3 423.446
R22 Y.n1 Y.n0 102.74
R23 Y.n3 Y.n2 92.5
R24 Y.n3 Y.n1 73.656
R25 Y.n2 Y.t1 24.923
R26 Y.n2 Y.t4 24.923
R27 Y.n0 Y.t2 24.923
R28 Y.n0 Y.t0 24.923
R29 Y Y.n3 4.48
R30 VNB VNB.t4 12650
R31 VNB.t5 VNB.t0 5321.88
R32 VNB.t4 VNB.t5 2847.06
R33 VNB.t2 VNB.t3 2320.88
R34 VNB.t3 VNB.t1 2030.77
R35 VNB.t0 VNB.t2 2030.77
R36 a_27_410.n1 a_27_410.t1 371.328
R37 a_27_410.n1 a_27_410.n0 321.62
R38 a_27_410.n0 a_27_410.t3 241.534
R39 a_27_410.t0 a_27_410.n1 219.632
R40 a_27_410.n0 a_27_410.t2 169.234
R41 C_N.n0 C_N.t1 329.901
R42 C_N.n0 C_N.t0 132.281
R43 C_N.n1 C_N.n0 76
R44 C_N.n1 C_N 10.422
R45 C_N C_N.n1 2.011
R46 A.n0 A.t1 235.819
R47 A.n0 A.t0 163.519
R48 A A.n0 77.171
R49 VPWR.n0 VPWR.t2 327.591
R50 VPWR.n1 VPWR.n0 311.239
R51 VPWR.n1 VPWR.t0 195.388
R52 VPWR.n0 VPWR.t1 63.321
R53 VPWR VPWR.n1 0.141
R54 VPB.t5 VPB.t2 553.426
R55 VPB.t4 VPB.t5 287.071
R56 VPB.t0 VPB.t3 284.112
R57 VPB.t3 VPB.t1 248.598
R58 VPB.t2 VPB.t0 248.598
R59 VPB VPB.t4 189.408
R60 D_N.n0 D_N.t1 142.993
R61 D_N.n0 D_N.t0 126.926
R62 D_N D_N.n0 78.427
R63 a_205_93.n2 a_205_93.n1 344.005
R64 a_205_93.n0 a_205_93.t2 227.985
R65 a_205_93.n1 a_205_93.t1 175.707
R66 a_205_93.n0 a_205_93.t3 155.685
R67 a_205_93.n1 a_205_93.n0 76
R68 a_205_93.n3 a_205_93.n2 54.078
R69 a_205_93.n2 a_205_93.t0 33.487
R70 a_573_297.t0 a_573_297.t1 53.19
R71 a_393_297.t0 a_393_297.t1 53.19
R72 a_477_297.t0 a_477_297.t1 65.01
C0 Y VGND 0.31fF
C1 B VPWR 0.13fF
C2 C_N D_N 0.11fF
C3 B A 0.15fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__nor4bb_2.ext - technology: sky130A

.subckt sky130_fd_sc_hd__nor4bb_2 D_N C_N A Y B VGND VPWR VNB VPB
X0 Y.t1 a_27_410.t2 a_336_297.t1 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 Y.t4 A.t0 VGND.t3 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 a_336_297.t2 a_201_93.t2 a_418_297.t1 VPB.t8 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 Y.t8 a_201_93.t3 VGND.t8 VNB.t8 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 Y.t3 a_27_410.t3 VGND.t1 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 Y.t6 B.t0 VGND.t6 VNB.t6 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 a_418_297.t0 a_201_93.t4 a_336_297.t3 VPB.t9 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 VGND.t4 D_N.t0 a_27_410.t0 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 VPWR.t3 D_N.t1 a_27_410.t1 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9 VGND.t2 A.t1 Y.t5 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 VGND.t7 B.t1 Y.t7 VNB.t7 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 a_776_297.t3 A.t2 VPWR.t1 VPB.t5 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 a_201_93.t0 C_N.t0 VPWR.t2 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13 a_201_93.t1 C_N.t1 VGND.t5 VNB.t5 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14 VPWR.t0 A.t3 a_776_297.t2 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 a_776_297.t1 B.t2 a_418_297.t2 VPB.t6 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16 VGND.t9 a_201_93.t5 Y.t9 VNB.t9 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X17 a_336_297.t0 a_27_410.t4 Y.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X18 a_418_297.t3 B.t3 a_776_297.t0 VPB.t7 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X19 VGND.t0 a_27_410.t5 Y.t2 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
R0 a_27_410.n3 a_27_410.t1 371.574
R1 a_27_410.n3 a_27_410.n2 255.879
R2 a_27_410.t0 a_27_410.n3 220.623
R3 a_27_410.n0 a_27_410.t4 212.079
R4 a_27_410.n1 a_27_410.t2 212.079
R5 a_27_410.n0 a_27_410.t5 139.779
R6 a_27_410.n1 a_27_410.t3 139.779
R7 a_27_410.n2 a_27_410.n0 26.842
R8 a_27_410.n2 a_27_410.n1 23.465
R9 a_336_297.n1 a_336_297.t3 594.398
R10 a_336_297.t0 a_336_297.n1 574.181
R11 a_336_297.n1 a_336_297.n0 292.5
R12 a_336_297.n0 a_336_297.t1 26.595
R13 a_336_297.n0 a_336_297.t2 26.595
R14 Y Y.n0 307.269
R15 Y.n6 Y.n4 88.89
R16 Y.n3 Y.n1 88.89
R17 Y.n6 Y.n5 52.624
R18 Y.n3 Y.n2 52.624
R19 Y.n0 Y.t0 26.595
R20 Y.n0 Y.t1 26.595
R21 Y.n4 Y.t5 24.923
R22 Y.n4 Y.t4 24.923
R23 Y.n5 Y.t7 24.923
R24 Y.n5 Y.t6 24.923
R25 Y.n1 Y.t9 24.923
R26 Y.n1 Y.t8 24.923
R27 Y.n2 Y.t2 24.923
R28 Y.n2 Y.t3 24.923
R29 Y.n7 Y.n3 24.533
R30 Y.n7 Y.n6 20.266
R31  Y.n7 19.2
R32  Y 14.299
R33 VPB.t3 VPB.t9 627.414
R34 VPB.t0 VPB.t7 568.224
R35 VPB.t2 VPB.t3 287.071
R36 VPB.t4 VPB.t5 248.598
R37 VPB.t6 VPB.t4 248.598
R38 VPB.t7 VPB.t6 248.598
R39 VPB.t1 VPB.t0 248.598
R40 VPB.t8 VPB.t1 248.598
R41 VPB.t9 VPB.t8 248.598
R42 VPB VPB.t2 192.367
R43 A.n0 A.t2 212.079
R44 A.n1 A.t3 212.079
R45 A.n0 A.t1 139.779
R46 A.n1 A.t0 139.779
R47 A A.n2 81.76
R48 A.n2 A.n1 32.133
R49 A.n2 A.n0 29.212
R50 VGND.n10 VGND.t0 170.961
R51 VGND.n7 VGND.t6 165.357
R52 VGND.n21 VGND.t8 147.319
R53 VGND.n26 VGND.n25 135.794
R54 VGND.n2 VGND.n1 115.464
R55 VGND.n16 VGND.n15 115.464
R56 VGND.n0 VGND.t2 108.731
R57 VGND.n25 VGND.t5 38.571
R58 VGND.n25 VGND.t4 38.571
R59 VGND.n1 VGND.t3 24.923
R60 VGND.n1 VGND.t7 24.923
R61 VGND.n15 VGND.t1 24.923
R62 VGND.n15 VGND.t9 24.923
R63 VGND.n17 VGND.n16 8.658
R64 VGND.n27 VGND.n26 6.405
R65 VGND.n4 VGND.n3 4.65
R66 VGND.n6 VGND.n5 4.65
R67 VGND.n9 VGND.n8 4.65
R68 VGND.n12 VGND.n11 4.65
R69 VGND.n14 VGND.n13 4.65
R70 VGND.n18 VGND.n17 4.65
R71 VGND.n20 VGND.n19 4.65
R72 VGND.n22 VGND.n21 4.65
R73 VGND.n24 VGND.n23 4.65
R74 VGND.n3 VGND.n2 2.635
R75 VGND.n8 VGND.n7 2.3
R76 VGND.n4 VGND.n0 0.767
R77 VGND.n11 VGND.n10 0.7
R78 VGND.n27 VGND.n24 0.132
R79 VGND VGND.n27 0.129
R80 VGND.n6 VGND.n4 0.119
R81 VGND.n9 VGND.n6 0.119
R82 VGND.n12 VGND.n9 0.119
R83 VGND.n14 VGND.n12 0.119
R84 VGND.n18 VGND.n14 0.119
R85 VGND.n20 VGND.n18 0.119
R86 VGND.n22 VGND.n20 0.119
R87 VGND.n24 VGND.n22 0.119
R88 VNB VNB.t4 12682.4
R89 VNB.t5 VNB.t8 6129.28
R90 VNB.t0 VNB.t6 4641.76
R91 VNB.t4 VNB.t5 2717.65
R92 VNB.t3 VNB.t2 2030.77
R93 VNB.t7 VNB.t3 2030.77
R94 VNB.t6 VNB.t7 2030.77
R95 VNB.t1 VNB.t0 2030.77
R96 VNB.t9 VNB.t1 2030.77
R97 VNB.t8 VNB.t9 2030.77
R98 a_201_93.t0 a_201_93.n3 398.797
R99 a_201_93.n0 a_201_93.t2 212.079
R100 a_201_93.n1 a_201_93.t4 212.079
R101 a_201_93.n3 a_201_93.t1 171.718
R102 a_201_93.n0 a_201_93.t5 139.779
R103 a_201_93.n1 a_201_93.t3 139.779
R104 a_201_93.n3 a_201_93.n2 72.207
R105 a_201_93.n2 a_201_93.n0 44.385
R106 a_201_93.n2 a_201_93.n1 12.82
R107 a_418_297.n1 a_418_297.n0 600.15
R108 a_418_297.n0 a_418_297.t2 26.595
R109 a_418_297.n0 a_418_297.t3 26.595
R110 a_418_297.t1 a_418_297.n1 26.595
R111 a_418_297.n1 a_418_297.t0 26.595
R112 B.n0 B.t2 212.079
R113 B.n1 B.t3 212.079
R114 B.n0 B.t1 139.779
R115 B.n1 B.t0 139.779
R116 B B.n2 87.2
R117 B.n2 B.n1 32.863
R118 B.n2 B.n0 28.481
R119 D_N.n0 D_N.t1 329.901
R120 D_N.n0 D_N.t0 132.281
R121 D_N.n1 D_N.n0 76
R122  D_N.n1 10.276
R123 D_N.n1 D_N 1.983
R124 VPWR.n1 VPWR.t2 327.591
R125 VPWR.n2 VPWR.n1 311.239
R126 VPWR.n2 VPWR.n0 181.605
R127 VPWR.n1 VPWR.t3 63.321
R128 VPWR.n0 VPWR.t1 26.595
R129 VPWR.n0 VPWR.t0 26.595
R130 VPWR VPWR.n2 0.143
R131 a_776_297.n0 a_776_297.t0 574.021
R132 a_776_297.n0 a_776_297.t3 199.067
R133 a_776_297.n1 a_776_297.n0 89.753
R134 a_776_297.n1 a_776_297.t2 26.595
R135 a_776_297.t1 a_776_297.n1 26.595
R136 C_N.n0 C_N.t0 141.945
R137 C_N.n0 C_N.t1 125.878
R138 C_N C_N.n0 78.47
C0 VPWR VGND 0.13fF
C1 B Y 0.21fF
C2 D_N C_N 0.11fF
C3 Y VGND 0.99fF
C4 VPB VPWR 0.12fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__nor4bb_4.ext - technology: sky130A

.subckt sky130_fd_sc_hd__nor4bb_4 D_N Y A B C_N VGND VPWR VNB VPB
X0 Y.t9 B.t0 VGND.t9 VNB.t9 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 a_729_297.t7 a_27_297.t2 a_311_297.t7 VPB.t14 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 Y.t8 B.t1 VGND.t8 VNB.t8 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 Y.t4 A.t0 VGND.t4 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 a_197_47.t0 D_N.t0 VPWR.t0 VPB.t17 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 a_311_297.t6 a_27_297.t3 a_729_297.t6 VPB.t13 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 Y.t5 A.t1 VGND.t5 VNB.t5 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 a_729_297.t3 B.t2 a_1087_297.t7 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 VGND.t10 a_197_47.t2 Y.t10 VNB.t10 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 VGND.t11 a_197_47.t3 Y.t11 VNB.t11 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 a_729_297.t5 a_27_297.t4 a_311_297.t5 VPB.t12 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 a_1087_297.t6 B.t3 a_729_297.t2 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 VGND.t0 a_27_297.t5 Y.t0 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 a_197_47.t1 D_N.t1 VGND.t15 VNB.t15 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14 VGND.t1 a_27_297.t6 Y.t1 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X15 VGND.t14 C_N.t0 a_27_297.t1 VNB.t14 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X16 a_729_297.t1 B.t4 a_1087_297.t5 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17 VGND.t16 A.t2 Y.t18 VNB.t16 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X18 VGND.t17 A.t3 Y.t19 VNB.t17 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X19 a_1087_297.t3 A.t4 VPWR.t4 VPB.t15 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X20 Y.t2 a_27_297.t7 VGND.t2 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X21 Y.t3 a_27_297.t8 VGND.t3 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X22 VPWR.t3 A.t5 a_1087_297.t2 VPB.t16 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X23 VPWR.t5 C_N.t1 a_27_297.t0 VPB.t8 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X24 a_311_297.t0 a_197_47.t4 Y.t12 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X25 Y.t13 a_197_47.t5 a_311_297.t1 VPB.t5 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X26 a_1087_297.t1 A.t6 VPWR.t2 VPB.t9 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X27 VPWR.t1 A.t7 a_1087_297.t0 VPB.t10 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X28 a_311_297.t2 a_197_47.t6 Y.t14 VPB.t6 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X29 a_1087_297.t4 B.t5 a_729_297.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X30 VGND.t7 B.t6 Y.t7 VNB.t7 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X31 Y.t15 a_197_47.t7 a_311_297.t3 VPB.t7 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X32 VGND.t6 B.t7 Y.t6 VNB.t6 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X33 Y.t16 a_197_47.t8 VGND.t12 VNB.t12 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X34 a_311_297.t4 a_27_297.t9 a_729_297.t4 VPB.t11 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X35 Y.t17 a_197_47.t9 VGND.t13 VNB.t13 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
R0 B.n0 B.t5 212.079
R1 B.n2 B.t2 212.079
R2 B.n5 B.t3 212.079
R3 B.n8 B.t4 212.079
R4 B.n0 B.t7 139.779
R5 B.n2 B.t1 139.779
R6 B.n5 B.t6 139.779
R7 B.n8 B.t0 139.779
R8 B.n4 B.n1 96.723
R9 B B.n9 88.19
R10 B.n4 B.n3 76
R11 B.n7 B.n6 76
R12 B.n9 B.n8 21.909
R13 B.n7 B.n4 20.723
R14 B.n1 B.n0 13.145
R15 B.n6 B.n5 10.224
R16 B B.n7 8.533
R17 B.n3 B.n2 1.46
R18 VGND.n45 VGND.t12 193.925
R19 VGND.n2 VGND.n1 115.464
R20 VGND.n8 VGND.n7 115.464
R21 VGND.n14 VGND.n13 115.464
R22 VGND.n28 VGND.n27 115.464
R23 VGND.n34 VGND.n33 115.464
R24 VGND.n40 VGND.n39 115.464
R25 VGND.n51 VGND.n50 115.464
R26 VGND.n0 VGND.t17 108.053
R27 VGND.n20 VGND.n19 92.5
R28 VGND.n22 VGND.n21 92.5
R29 VGND.n19 VGND.t9 24.923
R30 VGND.n21 VGND.t1 24.923
R31 VGND.n1 VGND.t5 24.923
R32 VGND.n1 VGND.t16 24.923
R33 VGND.n7 VGND.t4 24.923
R34 VGND.n7 VGND.t6 24.923
R35 VGND.n13 VGND.t8 24.923
R36 VGND.n13 VGND.t7 24.923
R37 VGND.n27 VGND.t3 24.923
R38 VGND.n27 VGND.t0 24.923
R39 VGND.n33 VGND.t2 24.923
R40 VGND.n33 VGND.t11 24.923
R41 VGND.n39 VGND.t13 24.923
R42 VGND.n39 VGND.t10 24.923
R43 VGND.n50 VGND.t15 24.923
R44 VGND.n50 VGND.t14 24.923
R45 VGND.n15 VGND.n14 14.305
R46 VGND.n29 VGND.n28 12.8
R47 VGND.n9 VGND.n8 8.282
R48 VGND.n35 VGND.n34 6.776
R49 VGND.n23 VGND.n20 5.4
R50 VGND.n46 VGND.n45 5.27
R51 VGND.n23 VGND.n22 5
R52 VGND.n52 VGND.n51 4.899
R53 VGND.n4 VGND.n3 4.65
R54 VGND.n6 VGND.n5 4.65
R55 VGND.n10 VGND.n9 4.65
R56 VGND.n12 VGND.n11 4.65
R57 VGND.n16 VGND.n15 4.65
R58 VGND.n18 VGND.n17 4.65
R59 VGND.n24 VGND.n23 4.65
R60 VGND.n26 VGND.n25 4.65
R61 VGND.n30 VGND.n29 4.65
R62 VGND.n32 VGND.n31 4.65
R63 VGND.n36 VGND.n35 4.65
R64 VGND.n38 VGND.n37 4.65
R65 VGND.n42 VGND.n41 4.65
R66 VGND.n44 VGND.n43 4.65
R67 VGND.n47 VGND.n46 4.65
R68 VGND.n49 VGND.n48 4.65
R69 VGND.n3 VGND.n2 2.258
R70 VGND.n4 VGND.n0 0.774
R71 VGND.n41 VGND.n40 0.752
R72 VGND.n52 VGND.n49 0.132
R73 VGND VGND.n52 0.127
R74 VGND.n6 VGND.n4 0.119
R75 VGND.n10 VGND.n6 0.119
R76 VGND.n12 VGND.n10 0.119
R77 VGND.n16 VGND.n12 0.119
R78 VGND.n18 VGND.n16 0.119
R79 VGND.n24 VGND.n18 0.119
R80 VGND.n26 VGND.n24 0.119
R81 VGND.n30 VGND.n26 0.119
R82 VGND.n32 VGND.n30 0.119
R83 VGND.n36 VGND.n32 0.119
R84 VGND.n38 VGND.n36 0.119
R85 VGND.n42 VGND.n38 0.119
R86 VGND.n44 VGND.n42 0.119
R87 VGND.n47 VGND.n44 0.119
R88 VGND.n49 VGND.n47 0.119
R89 Y Y.n17 327.81
R90 Y.n16 Y.n15 292.5
R91 Y.n13 Y.n12 100.623
R92 Y.n2 Y.n0 88.89
R93 Y.n8 Y.n6 73.244
R94 Y.n2 Y.n1 52.624
R95 Y.n4 Y.n3 52.624
R96 Y.n6 Y.n5 52.624
R97 Y.n8 Y.n7 52.624
R98 Y.n10 Y.n9 52.624
R99 Y.n13 Y.n11 49.285
R100 Y.n16 Y.n14 45.462
R101 Y.n14 Y.n10 36.622
R102 Y.n4 Y.n2 36.266
R103 Y.n6 Y.n4 36.266
R104 Y.n10 Y.n8 36.266
R105 Y.n17 Y.t14 26.595
R106 Y.n17 Y.t15 26.595
R107 Y.n15 Y.t12 26.595
R108 Y.n15 Y.t13 26.595
R109 Y.n11 Y.t11 24.923
R110 Y.n11 Y.t17 24.923
R111 Y.n12 Y.t10 24.923
R112 Y.n12 Y.t16 24.923
R113 Y.n0 Y.t19 24.923
R114 Y.n0 Y.t5 24.923
R115 Y.n1 Y.t18 24.923
R116 Y.n1 Y.t4 24.923
R117 Y.n3 Y.t6 24.923
R118 Y.n3 Y.t8 24.923
R119 Y.n5 Y.t7 24.923
R120 Y.n5 Y.t9 24.923
R121 Y.n7 Y.t1 24.923
R122 Y.n7 Y.t3 24.923
R123 Y.n9 Y.t0 24.923
R124 Y.n9 Y.t2 24.923
R125 Y.n14 Y.n13 11.377
R126 Y Y.n16 1.765
R127 VNB VNB.t14 6150.61
R128 VNB.t15 VNB.t12 4738.46
R129 VNB.t1 VNB.t9 4545.05
R130 VNB.t5 VNB.t17 2030.77
R131 VNB.t16 VNB.t5 2030.77
R132 VNB.t4 VNB.t16 2030.77
R133 VNB.t6 VNB.t4 2030.77
R134 VNB.t8 VNB.t6 2030.77
R135 VNB.t7 VNB.t8 2030.77
R136 VNB.t9 VNB.t7 2030.77
R137 VNB.t3 VNB.t1 2030.77
R138 VNB.t0 VNB.t3 2030.77
R139 VNB.t2 VNB.t0 2030.77
R140 VNB.t11 VNB.t2 2030.77
R141 VNB.t13 VNB.t11 2030.77
R142 VNB.t10 VNB.t13 2030.77
R143 VNB.t12 VNB.t10 2030.77
R144 VNB.t14 VNB.t15 2030.77
R145 a_27_297.n11 a_27_297.n10 263.527
R146 a_27_297.n0 a_27_297.t9 212.079
R147 a_27_297.n2 a_27_297.t2 212.079
R148 a_27_297.n5 a_27_297.t3 212.079
R149 a_27_297.n8 a_27_297.t4 212.079
R150 a_27_297.n11 a_27_297.t1 156.49
R151 a_27_297.n0 a_27_297.t6 139.779
R152 a_27_297.n2 a_27_297.t8 139.779
R153 a_27_297.n5 a_27_297.t5 139.779
R154 a_27_297.n8 a_27_297.t7 139.779
R155 a_27_297.t0 a_27_297.n11 136.044
R156 a_27_297.n4 a_27_297.n1 96.723
R157 a_27_297.n10 a_27_297.n9 76
R158 a_27_297.n4 a_27_297.n3 76
R159 a_27_297.n7 a_27_297.n6 76
R160 a_27_297.n9 a_27_297.n8 21.909
R161 a_27_297.n7 a_27_297.n4 20.723
R162 a_27_297.n10 a_27_297.n7 20.723
R163 a_27_297.n1 a_27_297.n0 13.145
R164 a_27_297.n6 a_27_297.n5 10.224
R165 a_27_297.n3 a_27_297.n2 1.46
R166 a_311_297.n3 a_311_297.t3 574.181
R167 a_311_297.n3 a_311_297.n2 292.5
R168 a_311_297.n5 a_311_297.n4 292.5
R169 a_311_297.n1 a_311_297.t4 224.711
R170 a_311_297.n1 a_311_297.n0 154.573
R171 a_311_297.n4 a_311_297.n1 49.859
R172 a_311_297.n4 a_311_297.n3 43.008
R173 a_311_297.n2 a_311_297.t1 26.595
R174 a_311_297.n2 a_311_297.t2 26.595
R175 a_311_297.n0 a_311_297.t7 26.595
R176 a_311_297.n0 a_311_297.t6 26.595
R177 a_311_297.n5 a_311_297.t5 26.595
R178 a_311_297.t0 a_311_297.n5 26.595
R179 a_729_297.n5 a_729_297.n4 200.554
R180 a_729_297.n2 a_729_297.n0 198.996
R181 a_729_297.n2 a_729_297.n1 154.573
R182 a_729_297.n4 a_729_297.n3 154.573
R183 a_729_297.n4 a_729_297.n2 83.576
R184 a_729_297.n0 a_729_297.t0 26.595
R185 a_729_297.n0 a_729_297.t3 26.595
R186 a_729_297.n1 a_729_297.t2 26.595
R187 a_729_297.n1 a_729_297.t1 26.595
R188 a_729_297.n3 a_729_297.t4 26.595
R189 a_729_297.n3 a_729_297.t7 26.595
R190 a_729_297.t6 a_729_297.n5 26.595
R191 a_729_297.n5 a_729_297.t5 26.595
R192 VPB.t17 VPB.t7 580.062
R193 VPB.t11 VPB.t1 556.386
R194 VPB.t16 VPB.t15 248.598
R195 VPB.t9 VPB.t16 248.598
R196 VPB.t10 VPB.t9 248.598
R197 VPB.t0 VPB.t10 248.598
R198 VPB.t3 VPB.t0 248.598
R199 VPB.t2 VPB.t3 248.598
R200 VPB.t1 VPB.t2 248.598
R201 VPB.t14 VPB.t11 248.598
R202 VPB.t13 VPB.t14 248.598
R203 VPB.t12 VPB.t13 248.598
R204 VPB.t4 VPB.t12 248.598
R205 VPB.t5 VPB.t4 248.598
R206 VPB.t6 VPB.t5 248.598
R207 VPB.t7 VPB.t6 248.598
R208 VPB.t8 VPB.t17 248.598
R209 VPB VPB.t8 201.246
R210 A.n0 A.t4 212.079
R211 A.n2 A.t5 212.079
R212 A.n7 A.t6 212.079
R213 A.n5 A.t7 212.079
R214 A.n0 A.t3 139.779
R215 A.n2 A.t1 139.779
R216 A.n7 A.t2 139.779
R217 A.n5 A.t0 139.779
R218 A.n9 A.n6 96.723
R219 A.n4 A.n1 96.723
R220 A.n4 A.n3 76
R221 A.n9 A.n8 76
R222 A.n6 A.n5 21.909
R223 A A.n4 19.504
R224 A.n1 A.n0 13.145
R225 A.n8 A.n7 10.224
R226 A.n3 A.n2 1.46
R227 A A.n9 1.219
R228 D_N.n0 D_N.t0 229.752
R229 D_N.n0 D_N.t1 157.452
R230 D_N D_N.n0 78.07
R231 VPWR.n33 VPWR.n32 308.79
R232 VPWR.n3 VPWR.n2 175.611
R233 VPWR.n1 VPWR.n0 171.981
R234 VPWR.n2 VPWR.t4 26.595
R235 VPWR.n2 VPWR.t3 26.595
R236 VPWR.n0 VPWR.t2 26.595
R237 VPWR.n0 VPWR.t1 26.595
R238 VPWR.n32 VPWR.t0 26.595
R239 VPWR.n32 VPWR.t5 26.595
R240 VPWR.n5 VPWR.n4 4.65
R241 VPWR.n7 VPWR.n6 4.65
R242 VPWR.n9 VPWR.n8 4.65
R243 VPWR.n11 VPWR.n10 4.65
R244 VPWR.n13 VPWR.n12 4.65
R245 VPWR.n15 VPWR.n14 4.65
R246 VPWR.n17 VPWR.n16 4.65
R247 VPWR.n19 VPWR.n18 4.65
R248 VPWR.n21 VPWR.n20 4.65
R249 VPWR.n23 VPWR.n22 4.65
R250 VPWR.n25 VPWR.n24 4.65
R251 VPWR.n27 VPWR.n26 4.65
R252 VPWR.n29 VPWR.n28 4.65
R253 VPWR.n31 VPWR.n30 4.65
R254 VPWR.n34 VPWR.n33 3.966
R255 VPWR.n3 VPWR.n1 3.784
R256 VPWR.n5 VPWR.n3 0.233
R257 VPWR.n34 VPWR.n31 0.137
R258 VPWR VPWR.n34 0.122
R259 VPWR.n7 VPWR.n5 0.119
R260 VPWR.n9 VPWR.n7 0.119
R261 VPWR.n11 VPWR.n9 0.119
R262 VPWR.n13 VPWR.n11 0.119
R263 VPWR.n15 VPWR.n13 0.119
R264 VPWR.n17 VPWR.n15 0.119
R265 VPWR.n19 VPWR.n17 0.119
R266 VPWR.n21 VPWR.n19 0.119
R267 VPWR.n23 VPWR.n21 0.119
R268 VPWR.n25 VPWR.n23 0.119
R269 VPWR.n27 VPWR.n25 0.119
R270 VPWR.n29 VPWR.n27 0.119
R271 VPWR.n31 VPWR.n29 0.119
R272 a_197_47.t0 a_197_47.n7 603.514
R273 a_197_47.n0 a_197_47.t4 212.079
R274 a_197_47.n1 a_197_47.t5 212.079
R275 a_197_47.n2 a_197_47.t6 212.079
R276 a_197_47.n4 a_197_47.t7 212.079
R277 a_197_47.n0 a_197_47.t3 139.779
R278 a_197_47.n1 a_197_47.t9 139.779
R279 a_197_47.n2 a_197_47.t2 139.779
R280 a_197_47.n4 a_197_47.t8 139.779
R281 a_197_47.n7 a_197_47.t1 124.898
R282 a_197_47.n6 a_197_47.n5 76
R283 a_197_47.n1 a_197_47.n0 61.345
R284 a_197_47.n6 a_197_47.n3 59.578
R285 a_197_47.n7 a_197_47.n6 33.882
R286 a_197_47.n3 a_197_47.n1 29.505
R287 a_197_47.n3 a_197_47.n2 20.989
R288 a_197_47.n5 a_197_47.n4 16.066
R289 a_1087_297.n2 a_1087_297.t5 224.108
R290 a_1087_297.t3 a_1087_297.n5 179.121
R291 a_1087_297.n2 a_1087_297.n1 154.573
R292 a_1087_297.n5 a_1087_297.n4 110.76
R293 a_1087_297.n3 a_1087_297.n0 90.234
R294 a_1087_297.n3 a_1087_297.n2 64.95
R295 a_1087_297.n5 a_1087_297.n3 64.95
R296 a_1087_297.n0 a_1087_297.t0 26.595
R297 a_1087_297.n0 a_1087_297.t4 26.595
R298 a_1087_297.n1 a_1087_297.t7 26.595
R299 a_1087_297.n1 a_1087_297.t6 26.595
R300 a_1087_297.n4 a_1087_297.t2 26.595
R301 a_1087_297.n4 a_1087_297.t1 26.595
R302 C_N.n0 C_N.t1 231.014
R303 C_N.n0 C_N.t0 158.714
R304 C_N C_N.n0 81.737
C0 VPWR VGND 0.19fF
C1 B Y 0.36fF
C2 Y VGND 1.87fF
C3 A Y 0.24fF
C4 VPB VPWR 0.17fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__o2bb2a_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__o2bb2a_1 A1_N X A2_N B2 B1 VPWR VGND VNB VPB
X0 a_206_369.t2 A1_N.t0 VPWR.t4 VPB.t5 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1 a_206_369.t0 A2_N.t0 a_205_47.t0 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 VGND.t0 B2.t0 a_489_47.t0 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3 a_585_369.t0 B2.t1 a_76_199.t0 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 a_489_47.t1 a_206_369.t3 a_76_199.t1 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 a_489_47.t2 B1.t0 VGND.t2 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 VPWR.t1 A2_N.t1 a_206_369.t1 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7 a_76_199.t2 a_206_369.t4 VPWR.t3 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 a_205_47.t1 A1_N.t1 VGND.t3 VNB.t5 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9 VPWR.t2 a_76_199.t3 X.t1 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 VPWR.t0 B1.t1 a_585_369.t1 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11 VGND.t1 a_76_199.t4 X.t0 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
R0 A1_N.n0 A1_N.t0 264.028
R1 A1_N.n0 A1_N.t1 206.188
R2 A1_N A1_N.n0 79.52
R3 VPWR.n2 VPWR.t0 384.491
R4 VPWR.n8 VPWR.n7 349.688
R5 VPWR.n1 VPWR.n0 292.5
R6 VPWR.n0 VPWR.t3 135.266
R7 VPWR.n0 VPWR.t1 118.547
R8 VPWR.n7 VPWR.t4 96.154
R9 VPWR.n7 VPWR.t2 32.743
R10 VPWR.n2 VPWR.n1 7.581
R11 VPWR.n4 VPWR.n3 4.65
R12 VPWR.n6 VPWR.n5 4.65
R13 VPWR.n9 VPWR.n8 3.932
R14 VPWR.n4 VPWR.n2 0.144
R15 VPWR.n9 VPWR.n6 0.137
R16 VPWR VPWR.n9 0.121
R17 VPWR.n6 VPWR.n4 0.119
R18 a_206_369.n2 a_206_369.n0 495.257
R19 a_206_369.n1 a_206_369.t3 292.413
R20 a_206_369.t0 a_206_369.n2 212.915
R21 a_206_369.n2 a_206_369.n1 140.996
R22 a_206_369.n1 a_206_369.t4 120.429
R23 a_206_369.n0 a_206_369.t1 93.809
R24 a_206_369.n0 a_206_369.t2 93.809
R25 VPB.t2 VPB.t0 517.912
R26 VPB.t5 VPB.t2 325.545
R27 VPB.t3 VPB.t5 287.071
R28 VPB.t0 VPB.t4 278.193
R29 VPB.t4 VPB.t1 213.084
R30 VPB VPB.t3 189.408
R31 A2_N.n0 A2_N.t1 334.297
R32 A2_N.n0 A2_N.t0 131.857
R33 A2_N A2_N.n0 114.921
R34 a_205_47.t0 a_205_47.t1 90
R35 VNB.t4 VNB.t0 6179.41
R36 VNB VNB.t2 6053.91
R37 VNB.t5 VNB.t4 3008.82
R38 VNB.t1 VNB.t3 2717.65
R39 VNB.t0 VNB.t1 2717.65
R40 VNB.t2 VNB.t5 2279.52
R41 B2.n0 B2.t1 264.028
R42 B2.n0 B2.t0 206.188
R43 B2 B2.n0 95.017
R44 a_489_47.n0 a_489_47.t2 291.038
R45 a_489_47.t0 a_489_47.n0 38.571
R46 a_489_47.n0 a_489_47.t1 38.571
R47 VGND.n2 VGND.n1 130.241
R48 VGND.n2 VGND.n0 120.386
R49 VGND.n1 VGND.t3 48.571
R50 VGND.n0 VGND.t2 38.571
R51 VGND.n0 VGND.t0 38.571
R52 VGND.n1 VGND.t1 33.077
R53 VGND VGND.n2 0.145
R54 a_76_199.n2 a_76_199.n1 295.549
R55 a_76_199.n1 a_76_199.n0 243.151
R56 a_76_199.n0 a_76_199.t3 241.534
R57 a_76_199.n1 a_76_199.t1 211.49
R58 a_76_199.n0 a_76_199.t4 169.234
R59 a_76_199.t0 a_76_199.n2 86.773
R60 a_76_199.n2 a_76_199.t2 63.321
R61 a_585_369.t0 a_585_369.t1 98.5
R62 B1.n0 B1.t1 252.648
R63 B1.n0 B1.t0 194.808
R64 B1.n1 B1.n0 76
R65  B1.n1 10.573
R66 B1.n1 B1 2.04
R67 X.n0 X.t0 175.311
R68 X.n0 X.t1 172.965
R69 X X.n0 4.065
C0 B2 B1 0.18fF
C1 X VGND 0.10fF
C2 VPWR B2 0.14fF
C3 A1_N A2_N 0.11fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__o2bb2a_2.ext - technology: sky130A

.subckt sky130_fd_sc_hd__o2bb2a_2 A1_N X A2_N B2 B1 VGND VPWR VNB VPB
X0 a_294_47.t1 A1_N.t0 VGND.t2 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1 VPWR.t2 A2_N.t0 a_295_369.t0 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X2 VPWR.t5 B1.t0 a_665_369.t0 VPB.t6 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X3 VGND.t4 a_84_21.t3 X.t3 VNB.t6 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 X.t2 a_84_21.t4 VGND.t1 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 a_581_47.t2 a_295_369.t3 a_84_21.t2 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 VPWR.t0 a_84_21.t5 X.t1 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 a_665_369.t1 B2.t0 a_84_21.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X8 VGND.t0 B2.t1 a_581_47.t0 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9 a_295_369.t1 A2_N.t1 a_294_47.t0 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10 X.t0 a_84_21.t6 VPWR.t1 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 a_84_21.t1 a_295_369.t4 VPWR.t4 VPB.t5 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X12 a_295_369.t2 A1_N.t1 VPWR.t3 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X13 a_581_47.t1 B1.t1 VGND.t3 VNB.t5 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
R0 A1_N.n0 A1_N.t1 299.374
R1 A1_N.n0 A1_N.t0 206.188
R2 A1_N A1_N.n0 80.8
R3 VGND.n2 VGND.n1 125.629
R4 VGND.n3 VGND.n0 120.377
R5 VGND.n6 VGND.t1 104.879
R6 VGND.n1 VGND.t2 48.571
R7 VGND.n0 VGND.t3 38.571
R8 VGND.n0 VGND.t0 38.571
R9 VGND.n1 VGND.t4 33.077
R10 VGND.n7 VGND.n6 4.65
R11 VGND.n5 VGND.n4 4.65
R12 VGND.n3 VGND.n2 4.14
R13 VGND.n5 VGND.n3 0.134
R14 VGND.n7 VGND.n5 0.119
R15 VGND VGND.n7 0.024
R16 a_294_47.t0 a_294_47.t1 90
R17 VNB.t3 VNB.t0 6276.47
R18 VNB VNB.t2 6247.32
R19 VNB.t4 VNB.t3 3008.82
R20 VNB.t1 VNB.t5 2717.65
R21 VNB.t0 VNB.t1 2717.65
R22 VNB.t6 VNB.t4 2279.52
R23 VNB.t2 VNB.t6 2030.77
R24 A2_N.n0 A2_N.t0 369.643
R25 A2_N.n0 A2_N.t1 131.857
R26 A2_N A2_N.n0 116.355
R27 a_295_369.n2 a_295_369.n1 496.279
R28 a_295_369.n0 a_295_369.t3 295.334
R29 a_295_369.n1 a_295_369.t1 214.333
R30 a_295_369.n0 a_295_369.t4 154.239
R31 a_295_369.n1 a_295_369.n0 139.536
R32 a_295_369.t0 a_295_369.n2 61.562
R33 a_295_369.n2 a_295_369.t2 61.562
R34 VPWR.n8 VPWR.n7 308.015
R35 VPWR.n1 VPWR.n0 292.5
R36 VPWR.n2 VPWR.t5 233.762
R37 VPWR.n12 VPWR.t1 155.155
R38 VPWR.n0 VPWR.t4 113.89
R39 VPWR.n0 VPWR.t2 104.656
R40 VPWR.n7 VPWR.t3 61.562
R41 VPWR.n7 VPWR.t0 30.594
R42 VPWR.n2 VPWR.n1 7.814
R43 VPWR.n4 VPWR.n3 4.65
R44 VPWR.n6 VPWR.n5 4.65
R45 VPWR.n9 VPWR.n8 4.65
R46 VPWR.n11 VPWR.n10 4.65
R47 VPWR.n13 VPWR.n12 4.65
R48 VPWR.n4 VPWR.n2 0.143
R49 VPWR.n6 VPWR.n4 0.119
R50 VPWR.n9 VPWR.n6 0.119
R51 VPWR.n11 VPWR.n9 0.119
R52 VPWR.n13 VPWR.n11 0.119
R53 VPWR VPWR.n13 0.024
R54 VPB.t3 VPB.t5 509.034
R55 VPB.t4 VPB.t3 325.545
R56 VPB.t1 VPB.t4 287.071
R57 VPB.t5 VPB.t0 260.436
R58 VPB.t0 VPB.t6 248.598
R59 VPB.t2 VPB.t1 248.598
R60 VPB VPB.t2 213.084
R61 B1.n0 B1.t0 288.414
R62 B1.n0 B1.t1 195.228
R63 B1.n1 B1.n0 76
R64  B1.n1 10.573
R65 B1.n1 B1 2.04
R66 a_665_369.t0 a_665_369.t1 83.109
R67 a_84_21.n2 a_84_21.n1 250.1
R68 a_84_21.n1 a_84_21.t5 212.079
R69 a_84_21.n0 a_84_21.t6 212.079
R70 a_84_21.n2 a_84_21.t2 211.998
R71 a_84_21.n3 a_84_21.n2 149.808
R72 a_84_21.n1 a_84_21.t3 139.779
R73 a_84_21.n0 a_84_21.t4 139.779
R74 a_84_21.n1 a_84_21.n0 61.345
R75 a_84_21.t0 a_84_21.n3 47.71
R76 a_84_21.n3 a_84_21.t1 41.554
R77 X.n2 X.n1 146.372
R78 X.n2 X.n0 139.021
R79 X.n1 X.t1 26.595
R80 X.n1 X.t0 26.595
R81 X.n0 X.t3 24.923
R82 X.n0 X.t2 24.923
R83 X X.n2 4.145
R84 a_581_47.n0 a_581_47.t1 294.363
R85 a_581_47.t0 a_581_47.n0 38.571
R86 a_581_47.n0 a_581_47.t2 38.571
R87 B2.n0 B2.t0 299.374
R88 B2.n0 B2.t1 206.188
R89 B2 B2.n0 94.763
C0 VPWR VGND 0.11fF
C1 X VGND 0.21fF
C2 B2 B1 0.16fF
C3 A1_N A2_N 0.12fF
C4 VPWR X 0.24fF
C5 B2 VPWR 0.12fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__o2bb2a_4.ext - technology: sky130A

.subckt sky130_fd_sc_hd__o2bb2a_4 A2_N A1_N X B2 B1 VGND VPWR VNB VPB
X0 a_27_47.t1 a_415_21.t6 a_193_297.t1 VNB.t6 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 VPWR.t3 A2_N.t0 a_415_21.t1 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 a_415_21.t0 A1_N.t0 VPWR.t1 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 a_415_21.t2 A2_N.t1 a_717_47.t1 VNB.t7 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 a_193_297.t3 a_415_21.t7 VPWR.t9 VPB.t9 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 VPWR.t0 B1.t0 a_109_297.t1 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 VPWR.t7 a_193_297.t6 X.t7 VPB.t7 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 X.t3 a_193_297.t7 VGND.t7 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 a_109_297.t2 B2.t0 a_193_297.t4 VPB.t10 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 X.t6 a_193_297.t8 VPWR.t6 VPB.t6 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 a_717_47.t3 A1_N.t1 VGND.t3 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 a_717_47.t0 A2_N.t2 a_415_21.t4 VNB.t12 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 X.t2 a_193_297.t9 VGND.t6 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 a_193_297.t5 B2.t1 a_109_297.t3 VPB.t11 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14 a_27_47.t2 B2.t2 VGND.t8 VNB.t8 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X15 a_27_47.t4 B1.t1 VGND.t1 VNB.t10 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X16 VGND.t5 a_193_297.t10 X.t1 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X17 VGND.t2 A1_N.t2 a_717_47.t2 VNB.t13 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X18 VGND.t4 a_193_297.t11 X.t0 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X19 VGND.t9 B2.t3 a_27_47.t3 VNB.t9 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X20 a_193_297.t0 a_415_21.t8 a_27_47.t0 VNB.t5 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X21 VPWR.t5 a_193_297.t12 X.t5 VPB.t5 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X22 VPWR.t8 a_415_21.t9 a_193_297.t2 VPB.t8 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X23 X.t4 a_193_297.t13 VPWR.t4 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X24 VPWR.t11 A1_N.t3 a_415_21.t5 VPB.t13 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X25 a_109_297.t0 B1.t2 VPWR.t10 VPB.t12 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X26 a_415_21.t3 A2_N.t3 VPWR.t2 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X27 VGND.t0 B1.t3 a_27_47.t5 VNB.t11 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
R0 a_415_21.n6 a_415_21.n5 292.5
R1 a_415_21.n2 a_415_21.t9 212.079
R2 a_415_21.n1 a_415_21.t7 212.079
R3 a_415_21.n5 a_415_21.n0 201.489
R4 a_415_21.n4 a_415_21.n3 182.887
R5 a_415_21.n2 a_415_21.t6 139.779
R6 a_415_21.n1 a_415_21.t8 139.779
R7 a_415_21.n4 a_415_21.n2 119.848
R8 a_415_21.n5 a_415_21.n4 84.873
R9 a_415_21.n2 a_415_21.n1 61.345
R10 a_415_21.n0 a_415_21.t5 26.595
R11 a_415_21.n0 a_415_21.t3 26.595
R12 a_415_21.n6 a_415_21.t1 26.595
R13 a_415_21.t0 a_415_21.n6 26.595
R14 a_415_21.n3 a_415_21.t4 24.923
R15 a_415_21.n3 a_415_21.t2 24.923
R16 a_193_297.n12 a_193_297.n0 362.895
R17 a_193_297.n1 a_193_297.t6 212.079
R18 a_193_297.n3 a_193_297.t8 212.079
R19 a_193_297.n6 a_193_297.t12 212.079
R20 a_193_297.n7 a_193_297.t13 212.079
R21 a_193_297.n1 a_193_297.t11 139.779
R22 a_193_297.n3 a_193_297.t9 139.779
R23 a_193_297.n6 a_193_297.t10 139.779
R24 a_193_297.n7 a_193_297.t7 139.779
R25 a_193_297.n11 a_193_297.n10 124.292
R26 a_193_297.n13 a_193_297.n12 122.803
R27 a_193_297.n5 a_193_297.n2 101.6
R28 a_193_297.n5 a_193_297.n4 76
R29 a_193_297.n9 a_193_297.n8 76
R30 a_193_297.n8 a_193_297.n7 49.66
R31 a_193_297.n2 a_193_297.n1 35.054
R32 a_193_297.n11 a_193_297.n9 33.657
R33 a_193_297.n0 a_193_297.t4 26.595
R34 a_193_297.n0 a_193_297.t5 26.595
R35 a_193_297.t2 a_193_297.n13 26.595
R36 a_193_297.n13 a_193_297.t3 26.595
R37 a_193_297.n9 a_193_297.n5 25.6
R38 a_193_297.n10 a_193_297.t1 24.923
R39 a_193_297.n10 a_193_297.t0 24.923
R40 a_193_297.n4 a_193_297.n3 23.369
R41 a_193_297.n8 a_193_297.n6 11.684
R42 a_193_297.n12 a_193_297.n11 5.404
R43 a_27_47.t1 a_27_47.n3 224.124
R44 a_27_47.n1 a_27_47.t5 128.218
R45 a_27_47.n1 a_27_47.n0 52.624
R46 a_27_47.n3 a_27_47.n1 51.157
R47 a_27_47.n3 a_27_47.n2 42.273
R48 a_27_47.n2 a_27_47.t0 24.923
R49 a_27_47.n2 a_27_47.t4 24.923
R50 a_27_47.n0 a_27_47.t3 24.923
R51 a_27_47.n0 a_27_47.t2 24.923
R52 VNB VNB.t11 6078.09
R53 VNB.t6 VNB.t0 4545.05
R54 VNB.t3 VNB.t1 2030.77
R55 VNB.t2 VNB.t3 2030.77
R56 VNB.t4 VNB.t2 2030.77
R57 VNB.t13 VNB.t4 2030.77
R58 VNB.t12 VNB.t13 2030.77
R59 VNB.t7 VNB.t12 2030.77
R60 VNB.t0 VNB.t7 2030.77
R61 VNB.t5 VNB.t6 2030.77
R62 VNB.t10 VNB.t5 2030.77
R63 VNB.t9 VNB.t10 2030.77
R64 VNB.t8 VNB.t9 2030.77
R65 VNB.t11 VNB.t8 2030.77
R66 A2_N.n0 A2_N.t3 212.079
R67 A2_N.n1 A2_N.t0 212.079
R68 A2_N.n0 A2_N.t2 139.779
R69 A2_N.n1 A2_N.t1 139.779
R70 A2_N A2_N.n2 95.2
R71 A2_N.n2 A2_N.n1 31.403
R72 A2_N.n2 A2_N.n0 29.942
R73 VPWR.n26 VPWR.n25 314.004
R74 VPWR.n12 VPWR.n11 314.004
R75 VPWR.n1 VPWR.n0 312.468
R76 VPWR.n20 VPWR.n19 292.5
R77 VPWR.n16 VPWR.n15 292.5
R78 VPWR.n35 VPWR.t10 204.191
R79 VPWR.n2 VPWR.t7 200.67
R80 VPWR.n6 VPWR.n5 171.981
R81 VPWR.n15 VPWR.t1 26.595
R82 VPWR.n19 VPWR.t8 26.595
R83 VPWR.n25 VPWR.t9 26.595
R84 VPWR.n25 VPWR.t0 26.595
R85 VPWR.n11 VPWR.t2 26.595
R86 VPWR.n11 VPWR.t3 26.595
R87 VPWR.n5 VPWR.t4 26.595
R88 VPWR.n5 VPWR.t11 26.595
R89 VPWR.n0 VPWR.t6 26.595
R90 VPWR.n0 VPWR.t5 26.595
R91 VPWR.n13 VPWR.n12 7.905
R92 VPWR.n4 VPWR.n3 4.65
R93 VPWR.n8 VPWR.n7 4.65
R94 VPWR.n10 VPWR.n9 4.65
R95 VPWR.n14 VPWR.n13 4.65
R96 VPWR.n18 VPWR.n17 4.65
R97 VPWR.n22 VPWR.n21 4.65
R98 VPWR.n24 VPWR.n23 4.65
R99 VPWR.n28 VPWR.n27 4.65
R100 VPWR.n30 VPWR.n29 4.65
R101 VPWR.n32 VPWR.n31 4.65
R102 VPWR.n34 VPWR.n33 4.65
R103 VPWR.n36 VPWR.n35 4.65
R104 VPWR.n17 VPWR.n16 4.27
R105 VPWR.n21 VPWR.n20 4.011
R106 VPWR.n2 VPWR.n1 3.784
R107 VPWR.n7 VPWR.n6 1.882
R108 VPWR.n27 VPWR.n26 0.376
R109 VPWR.n4 VPWR.n2 0.233
R110 VPWR.n8 VPWR.n4 0.119
R111 VPWR.n10 VPWR.n8 0.119
R112 VPWR.n14 VPWR.n10 0.119
R113 VPWR.n18 VPWR.n14 0.119
R114 VPWR.n22 VPWR.n18 0.119
R115 VPWR.n24 VPWR.n22 0.119
R116 VPWR.n28 VPWR.n24 0.119
R117 VPWR.n30 VPWR.n28 0.119
R118 VPWR.n32 VPWR.n30 0.119
R119 VPWR.n34 VPWR.n32 0.119
R120 VPWR.n36 VPWR.n34 0.119
R121 VPWR VPWR.n36 0.022
R122 VPB.t8 VPB.t1 556.386
R123 VPB.t6 VPB.t7 248.598
R124 VPB.t5 VPB.t6 248.598
R125 VPB.t4 VPB.t5 248.598
R126 VPB.t13 VPB.t4 248.598
R127 VPB.t2 VPB.t13 248.598
R128 VPB.t3 VPB.t2 248.598
R129 VPB.t1 VPB.t3 248.598
R130 VPB.t9 VPB.t8 248.598
R131 VPB.t0 VPB.t9 248.598
R132 VPB.t10 VPB.t0 248.598
R133 VPB.t11 VPB.t10 248.598
R134 VPB.t12 VPB.t11 248.598
R135 VPB VPB.t12 192.367
R136 A1_N.n1 A1_N.t3 241.534
R137 A1_N.n0 A1_N.t0 236.179
R138 A1_N.n2 A1_N.n0 175.788
R139 A1_N.n1 A1_N.t2 169.234
R140 A1_N.n0 A1_N.t1 163.879
R141 A1_N.n2 A1_N.n1 76
R142 A1_N A1_N.n2 1.955
R143 a_717_47.n1 a_717_47.n0 199.576
R144 a_717_47.n0 a_717_47.t2 24.923
R145 a_717_47.n0 a_717_47.t0 24.923
R146 a_717_47.t1 a_717_47.n1 24.923
R147 a_717_47.n1 a_717_47.t3 24.923
R148 B1.n1 B1.t2 241.534
R149 B1.n0 B1.t0 241.534
R150 B1.n1 B1.t3 169.234
R151 B1.n0 B1.t1 169.234
R152 B1.n2 B1.n0 168.803
R153 B1.n2 B1.n1 76
R154 B1 B1.n2 6.281
R155 a_109_297.n1 a_109_297.n0 496.201
R156 a_109_297.n0 a_109_297.t3 26.595
R157 a_109_297.n0 a_109_297.t0 26.595
R158 a_109_297.t1 a_109_297.n1 26.595
R159 a_109_297.n1 a_109_297.t2 26.595
R160 X.n2 X.n0 203.821
R161 X.n2 X.n1 98.532
R162 X.n5 X.n3 88.89
R163 X.n5 X.n4 52.624
R164 X X.n2 29.062
R165 X.n1 X.t7 26.595
R166 X.n1 X.t6 26.595
R167 X.n0 X.t5 26.595
R168 X.n0 X.t4 26.595
R169  X.n5 26.392
R170 X.n3 X.t1 24.923
R171 X.n3 X.t3 24.923
R172 X.n4 X.t0 24.923
R173 X.n4 X.t2 24.923
R174  X 14.268
R175 VGND.n0 VGND.t4 197.839
R176 VGND.n15 VGND.t3 193.925
R177 VGND.n2 VGND.n1 115.464
R178 VGND.n25 VGND.n24 115.464
R179 VGND.n31 VGND.n30 115.464
R180 VGND.n8 VGND.n7 74.837
R181 VGND.n1 VGND.t6 24.923
R182 VGND.n1 VGND.t5 24.923
R183 VGND.n7 VGND.t7 24.923
R184 VGND.n7 VGND.t2 24.923
R185 VGND.n24 VGND.t1 24.923
R186 VGND.n24 VGND.t9 24.923
R187 VGND.n30 VGND.t8 24.923
R188 VGND.n30 VGND.t0 24.923
R189 VGND.n9 VGND.n8 11.294
R190 VGND.n16 VGND.n15 11.294
R191 VGND.n26 VGND.n25 6.776
R192 VGND.n3 VGND.n2 5.27
R193 VGND.n4 VGND.n3 4.65
R194 VGND.n6 VGND.n5 4.65
R195 VGND.n10 VGND.n9 4.65
R196 VGND.n12 VGND.n11 4.65
R197 VGND.n14 VGND.n13 4.65
R198 VGND.n17 VGND.n16 4.65
R199 VGND.n19 VGND.n18 4.65
R200 VGND.n21 VGND.n20 4.65
R201 VGND.n23 VGND.n22 4.65
R202 VGND.n27 VGND.n26 4.65
R203 VGND.n29 VGND.n28 4.65
R204 VGND.n33 VGND.n32 4.65
R205 VGND.n32 VGND.n31 0.752
R206 VGND.n4 VGND.n0 0.657
R207 VGND.n6 VGND.n4 0.119
R208 VGND.n10 VGND.n6 0.119
R209 VGND.n12 VGND.n10 0.119
R210 VGND.n14 VGND.n12 0.119
R211 VGND.n17 VGND.n14 0.119
R212 VGND.n19 VGND.n17 0.119
R213 VGND.n21 VGND.n19 0.119
R214 VGND.n23 VGND.n21 0.119
R215 VGND.n27 VGND.n23 0.119
R216 VGND.n29 VGND.n27 0.119
R217 VGND.n33 VGND.n29 0.119
R218 VGND.n34 VGND.n33 0.119
R219 VGND VGND.n34 0.022
R220 B2.n0 B2.t0 212.079
R221 B2.n1 B2.t1 212.079
R222 B2.n0 B2.t3 139.779
R223 B2.n1 B2.t2 139.779
R224 B2 B2.n2 77.303
R225 B2.n2 B2.n0 30.672
R226 B2.n2 B2.n1 30.672
C0 X VPWR 0.52fF
C1 A1_N A2_N 0.35fF
C2 X VGND 0.47fF
C3 VGND VPWR 0.12fF
C4 VPB VPWR 0.15fF
C5 B1 B2 0.30fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__o2bb2ai_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__o2bb2ai_1 Y A1_N A2_N B2 B1 VGND VPWR VNB VPB
X0 VPWR.t2 A2_N.t0 a_112_297.t0 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 Y.t1 a_112_297.t3 VPWR.t0 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 VGND.t2 B2.t0 a_394_47.t2 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 a_112_297.t1 A2_N.t1 a_112_47.t1 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 a_112_47.t0 A1_N.t0 VGND.t0 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 a_112_297.t2 A1_N.t1 VPWR.t3 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 VPWR.t1 B1.t0 a_478_297.t0 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 a_394_47.t0 a_112_297.t4 Y.t2 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 a_394_47.t1 B1.t1 VGND.t1 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 a_478_297.t1 B2.t1 Y.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
R0 A2_N.n0 A2_N.t0 241.534
R1 A2_N.n0 A2_N.t1 169.234
R2 A2_N A2_N.n0 87.635
R3 a_112_297.n2 a_112_297.n1 222.526
R4 a_112_297.n0 a_112_297.t3 212.079
R5 a_112_297.n1 a_112_297.n0 150.49
R6 a_112_297.n0 a_112_297.t4 139.779
R7 a_112_297.n1 a_112_297.t1 117.89
R8 a_112_297.t0 a_112_297.n2 26.595
R9 a_112_297.n2 a_112_297.t2 26.595
R10 VPWR.n2 VPWR.t1 158.489
R11 VPWR.n9 VPWR.t3 154.252
R12 VPWR.n4 VPWR.n3 146.25
R13 VPWR.n1 VPWR.n0 146.25
R14 VPWR.n0 VPWR.t0 42.355
R15 VPWR.n3 VPWR.t2 34.475
R16 VPWR.n6 VPWR.n5 4.65
R17 VPWR.n8 VPWR.n7 4.65
R18 VPWR.n10 VPWR.n9 4.65
R19 VPWR.n2 VPWR.n1 4.044
R20 VPWR.n6 VPWR.n2 0.148
R21 VPWR.n8 VPWR.n6 0.119
R22 VPWR.n10 VPWR.n8 0.119
R23 VPWR.n5 VPWR.n4 0.065
R24 VPWR VPWR.n10 0.022
R25 VPB.t3 VPB.t1 585.981
R26 VPB.t0 VPB.t2 248.598
R27 VPB.t1 VPB.t0 248.598
R28 VPB.t4 VPB.t3 248.598
R29 VPB VPB.t4 201.246
R30 Y.n1 Y.t2 197.716
R31 Y Y.n0 156.262
R32 Y.n0 Y.t0 26.595
R33 Y.n0 Y.t1 26.595
R34 Y Y.n1 6.4
R35 B2.n0 B2.t1 241.534
R36 B2.n0 B2.t0 169.234
R37 B2 B2.n0 96.043
R38 a_394_47.n0 a_394_47.t1 229.986
R39 a_394_47.n0 a_394_47.t2 24.923
R40 a_394_47.t0 a_394_47.n0 24.923
R41 VGND.n1 VGND.n0 120.07
R42 VGND.n1 VGND.t0 105.248
R43 VGND.n0 VGND.t1 24.923
R44 VGND.n0 VGND.t2 24.923
R45 VGND VGND.n1 0.044
R46 VNB VNB.t1 6150.61
R47 VNB.t2 VNB.t0 5076.92
R48 VNB.t4 VNB.t3 2030.77
R49 VNB.t0 VNB.t4 2030.77
R50 VNB.t1 VNB.t2 1740.66
R51 a_112_47.t0 a_112_47.t1 38.769
R52 A1_N.n0 A1_N.t1 229.558
R53 A1_N.n0 A1_N.t0 157.258
R54 A1_N A1_N.n0 81.333
R55 B1.n0 B1.t0 229.558
R56 B1.n0 B1.t1 157.258
R57 B1 B1.n0 78.011
R58 a_478_297.t0 a_478_297.t1 53.19
C0 VPWR Y 0.20fF
C1 B2 VPWR 0.17fF
C2 B2 Y 0.16fF
C3 A1_N A2_N 0.11fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__o2bb2ai_2.ext - technology: sky130A

.subckt sky130_fd_sc_hd__o2bb2ai_2 B2 Y A1_N A2_N B1 VGND VPWR VNB VPB
X0 a_113_297.t1 A2_N.t0 VPWR.t3 VPB.t5 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_113_47.t1 A2_N.t1 a_113_297.t3 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 VPWR.t5 B1.t0 a_730_297.t3 VPB.t7 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 VPWR.t2 A2_N.t2 a_113_297.t0 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 a_730_297.t0 B2.t0 Y.t5 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 a_471_47.t3 B2.t1 VGND.t1 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 a_471_47.t5 B1.t1 VGND.t3 VNB.t6 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 Y.t4 B2.t2 a_730_297.t1 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 a_113_297.t2 A2_N.t3 a_113_47.t0 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 a_113_47.t2 A1_N.t0 VGND.t4 VNB.t8 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 VGND.t5 A1_N.t1 a_113_47.t3 VNB.t9 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 VGND.t0 B2.t3 a_471_47.t2 VNB.t5 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 VPWR.t0 a_113_297.t6 Y.t1 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13 a_113_297.t5 A1_N.t2 VPWR.t7 VPB.t9 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14 Y.t0 a_113_297.t7 VPWR.t1 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 a_730_297.t2 B1.t2 VPWR.t6 VPB.t8 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16 Y.t2 a_113_297.t8 a_471_47.t1 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X17 a_471_47.t0 a_113_297.t9 Y.t3 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X18 VPWR.t4 A1_N.t3 a_113_297.t4 VPB.t6 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X19 VGND.t2 B1.t3 a_471_47.t4 VNB.t7 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
R0 A2_N.n0 A2_N.t0 212.079
R1 A2_N.n1 A2_N.t2 212.079
R2 A2_N.n0 A2_N.t1 139.779
R3 A2_N.n1 A2_N.t3 139.779
R4 A2_N A2_N.n2 77.163
R5 A2_N.n2 A2_N.n0 31.403
R6 A2_N.n2 A2_N.n1 29.942
R7 VPWR.n16 VPWR.n15 314.004
R8 VPWR.n1 VPWR.n0 311.363
R9 VPWR.n10 VPWR.n9 292.5
R10 VPWR.n6 VPWR.n5 292.5
R11 VPWR.n2 VPWR.t5 212.532
R12 VPWR.n20 VPWR.t7 198.576
R13 VPWR.n0 VPWR.t6 33.49
R14 VPWR.n5 VPWR.t1 26.595
R15 VPWR.n9 VPWR.t4 26.595
R16 VPWR.n15 VPWR.t3 26.595
R17 VPWR.n15 VPWR.t2 26.595
R18 VPWR.n0 VPWR.t0 26.595
R19 VPWR.n4 VPWR.n3 4.65
R20 VPWR.n8 VPWR.n7 4.65
R21 VPWR.n12 VPWR.n11 4.65
R22 VPWR.n14 VPWR.n13 4.65
R23 VPWR.n17 VPWR.n16 4.65
R24 VPWR.n19 VPWR.n18 4.65
R25 VPWR.n21 VPWR.n20 4.65
R26 VPWR.n2 VPWR.n1 4.099
R27 VPWR.n11 VPWR.n10 2.101
R28 VPWR.n7 VPWR.n6 0.764
R29 VPWR.n4 VPWR.n2 0.138
R30 VPWR.n8 VPWR.n4 0.119
R31 VPWR.n12 VPWR.n8 0.119
R32 VPWR.n14 VPWR.n12 0.119
R33 VPWR.n17 VPWR.n14 0.119
R34 VPWR.n19 VPWR.n17 0.119
R35 VPWR.n21 VPWR.n19 0.119
R36 VPWR VPWR.n21 0.02
R37 a_113_297.n6 a_113_297.n5 292.5
R38 a_113_297.n0 a_113_297.t6 212.079
R39 a_113_297.n1 a_113_297.t7 212.079
R40 a_113_297.n5 a_113_297.n4 201.489
R41 a_113_297.n3 a_113_297.n2 177.056
R42 a_113_297.n0 a_113_297.t9 139.779
R43 a_113_297.n1 a_113_297.t8 139.779
R44 a_113_297.n3 a_113_297.n1 106.672
R45 a_113_297.n5 a_113_297.n3 81.975
R46 a_113_297.n1 a_113_297.n0 61.345
R47 a_113_297.n4 a_113_297.t0 26.595
R48 a_113_297.n4 a_113_297.t5 26.595
R49 a_113_297.n6 a_113_297.t4 26.595
R50 a_113_297.t1 a_113_297.n6 26.595
R51 a_113_297.n2 a_113_297.t3 24.923
R52 a_113_297.n2 a_113_297.t2 24.923
R53 VPB.t6 VPB.t0 562.305
R54 VPB.t1 VPB.t8 269.314
R55 VPB.t2 VPB.t7 248.598
R56 VPB.t3 VPB.t2 248.598
R57 VPB.t8 VPB.t3 248.598
R58 VPB.t0 VPB.t1 248.598
R59 VPB.t5 VPB.t6 248.598
R60 VPB.t4 VPB.t5 248.598
R61 VPB.t9 VPB.t4 248.598
R62 VPB VPB.t9 201.246
R63 a_113_47.n1 a_113_47.n0 199.576
R64 a_113_47.n0 a_113_47.t0 24.923
R65 a_113_47.n0 a_113_47.t2 24.923
R66 a_113_47.n1 a_113_47.t3 24.923
R67 a_113_47.t1 a_113_47.n1 24.923
R68 VNB VNB.t8 6150.61
R69 VNB.t9 VNB.t1 4593.41
R70 VNB.t0 VNB.t7 2200
R71 VNB.t5 VNB.t6 2030.77
R72 VNB.t2 VNB.t5 2030.77
R73 VNB.t7 VNB.t2 2030.77
R74 VNB.t1 VNB.t0 2030.77
R75 VNB.t4 VNB.t9 2030.77
R76 VNB.t3 VNB.t4 2030.77
R77 VNB.t8 VNB.t3 2030.77
R78 B1.n0 B1.t0 241.534
R79 B1.n1 B1.t2 241.534
R80 B1.n0 B1.t1 169.234
R81 B1.n1 B1.t3 169.234
R82 B1.n2 B1.n1 168.803
R83 B1.n2 B1.n0 76
R84 B1 B1.n2 7.348
R85 a_730_297.n1 a_730_297.n0 496.201
R86 a_730_297.n0 a_730_297.t3 26.595
R87 a_730_297.n0 a_730_297.t0 26.595
R88 a_730_297.n1 a_730_297.t1 26.595
R89 a_730_297.t2 a_730_297.n1 26.595
R90 B2.n0 B2.t0 212.079
R91 B2.n1 B2.t2 212.079
R92 B2.n0 B2.t3 139.779
R93 B2.n1 B2.t1 139.779
R94 B2 B2.n2 82.72
R95 B2.n2 B2.n0 30.672
R96 B2.n2 B2.n1 30.672
R97 Y.n2 Y.n1 364.632
R98 Y Y.n3 115.957
R99 Y.n2 Y.n0 98.704
R100 Y.n1 Y.t5 26.595
R101 Y.n1 Y.t4 26.595
R102 Y.n0 Y.t1 26.595
R103 Y.n0 Y.t0 26.595
R104 Y.n3 Y.t3 24.923
R105 Y.n3 Y.t2 24.923
R106 Y Y.n2 9.174
R107 VGND.n10 VGND.t5 193.925
R108 VGND.n3 VGND.n0 126.027
R109 VGND.n2 VGND.n1 115.464
R110 VGND.n19 VGND.t4 111.584
R111 VGND.n0 VGND.t3 24.923
R112 VGND.n0 VGND.t0 24.923
R113 VGND.n1 VGND.t1 24.923
R114 VGND.n1 VGND.t2 24.923
R115 VGND.n3 VGND.n2 13.328
R116 VGND.n20 VGND.n19 8.414
R117 VGND.n11 VGND.n10 8.282
R118 VGND.n5 VGND.n4 4.65
R119 VGND.n7 VGND.n6 4.65
R120 VGND.n9 VGND.n8 4.65
R121 VGND.n12 VGND.n11 4.65
R122 VGND.n14 VGND.n13 4.65
R123 VGND.n16 VGND.n15 4.65
R124 VGND.n18 VGND.n17 4.65
R125 VGND.n5 VGND.n3 0.357
R126 VGND.n7 VGND.n5 0.119
R127 VGND.n9 VGND.n7 0.119
R128 VGND.n12 VGND.n9 0.119
R129 VGND.n14 VGND.n12 0.119
R130 VGND.n16 VGND.n14 0.119
R131 VGND.n18 VGND.n16 0.119
R132 VGND.n20 VGND.n18 0.119
R133 VGND VGND.n20 0.02
R134 a_471_47.t1 a_471_47.n3 218.837
R135 a_471_47.n1 a_471_47.t5 128.218
R136 a_471_47.n1 a_471_47.n0 52.624
R137 a_471_47.n3 a_471_47.n1 49.688
R138 a_471_47.n3 a_471_47.n2 42.724
R139 a_471_47.n2 a_471_47.t4 31.384
R140 a_471_47.n2 a_471_47.t0 24.923
R141 a_471_47.n0 a_471_47.t2 24.923
R142 a_471_47.n0 a_471_47.t3 24.923
R143 A1_N.n1 A1_N.t2 236.179
R144 A1_N.n0 A1_N.t3 236.179
R145 A1_N.n2 A1_N.n0 168.803
R146 A1_N.n1 A1_N.t0 163.879
R147 A1_N.n0 A1_N.t1 163.879
R148 A1_N.n2 A1_N.n1 76
R149 A1_N A1_N.n2 7.348
C0 VPWR VGND 0.12fF
C1 B1 Y 0.23fF
C2 B1 B2 0.30fF
C3 VPWR VPB 0.11fF
C4 A1_N A2_N 0.34fF
C5 VPWR Y 0.26fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__o2bb2ai_4.ext - technology: sky130A

.subckt sky130_fd_sc_hd__o2bb2ai_4 A1_N B1 B2 A2_N Y VGND VPWR VNB VPB
X0 a_1241_297.t7 B1.t0 VPWR.t13 VPB.t17 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_113_47.t3 A2_N.t0 VPWR.t4 VPB.t8 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 a_807_47.t5 a_113_47.t12 Y.t11 VNB.t5 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 VGND.t3 B2.t0 a_807_47.t6 VNB.t6 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 a_113_47.t7 A2_N.t1 a_27_47.t3 VNB.t11 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 VGND.t2 B2.t1 a_807_47.t7 VNB.t7 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 VPWR.t5 A2_N.t2 a_113_47.t2 VPB.t9 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 VPWR.t12 B1.t1 a_1241_297.t6 VPB.t16 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 Y.t10 a_113_47.t13 a_807_47.t4 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 a_1241_297.t2 B2.t2 Y.t2 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 Y.t3 B2.t3 a_1241_297.t3 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 Y.t9 a_113_47.t14 a_807_47.t3 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 a_27_47.t2 A2_N.t3 a_113_47.t6 VNB.t10 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 a_807_47.t0 B2.t4 VGND.t1 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14 VPWR.t14 A1_N.t0 a_113_47.t10 VPB.t18 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 a_113_47.t5 A2_N.t4 a_27_47.t1 VNB.t9 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X16 a_27_47.t0 A2_N.t5 a_113_47.t4 VNB.t8 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X17 a_807_47.t1 B2.t5 VGND.t0 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X18 a_27_47.t5 A1_N.t1 VGND.t9 VNB.t17 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X19 a_807_47.t11 B1.t2 VGND.t8 VNB.t16 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X20 a_1241_297.t0 B2.t6 Y.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X21 VPWR.t0 a_113_47.t15 Y.t7 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X22 a_27_47.t6 A1_N.t2 VGND.t10 VNB.t18 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X23 a_807_47.t10 B1.t3 VGND.t7 VNB.t15 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X24 a_113_47.t11 A1_N.t3 VPWR.t15 VPB.t19 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X25 Y.t1 B2.t7 a_1241_297.t1 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X26 Y.t6 a_113_47.t16 VPWR.t1 VPB.t5 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X27 VPWR.t2 a_113_47.t17 Y.t5 VPB.t6 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X28 a_113_47.t1 A2_N.t6 VPWR.t6 VPB.t10 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X29 a_1241_297.t5 B1.t4 VPWR.t11 VPB.t15 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X30 VGND.t11 A1_N.t4 a_27_47.t7 VNB.t19 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X31 VGND.t6 B1.t5 a_807_47.t9 VNB.t14 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X32 Y.t4 a_113_47.t18 VPWR.t3 VPB.t7 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X33 VGND.t4 A1_N.t5 a_27_47.t4 VNB.t12 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X34 VGND.t5 B1.t6 a_807_47.t8 VNB.t13 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X35 VPWR.t10 B1.t7 a_1241_297.t4 VPB.t14 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X36 VPWR.t8 A1_N.t6 a_113_47.t8 VPB.t12 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X37 a_113_47.t9 A1_N.t7 VPWR.t9 VPB.t13 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X38 VPWR.t7 A2_N.t7 a_113_47.t0 VPB.t11 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X39 a_807_47.t2 a_113_47.t19 Y.t8 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
R0 B1.n0 B1.t4 212.079
R1 B1.n2 B1.t7 212.079
R2 B1.n6 B1.t0 212.079
R3 B1.n5 B1.t1 212.079
R4 B1.n0 B1.t3 139.779
R5 B1.n2 B1.t6 139.779
R6 B1.n6 B1.t2 139.779
R7 B1.n5 B1.t5 139.779
R8 B1.n4 B1.n1 96.723
R9 B1.n4 B1.n3 76
R10 B1 B1.n7 49.208
R11 B1.n7 B1.n5 30.363
R12 B1.n1 B1.n0 26.29
R13 B1.n7 B1.n6 19.893
R14 B1.n3 B1.n2 14.606
R15 B1 B1.n4 4.571
R16 VPWR.n45 VPWR.t6 198.576
R17 VPWR.n14 VPWR.t0 198.576
R18 VPWR.n3 VPWR.n0 176.868
R19 VPWR.n41 VPWR.n40 171.981
R20 VPWR.n36 VPWR.n35 171.981
R21 VPWR.n30 VPWR.n29 171.981
R22 VPWR.n19 VPWR.n18 171.981
R23 VPWR.n2 VPWR.n1 171.981
R24 VPWR.n25 VPWR.n24 63.687
R25 VPWR.n24 VPWR.t3 62.886
R26 VPWR.n24 VPWR.t14 62.885
R27 VPWR.n40 VPWR.t4 26.595
R28 VPWR.n40 VPWR.t5 26.595
R29 VPWR.n35 VPWR.t9 26.595
R30 VPWR.n35 VPWR.t7 26.595
R31 VPWR.n29 VPWR.t15 26.595
R32 VPWR.n29 VPWR.t8 26.595
R33 VPWR.n18 VPWR.t1 26.595
R34 VPWR.n18 VPWR.t2 26.595
R35 VPWR.n1 VPWR.t13 26.595
R36 VPWR.n1 VPWR.t12 26.595
R37 VPWR.n0 VPWR.t11 26.595
R38 VPWR.n0 VPWR.t10 26.595
R39 VPWR.n31 VPWR.n30 4.894
R40 VPWR.n5 VPWR.n4 4.65
R41 VPWR.n7 VPWR.n6 4.65
R42 VPWR.n9 VPWR.n8 4.65
R43 VPWR.n11 VPWR.n10 4.65
R44 VPWR.n13 VPWR.n12 4.65
R45 VPWR.n15 VPWR.n14 4.65
R46 VPWR.n17 VPWR.n16 4.65
R47 VPWR.n21 VPWR.n20 4.65
R48 VPWR.n23 VPWR.n22 4.65
R49 VPWR.n26 VPWR.n25 4.65
R50 VPWR.n28 VPWR.n27 4.65
R51 VPWR.n32 VPWR.n31 4.65
R52 VPWR.n34 VPWR.n33 4.65
R53 VPWR.n37 VPWR.n36 4.65
R54 VPWR.n39 VPWR.n38 4.65
R55 VPWR.n42 VPWR.n41 4.65
R56 VPWR.n44 VPWR.n43 4.65
R57 VPWR.n46 VPWR.n45 4.65
R58 VPWR.n3 VPWR.n2 3.941
R59 VPWR.n20 VPWR.n19 1.129
R60 VPWR.n5 VPWR.n3 0.285
R61 VPWR.n7 VPWR.n5 0.119
R62 VPWR.n9 VPWR.n7 0.119
R63 VPWR.n11 VPWR.n9 0.119
R64 VPWR.n13 VPWR.n11 0.119
R65 VPWR.n15 VPWR.n13 0.119
R66 VPWR.n17 VPWR.n15 0.119
R67 VPWR.n21 VPWR.n17 0.119
R68 VPWR.n23 VPWR.n21 0.119
R69 VPWR.n26 VPWR.n23 0.119
R70 VPWR.n28 VPWR.n26 0.119
R71 VPWR.n32 VPWR.n28 0.119
R72 VPWR.n34 VPWR.n32 0.119
R73 VPWR.n37 VPWR.n34 0.119
R74 VPWR.n39 VPWR.n37 0.119
R75 VPWR.n42 VPWR.n39 0.119
R76 VPWR.n44 VPWR.n42 0.119
R77 VPWR.n46 VPWR.n44 0.119
R78 VPWR VPWR.n46 0.024
R79 a_1241_297.n1 a_1241_297.t1 224.711
R80 a_1241_297.n3 a_1241_297.t5 179.288
R81 a_1241_297.n1 a_1241_297.n0 154.573
R82 a_1241_297.n3 a_1241_297.n2 110.76
R83 a_1241_297.n5 a_1241_297.n4 90.234
R84 a_1241_297.n4 a_1241_297.n1 64.951
R85 a_1241_297.n4 a_1241_297.n3 64.951
R86 a_1241_297.n0 a_1241_297.t3 26.595
R87 a_1241_297.n0 a_1241_297.t0 26.595
R88 a_1241_297.n2 a_1241_297.t4 26.595
R89 a_1241_297.n2 a_1241_297.t7 26.595
R90 a_1241_297.t6 a_1241_297.n5 26.595
R91 a_1241_297.n5 a_1241_297.t2 26.595
R92 VPB.t4 VPB.t1 556.386
R93 VPB.t18 VPB.t7 538.629
R94 VPB.t14 VPB.t15 248.598
R95 VPB.t17 VPB.t14 248.598
R96 VPB.t16 VPB.t17 248.598
R97 VPB.t2 VPB.t16 248.598
R98 VPB.t3 VPB.t2 248.598
R99 VPB.t0 VPB.t3 248.598
R100 VPB.t1 VPB.t0 248.598
R101 VPB.t5 VPB.t4 248.598
R102 VPB.t6 VPB.t5 248.598
R103 VPB.t7 VPB.t6 248.598
R104 VPB.t19 VPB.t18 248.598
R105 VPB.t12 VPB.t19 248.598
R106 VPB.t13 VPB.t12 248.598
R107 VPB.t11 VPB.t13 248.598
R108 VPB.t8 VPB.t11 248.598
R109 VPB.t9 VPB.t8 248.598
R110 VPB.t10 VPB.t9 248.598
R111 VPB VPB.t10 210.124
R112 A2_N.n0 A2_N.t7 212.079
R113 A2_N.n2 A2_N.t0 212.079
R114 A2_N.n7 A2_N.t2 212.079
R115 A2_N.n5 A2_N.t6 212.079
R116 A2_N.n0 A2_N.t5 139.779
R117 A2_N.n2 A2_N.t1 139.779
R118 A2_N.n7 A2_N.t3 139.779
R119 A2_N.n5 A2_N.t4 139.779
R120 A2_N.n9 A2_N.n6 96.723
R121 A2_N.n4 A2_N.n1 96.723
R122 A2_N.n4 A2_N.n3 76
R123 A2_N.n9 A2_N.n8 76
R124 A2_N.n1 A2_N.n0 20.448
R125 A2_N.n6 A2_N.n5 14.606
R126 A2_N A2_N.n4 13.104
R127 A2_N.n3 A2_N.n2 8.763
R128 A2_N A2_N.n9 7.619
R129 A2_N.n8 A2_N.n7 2.921
R130 a_113_47.n15 a_113_47.t18 216.46
R131 a_113_47.n5 a_113_47.t15 212.079
R132 a_113_47.n8 a_113_47.t16 212.079
R133 a_113_47.n11 a_113_47.t17 212.079
R134 a_113_47.n5 a_113_47.t19 144.16
R135 a_113_47.n15 a_113_47.t14 139.779
R136 a_113_47.n12 a_113_47.t12 139.779
R137 a_113_47.n7 a_113_47.t13 139.779
R138 a_113_47.n2 a_113_47.n0 133.853
R139 a_113_47.n4 a_113_47.n3 110.761
R140 a_113_47.n23 a_113_47.n22 110.761
R141 a_113_47.n19 a_113_47.n18 110.76
R142 a_113_47.n21 a_113_47.n20 110.76
R143 a_113_47.n4 a_113_47.n2 97.997
R144 a_113_47.n10 a_113_47.n6 96.723
R145 a_113_47.n2 a_113_47.n1 92.5
R146 a_113_47.n19 a_113_47.n17 87.717
R147 a_113_47.n17 a_113_47.n16 76
R148 a_113_47.n10 a_113_47.n9 76
R149 a_113_47.n14 a_113_47.n13 76
R150 a_113_47.n21 a_113_47.n19 44.423
R151 a_113_47.n22 a_113_47.n4 44.423
R152 a_113_47.n22 a_113_47.n21 44.423
R153 a_113_47.n18 a_113_47.t10 26.595
R154 a_113_47.n18 a_113_47.t11 26.595
R155 a_113_47.n20 a_113_47.t8 26.595
R156 a_113_47.n20 a_113_47.t9 26.595
R157 a_113_47.n3 a_113_47.t2 26.595
R158 a_113_47.n3 a_113_47.t1 26.595
R159 a_113_47.n23 a_113_47.t0 26.595
R160 a_113_47.t3 a_113_47.n23 26.595
R161 a_113_47.n0 a_113_47.t4 24.923
R162 a_113_47.n0 a_113_47.t7 24.923
R163 a_113_47.n1 a_113_47.t6 24.923
R164 a_113_47.n1 a_113_47.t5 24.923
R165 a_113_47.n14 a_113_47.n10 20.723
R166 a_113_47.n17 a_113_47.n14 20.723
R167 a_113_47.n6 a_113_47.n5 17.527
R168 a_113_47.n16 a_113_47.n15 13.145
R169 a_113_47.n9 a_113_47.n8 5.842
R170 a_113_47.n8 a_113_47.n7 4.381
R171 a_113_47.n12 a_113_47.n11 4.381
R172 a_113_47.n13 a_113_47.n12 1.46
R173 Y.n2 Y.n0 155.184
R174 Y.n8 Y.n7 154.573
R175 Y.n10 Y.n9 146.375
R176 Y.n5 Y.n4 133.853
R177 Y.n2 Y.n1 110.76
R178 Y.n5 Y.n3 92.5
R179 Y.n6 Y.n5 57.371
R180 Y.n10 Y.n8 52.621
R181 Y.n8 Y.n6 35.388
R182 Y.n6 Y.n2 27.105
R183 Y.n9 Y.t2 26.595
R184 Y.n9 Y.t3 26.595
R185 Y.n0 Y.t5 26.595
R186 Y.n0 Y.t4 26.595
R187 Y.n1 Y.t7 26.595
R188 Y.n1 Y.t6 26.595
R189 Y.n7 Y.t0 26.595
R190 Y.n7 Y.t1 26.595
R191 Y.n3 Y.t8 24.923
R192 Y.n3 Y.t10 24.923
R193 Y.n4 Y.t11 24.923
R194 Y.n4 Y.t9 24.923
R195 Y Y.n10 4.228
R196 a_807_47.n10 a_807_47.t3 174.141
R197 a_807_47.n1 a_807_47.t10 128.218
R198 a_807_47.n7 a_807_47.n6 92.5
R199 a_807_47.n9 a_807_47.n8 92.5
R200 a_807_47.n11 a_807_47.n10 92.5
R201 a_807_47.n7 a_807_47.n5 69.223
R202 a_807_47.n1 a_807_47.n0 52.624
R203 a_807_47.n3 a_807_47.n2 52.624
R204 a_807_47.n5 a_807_47.n4 52.624
R205 a_807_47.n10 a_807_47.n9 48.872
R206 a_807_47.n3 a_807_47.n1 36.266
R207 a_807_47.n5 a_807_47.n3 36.266
R208 a_807_47.n9 a_807_47.n7 28.509
R209 a_807_47.n6 a_807_47.t6 24.923
R210 a_807_47.n8 a_807_47.t2 24.923
R211 a_807_47.n4 a_807_47.t7 24.923
R212 a_807_47.n4 a_807_47.t0 24.923
R213 a_807_47.n0 a_807_47.t8 24.923
R214 a_807_47.n0 a_807_47.t11 24.923
R215 a_807_47.n2 a_807_47.t9 24.923
R216 a_807_47.n2 a_807_47.t1 24.923
R217 a_807_47.n11 a_807_47.t4 24.923
R218 a_807_47.t5 a_807_47.n11 24.923
R219 VNB VNB.t9 6223.14
R220 VNB.t18 VNB.t3 4545.05
R221 VNB.t2 VNB.t6 4400
R222 VNB.t13 VNB.t15 2030.77
R223 VNB.t16 VNB.t13 2030.77
R224 VNB.t14 VNB.t16 2030.77
R225 VNB.t1 VNB.t14 2030.77
R226 VNB.t7 VNB.t1 2030.77
R227 VNB.t0 VNB.t7 2030.77
R228 VNB.t6 VNB.t0 2030.77
R229 VNB.t4 VNB.t2 2030.77
R230 VNB.t5 VNB.t4 2030.77
R231 VNB.t3 VNB.t5 2030.77
R232 VNB.t12 VNB.t18 2030.77
R233 VNB.t17 VNB.t12 2030.77
R234 VNB.t19 VNB.t17 2030.77
R235 VNB.t8 VNB.t19 2030.77
R236 VNB.t11 VNB.t8 2030.77
R237 VNB.t10 VNB.t11 2030.77
R238 VNB.t9 VNB.t10 2030.77
R239 B2.n0 B2.t2 212.079
R240 B2.n2 B2.t3 212.079
R241 B2.n7 B2.t6 212.079
R242 B2.n5 B2.t7 212.079
R243 B2.n0 B2.t5 139.779
R244 B2.n2 B2.t1 139.779
R245 B2.n7 B2.t4 139.779
R246 B2.n5 B2.t0 139.779
R247 B2.n9 B2.n6 96.723
R248 B2.n4 B2.n1 96.723
R249 B2.n4 B2.n3 76
R250 B2.n9 B2.n8 76
R251 B2.n1 B2.n0 21.909
R252 B2 B2.n4 16.152
R253 B2.n6 B2.n5 13.145
R254 B2.n3 B2.n2 10.224
R255 B2 B2.n9 4.571
R256 B2.n8 B2.n7 1.46
R257 VGND.n3 VGND.n0 125.514
R258 VGND.n7 VGND.n6 115.464
R259 VGND.n2 VGND.n1 115.464
R260 VGND.n12 VGND.n11 115.464
R261 VGND.n30 VGND.n29 115.464
R262 VGND.n34 VGND.n33 115.464
R263 VGND.n6 VGND.t0 24.923
R264 VGND.n6 VGND.t2 24.923
R265 VGND.n0 VGND.t7 24.923
R266 VGND.n0 VGND.t5 24.923
R267 VGND.n1 VGND.t8 24.923
R268 VGND.n1 VGND.t6 24.923
R269 VGND.n11 VGND.t1 24.923
R270 VGND.n11 VGND.t3 24.923
R271 VGND.n29 VGND.t10 24.923
R272 VGND.n29 VGND.t4 24.923
R273 VGND.n33 VGND.t9 24.923
R274 VGND.n33 VGND.t11 24.923
R275 VGND.n31 VGND.n30 17.317
R276 VGND.n35 VGND.n34 11.294
R277 VGND.n3 VGND.n2 9.978
R278 VGND.n13 VGND.n12 6.023
R279 VGND.n5 VGND.n4 4.65
R280 VGND.n8 VGND.n7 4.65
R281 VGND.n10 VGND.n9 4.65
R282 VGND.n14 VGND.n13 4.65
R283 VGND.n16 VGND.n15 4.65
R284 VGND.n18 VGND.n17 4.65
R285 VGND.n20 VGND.n19 4.65
R286 VGND.n22 VGND.n21 4.65
R287 VGND.n24 VGND.n23 4.65
R288 VGND.n26 VGND.n25 4.65
R289 VGND.n28 VGND.n27 4.65
R290 VGND.n32 VGND.n31 4.65
R291 VGND.n36 VGND.n35 4.65
R292 VGND VGND.n37 0.488
R293 VGND.n5 VGND.n3 0.318
R294 VGND.n37 VGND.n36 0.134
R295 VGND.n8 VGND.n5 0.119
R296 VGND.n10 VGND.n8 0.119
R297 VGND.n14 VGND.n10 0.119
R298 VGND.n16 VGND.n14 0.119
R299 VGND.n18 VGND.n16 0.119
R300 VGND.n20 VGND.n18 0.119
R301 VGND.n22 VGND.n20 0.119
R302 VGND.n24 VGND.n22 0.119
R303 VGND.n26 VGND.n24 0.119
R304 VGND.n28 VGND.n26 0.119
R305 VGND.n32 VGND.n28 0.119
R306 VGND.n36 VGND.n32 0.119
R307 a_27_47.n4 a_27_47.t1 214.229
R308 a_27_47.n1 a_27_47.t6 128.218
R309 a_27_47.n5 a_27_47.n4 92.5
R310 a_27_47.n4 a_27_47.n3 53.163
R311 a_27_47.n1 a_27_47.n0 52.624
R312 a_27_47.n3 a_27_47.n1 48.574
R313 a_27_47.n3 a_27_47.n2 42.273
R314 a_27_47.n2 a_27_47.t7 24.923
R315 a_27_47.n2 a_27_47.t0 24.923
R316 a_27_47.n0 a_27_47.t4 24.923
R317 a_27_47.n0 a_27_47.t5 24.923
R318 a_27_47.t3 a_27_47.n5 24.923
R319 a_27_47.n5 a_27_47.t2 24.923
R320 A1_N.n0 A1_N.t0 212.079
R321 A1_N.n2 A1_N.t3 212.079
R322 A1_N.n7 A1_N.t6 212.079
R323 A1_N.n5 A1_N.t7 212.079
R324 A1_N.n0 A1_N.t2 139.779
R325 A1_N.n2 A1_N.t5 139.779
R326 A1_N.n7 A1_N.t1 139.779
R327 A1_N.n5 A1_N.t4 139.779
R328 A1_N.n9 A1_N.n6 96.723
R329 A1_N.n4 A1_N.n1 96.723
R330 A1_N.n4 A1_N.n3 76
R331 A1_N.n9 A1_N.n8 76
R332 A1_N.n1 A1_N.n0 21.909
R333 A1_N A1_N.n9 17.98
R334 A1_N.n6 A1_N.n5 13.145
R335 A1_N.n3 A1_N.n2 10.224
R336 A1_N A1_N.n4 2.742
R337 A1_N.n8 A1_N.n7 1.46
C0 VPWR Y 0.70fF
C1 VPB VPWR 0.20fF
C2 VPWR VGND 0.22fF
C3 B2 Y 0.24fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__o21a_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__o21a_1 X A1 B1 A2 VGND VPWR VNB VPB
X0 VPWR.t0 A1.t0 a_382_297.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_297_47.t1 B1.t0 a_79_21.t0 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 a_297_47.t0 A1.t1 VGND.t0 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 VGND.t1 A2.t0 a_297_47.t2 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 VPWR.t1 a_79_21.t3 X.t1 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 a_79_21.t1 B1.t1 VPWR.t2 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 a_382_297.t1 A2.t1 a_79_21.t2 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 VGND.t2 a_79_21.t4 X.t0 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
R0 A1.n0 A1.t0 226.389
R1 A1.n0 A1.t1 158.274
R2 A1 A1.n0 91.86
R3 a_382_297.t0 a_382_297.t1 60.085
R4 VPWR.n5 VPWR.t0 195.082
R5 VPWR.n3 VPWR.n2 193.648
R6 VPWR.n4 VPWR.n1 180.045
R7 VPWR.n0 VPWR.t1 28.565
R8 VPWR.n2 VPWR.t2 27.58
R9 VPWR.n1 VPWR.n0 22.434
R10 VPWR.n5 VPWR.n4 8.81
R11 VPWR.n4 VPWR.n3 4.058
R12 VPWR VPWR.n5 0.204
R13 VPB.t1 VPB.t3 476.479
R14 VPB.t3 VPB.t2 319.626
R15 VPB.t2 VPB.t0 269.314
R16 VPB VPB.t1 204.205
R17 B1.n0 B1.t1 239.984
R18 B1.n0 B1.t0 167.684
R19 B1 B1.n0 92.973
R20 a_79_21.n0 a_79_21.t3 231.014
R21 a_79_21.n0 a_79_21.t4 158.714
R22 a_79_21.n2 a_79_21.n1 158.35
R23 a_79_21.n1 a_79_21.t0 116.128
R24 a_79_21.n1 a_79_21.n0 76
R25 a_79_21.t1 a_79_21.n2 41.37
R26 a_79_21.n2 a_79_21.t2 35.46
R27 a_297_47.t0 a_297_47.n0 225.987
R28 a_297_47.n0 a_297_47.t1 32.307
R29 a_297_47.n0 a_297_47.t2 24.923
R30 VNB VNB.t3 6078.09
R31 VNB.t3 VNB.t1 4545.05
R32 VNB.t1 VNB.t2 2224.18
R33 VNB.t2 VNB.t0 2030.77
R34 VGND.n1 VGND.t2 202.111
R35 VGND.n1 VGND.n0 119.396
R36 VGND.n0 VGND.t0 24.923
R37 VGND.n0 VGND.t1 24.923
R38 VGND VGND.n1 0.145
R39 A2.n0 A2.t1 241.534
R40 A2.n0 A2.t0 169.234
R41 A2 A2.n0 81.177
R42 X X.n0 158.036
R43 X.n1 X.t0 126.71
R44 X.n0 X.t1 26.595
R45 X X.n1 7.542
C0 A2 A1 0.12fF
C1 X VPWR 0.14fF
C2 A2 VPWR 0.11fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__o21a_2.ext - technology: sky130A

.subckt sky130_fd_sc_hd__o21a_2 A1 B1 A2 X VGND VPWR VNB VPB
X0 VPWR.t0 A1.t0 a_470_297.t1 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_79_21.t1 B1.t0 VPWR.t1 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 VGND.t2 a_79_21.t3 X.t3 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 VGND.t0 A2.t0 a_384_47.t1 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 a_470_297.t0 A2.t1 a_79_21.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 VPWR.t2 a_79_21.t4 X.t1 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 a_384_47.t2 B1.t1 a_79_21.t2 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 a_384_47.t0 A1.t1 VGND.t3 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 X.t0 a_79_21.t5 VPWR.t3 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 X.t2 a_79_21.t6 VGND.t1 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
R0 A1.n0 A1.t0 230.154
R1 A1.n0 A1.t1 157.854
R2 A1 A1.n0 78.109
R3 a_470_297.t0 a_470_297.t1 63.04
R4 VPWR.n6 VPWR.n5 292.5
R5 VPWR.n2 VPWR.n1 292.5
R6 VPWR.n11 VPWR.t3 268.15
R7 VPWR.n0 VPWR.t0 258.304
R8 VPWR.n1 VPWR.t1 27.58
R9 VPWR.n5 VPWR.t2 27.58
R10 VPWR.n4 VPWR.n3 4.65
R11 VPWR.n8 VPWR.n7 4.65
R12 VPWR.n10 VPWR.n9 4.65
R13 VPWR.n12 VPWR.n11 4.65
R14 VPWR.n7 VPWR.n6 0.825
R15 VPWR.n3 VPWR.n2 0.412
R16 VPWR.n4 VPWR.n0 0.213
R17 VPWR.n8 VPWR.n4 0.119
R18 VPWR.n10 VPWR.n8 0.119
R19 VPWR.n12 VPWR.n10 0.119
R20 VPWR VPWR.n12 0.02
R21 VPB.t3 VPB.t2 562.305
R22 VPB.t0 VPB.t1 278.193
R23 VPB.t2 VPB.t0 254.517
R24 VPB.t4 VPB.t3 251.557
R25 VPB VPB.t4 189.408
R26 B1.n0 B1.t0 232.213
R27 B1.n0 B1.t1 159.913
R28 B1 B1.n0 84.897
R29 a_79_21.n3 a_79_21.n2 237.955
R30 a_79_21.n1 a_79_21.t4 208.866
R31 a_79_21.n0 a_79_21.t5 208.866
R32 a_79_21.n1 a_79_21.t3 139.779
R33 a_79_21.n0 a_79_21.t6 139.779
R34 a_79_21.n2 a_79_21.t2 116.549
R35 a_79_21.n2 a_79_21.n1 107.08
R36 a_79_21.n1 a_79_21.n0 60.25
R37 a_79_21.t0 a_79_21.n3 27.58
R38 a_79_21.n3 a_79_21.t1 27.58
R39 X.n2 X.n0 173.004
R40 X.n2 X.n1 144.498
R41 X.n1 X.t1 27.58
R42 X.n1 X.t0 26.595
R43 X.n0 X.t3 25.846
R44 X.n0 X.t2 24.923
R45 X X.n2 8.13
R46 VGND.n1 VGND.t2 188.748
R47 VGND.n2 VGND.n0 110.98
R48 VGND.n5 VGND.t1 110.226
R49 VGND.n0 VGND.t3 29.538
R50 VGND.n0 VGND.t0 29.538
R51 VGND.n6 VGND.n5 4.65
R52 VGND.n4 VGND.n3 4.65
R53 VGND.n2 VGND.n1 3.99
R54 VGND.n4 VGND.n2 0.147
R55 VGND.n6 VGND.n4 0.119
R56 VGND VGND.n6 0.02
R57 VNB VNB.t1 6053.91
R58 VNB.t2 VNB.t4 4593.41
R59 VNB.t0 VNB.t3 2272.53
R60 VNB.t4 VNB.t0 2079.12
R61 VNB.t1 VNB.t2 2054.95
R62 A2.n0 A2.t1 236.179
R63 A2.n0 A2.t0 163.879
R64 A2 A2.n0 105.29
R65 a_384_47.t0 a_384_47.n0 264.53
R66 a_384_47.n0 a_384_47.t1 25.846
R67 a_384_47.n0 a_384_47.t2 25.846
C0 X VGND 0.14fF
C1 VPWR X 0.16fF
C2 B1 A2 0.13fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__o21a_4.ext - technology: sky130A

.subckt sky130_fd_sc_hd__o21a_4 A1 A2 B1 X VPWR VGND VNB VPB
X0 X.t3 a_80_21.t6 VGND.t7 VNB.t8 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 a_475_47.t1 A1.t0 VGND.t1 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 X.t7 a_80_21.t7 VPWR.t5 VPB.t7 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 VGND.t6 a_80_21.t8 X.t2 VNB.t7 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 a_762_297.t0 A1.t1 VPWR.t0 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 a_475_47.t2 B1.t0 a_80_21.t0 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 VGND.t2 A2.t0 a_475_47.t3 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 VGND.t5 a_80_21.t9 X.t1 VNB.t6 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 VPWR.t4 a_80_21.t10 X.t6 VPB.t6 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 X.t0 a_80_21.t11 VGND.t4 VNB.t5 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 a_80_21.t1 A2.t1 a_762_297.t1 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 a_80_21.t3 B1.t1 a_475_47.t5 VNB.t9 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 a_80_21.t4 B1.t2 VPWR.t6 VPB.t8 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13 a_475_47.t4 A2.t2 VGND.t3 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14 X.t5 a_80_21.t12 VPWR.t3 VPB.t5 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 VPWR.t1 A1.t2 a_934_297.t1 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16 a_934_297.t0 A2.t3 a_80_21.t2 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17 VPWR.t7 B1.t3 a_80_21.t5 VPB.t9 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X18 VPWR.t2 a_80_21.t13 X.t4 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X19 VGND.t0 A1.t3 a_475_47.t0 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
R0 a_80_21.n18 a_80_21.n17 227.922
R1 a_80_21.n13 a_80_21.t13 225.224
R2 a_80_21.n11 a_80_21.t12 212.079
R3 a_80_21.n7 a_80_21.t10 212.079
R4 a_80_21.n2 a_80_21.t7 212.079
R5 a_80_21.n1 a_80_21.t11 163.148
R6 a_80_21.n17 a_80_21.n16 150.789
R7 a_80_21.n15 a_80_21.n0 143.067
R8 a_80_21.n3 a_80_21.t9 139.779
R9 a_80_21.n6 a_80_21.t6 139.779
R10 a_80_21.n10 a_80_21.t8 139.779
R11 a_80_21.n5 a_80_21.n1 88.8
R12 a_80_21.n12 a_80_21.n11 76
R13 a_80_21.n9 a_80_21.n8 76
R14 a_80_21.n5 a_80_21.n4 76
R15 a_80_21.n14 a_80_21.n13 76
R16 a_80_21.n17 a_80_21.n15 56.679
R17 a_80_21.n16 a_80_21.t5 27.58
R18 a_80_21.n16 a_80_21.t4 27.58
R19 a_80_21.n18 a_80_21.t2 27.58
R20 a_80_21.t1 a_80_21.n18 27.58
R21 a_80_21.n0 a_80_21.t0 25.846
R22 a_80_21.n0 a_80_21.t3 25.846
R23 a_80_21.n11 a_80_21.n10 16.066
R24 a_80_21.n3 a_80_21.n2 16.066
R25 a_80_21.n8 a_80_21.n7 13.145
R26 a_80_21.n14 a_80_21.n12 12.8
R27 a_80_21.n12 a_80_21.n9 12.8
R28 a_80_21.n9 a_80_21.n5 12.8
R29 a_80_21.n4 a_80_21.n3 10.224
R30 a_80_21.n15 a_80_21.n14 8.282
R31 a_80_21.n8 a_80_21.n6 2.921
R32 VGND.n10 VGND.t6 188.748
R33 VGND.n19 VGND.t4 188.748
R34 VGND.n3 VGND.n0 109.976
R35 VGND.n15 VGND.n14 106.463
R36 VGND.n2 VGND.n1 106.052
R37 VGND.n1 VGND.t0 38.769
R38 VGND.n1 VGND.t3 27.692
R39 VGND.n0 VGND.t1 25.846
R40 VGND.n0 VGND.t2 25.846
R41 VGND.n14 VGND.t7 25.846
R42 VGND.n14 VGND.t5 25.846
R43 VGND.n20 VGND.n19 4.65
R44 VGND.n5 VGND.n4 4.65
R45 VGND.n7 VGND.n6 4.65
R46 VGND.n9 VGND.n8 4.65
R47 VGND.n11 VGND.n10 4.65
R48 VGND.n13 VGND.n12 4.65
R49 VGND.n16 VGND.n15 4.65
R50 VGND.n18 VGND.n17 4.65
R51 VGND.n3 VGND.n2 3.747
R52 VGND.n5 VGND.n3 0.248
R53 VGND.n7 VGND.n5 0.119
R54 VGND.n9 VGND.n7 0.119
R55 VGND.n11 VGND.n9 0.119
R56 VGND.n13 VGND.n11 0.119
R57 VGND.n16 VGND.n13 0.119
R58 VGND.n18 VGND.n16 0.119
R59 VGND.n20 VGND.n18 0.119
R60 VGND VGND.n20 0.02
R61 X.n2 X.n0 220.443
R62 X.n2 X.n1 168.766
R63 X.n5 X.n3 150.436
R64 X.n5 X.n4 92.5
R65 X X.n2 92.104
R66 X X.n5 29.609
R67 X.n0 X.t4 27.58
R68 X.n0 X.t5 27.58
R69 X.n1 X.t6 27.58
R70 X.n1 X.t7 27.58
R71 X.n4 X.t1 25.846
R72 X.n4 X.t0 25.846
R73 X.n3 X.t2 25.846
R74 X.n3 X.t3 25.846
R75 VNB VNB.t5 6078.09
R76 VNB.t7 VNB.t9 4593.41
R77 VNB.t0 VNB.t4 2465.93
R78 VNB.t2 VNB.t0 2465.93
R79 VNB.t3 VNB.t1 2079.12
R80 VNB.t4 VNB.t3 2079.12
R81 VNB.t9 VNB.t2 2079.12
R82 VNB.t8 VNB.t7 2079.12
R83 VNB.t6 VNB.t8 2079.12
R84 VNB.t5 VNB.t6 2079.12
R85 A1.n1 A1.t2 236.179
R86 A1.n0 A1.t1 233.287
R87 A1 A1.n0 175.712
R88 A1.n1 A1.t0 163.879
R89 A1.n0 A1.t3 160.987
R90 A1 A1.n1 85.859
R91 a_475_47.n2 a_475_47.t5 223.139
R92 a_475_47.t1 a_475_47.n3 183.098
R93 a_475_47.n3 a_475_47.n0 92.5
R94 a_475_47.n3 a_475_47.n2 64.327
R95 a_475_47.n2 a_475_47.n1 43.354
R96 a_475_47.n1 a_475_47.t2 40.615
R97 a_475_47.n0 a_475_47.t3 25.846
R98 a_475_47.n0 a_475_47.t4 25.846
R99 a_475_47.n1 a_475_47.t0 25.846
R100 VPWR.n10 VPWR.n9 306.397
R101 VPWR.n6 VPWR.n5 292.5
R102 VPWR.n2 VPWR.n1 292.5
R103 VPWR.n0 VPWR.t1 193.744
R104 VPWR.n21 VPWR.t5 192.21
R105 VPWR.n16 VPWR.n15 164.63
R106 VPWR.n9 VPWR.t2 31.52
R107 VPWR.n1 VPWR.t0 27.58
R108 VPWR.n5 VPWR.t7 27.58
R109 VPWR.n9 VPWR.t6 27.58
R110 VPWR.n15 VPWR.t3 27.58
R111 VPWR.n15 VPWR.t4 27.58
R112 VPWR.n7 VPWR.n6 5.866
R113 VPWR.n4 VPWR.n3 4.65
R114 VPWR.n8 VPWR.n7 4.65
R115 VPWR.n12 VPWR.n11 4.65
R116 VPWR.n14 VPWR.n13 4.65
R117 VPWR.n18 VPWR.n17 4.65
R118 VPWR.n20 VPWR.n19 4.65
R119 VPWR.n22 VPWR.n21 3.701
R120 VPWR.n11 VPWR.n10 3.388
R121 VPWR.n3 VPWR.n2 1.69
R122 VPWR.n17 VPWR.n16 0.376
R123 VPWR.n22 VPWR.n20 0.143
R124 VPWR.n4 VPWR.n0 0.143
R125 VPWR.n8 VPWR.n4 0.119
R126 VPWR.n12 VPWR.n8 0.119
R127 VPWR.n14 VPWR.n12 0.119
R128 VPWR.n18 VPWR.n14 0.119
R129 VPWR.n20 VPWR.n18 0.119
R130 VPWR VPWR.n22 0.115
R131 VPB.t9 VPB.t1 455.763
R132 VPB VPB.t7 381.775
R133 VPB.t4 VPB.t8 266.355
R134 VPB.t3 VPB.t0 254.517
R135 VPB.t2 VPB.t3 254.517
R136 VPB.t1 VPB.t2 254.517
R137 VPB.t8 VPB.t9 254.517
R138 VPB.t5 VPB.t4 254.517
R139 VPB.t6 VPB.t5 254.517
R140 VPB.t7 VPB.t6 254.517
R141 a_762_297.t0 a_762_297.t1 55.16
R142 B1.n3 B1.t2 228.875
R143 B1.n0 B1.t3 212.079
R144 B1.n1 B1.t0 162.418
R145 B1.n2 B1.t1 139.779
R146 B1 B1.n3 82.637
R147 B1 B1.n1 77.422
R148 B1.n3 B1.n2 9.493
R149 B1.n1 B1.n0 3.651
R150 A2.n0 A2.t3 212.079
R151 A2.n1 A2.t1 212.079
R152 A2.n0 A2.t0 139.779
R153 A2.n1 A2.t2 139.779
R154 A2 A2.n2 31.721
R155 A2.n2 A2.n1 28.046
R156 A2.n2 A2.n0 21.619
R157 a_934_297.t0 a_934_297.t1 55.16
C0 X VGND 0.19fF
C1 A1 A2 0.31fF
C2 VPWR X 0.49fF
C3 VPB VPWR 0.11fF
C4 VPWR VGND 0.12fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__o21ai_0.ext - technology: sky130A

.subckt sky130_fd_sc_hd__o21ai_0 VGND VPWR Y B1 A2 A1 VNB VPB
X0 a_120_369.t0 A1.t0 VPWR.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1 VGND.t1 A1.t1 a_32_47.t1 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 Y.t1 A2.t0 a_120_369.t1 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X3 a_32_47.t0 A2.t1 VGND.t0 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 VPWR.t1 B1.t0 Y.t0 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X5 Y.t2 B1.t1 a_32_47.t2 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
R0 A1.n0 A1.t0 253.565
R1 A1.n0 A1.t1 194.45
R2 A1 A1.n0 32.529
R3 VPWR.n0 VPWR.t0 233.129
R4 VPWR.n0 VPWR.t1 231.529
R5 VPWR VPWR.n0 0.06
R6 a_120_369.t0 a_120_369.t1 73.875
R7 VPB.t2 VPB.t1 254.517
R8 VPB.t0 VPB.t2 230.841
R9 VPB VPB.t0 224.922
R10 a_32_47.n0 a_32_47.t1 301.889
R11 a_32_47.n0 a_32_47.t2 40
R12 a_32_47.t0 a_32_47.n0 40
R13 VGND VGND.n0 110.021
R14 VGND.n0 VGND.t0 40
R15 VGND.n0 VGND.t1 40
R16 VNB VNB.t1 6664.71
R17 VNB.t0 VNB.t2 2782.35
R18 VNB.t1 VNB.t0 2782.35
R19 A2.n0 A2.t0 280.362
R20 A2.n0 A2.t1 219.31
R21 A2 A2.n0 88.533
R22 Y.n1 Y.t2 222.984
R23 Y.n1 Y.n0 146.997
R24 Y.n0 Y.t0 43.093
R25 Y.n0 Y.t1 43.093
R26 Y Y.n1 2.593
R27 B1.n0 B1.t1 309.516
R28 B1.n0 B1.t0 171.342
R29 B1 B1.n0 78.909
C0 VPWR Y 0.20fF
C1 A1 A2 0.13fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__o21ai_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__o21ai_1 VGND VPWR A2 A1 B1 Y VNB VPB
X0 Y.t2 A2.t0 a_109_297.t1 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 VPWR.t1 B1.t0 Y.t0 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=700000u l=150000u
X2 a_27_47.t1 A2.t1 VGND.t1 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 Y.t1 B1.t1 a_27_47.t2 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 a_109_297.t0 A1.t0 VPWR.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 VGND.t0 A1.t1 a_27_47.t0 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
R0 A2.n0 A2.t0 240.482
R1 A2.n0 A2.t1 168.182
R2 A2.n1 A2.n0 83.951
R3 A2 A2.n1 7.876
R4 A2.n1 A2 2.909
R5 a_109_297.t0 a_109_297.t1 41.37
R6 Y Y.t1 212.743
R7 Y.n1 Y.n0 147.104
R8 Y.n0 Y.t2 56.901
R9 Y.n0 Y.t0 46.435
R10 Y Y.n1 10.71
R11 Y.n1 Y 2.439
R12 VPB.t2 VPB.t1 319.626
R13 VPB.t0 VPB.t2 213.084
R14 VPB VPB.t0 189.408
R15 B1.n0 B1.t1 254.254
R16 B1.n0 B1.t0 181.954
R17 B1 B1.n0 78.666
R18 VPWR.n0 VPWR.t1 211.785
R19 VPWR.n0 VPWR.t0 150.438
R20 VPWR VPWR.n0 0.051
R21 VGND VGND.n0 110.006
R22 VGND.n0 VGND.t0 36
R23 VGND.n0 VGND.t1 24.923
R24 a_27_47.t0 a_27_47.n0 286.69
R25 a_27_47.n0 a_27_47.t2 24.923
R26 a_27_47.n0 a_27_47.t1 24.923
R27 VNB VNB.t0 6053.91
R28 VNB.t0 VNB.t1 2320.88
R29 VNB.t1 VNB.t2 2030.77
R30 A1.n0 A1.t0 234.481
R31 A1.n0 A1.t1 162.181
R32 A1 A1.n0 82.787
C0 A1 A2 0.11fF
C1 A2 Y 0.20fF
C2 VPWR Y 0.16fF
C3 A2 VPWR 0.11fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__o21ai_2.ext - technology: sky130A

.subckt sky130_fd_sc_hd__o21ai_2 B1 Y A2 A1 VGND VPWR VNB VPB
X0 VGND.t3 A2.t0 a_29_47.t3 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 Y.t1 B1.t0 a_29_47.t4 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 VPWR.t3 B1.t1 Y.t3 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 VPWR.t0 A1.t0 a_112_297.t1 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 a_29_47.t2 A2.t1 VGND.t2 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 Y.t5 A2.t2 a_112_297.t3 VPB.t5 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 VGND.t0 A1.t1 a_29_47.t0 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 a_112_297.t0 A1.t2 VPWR.t1 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 a_112_297.t2 A2.t3 Y.t4 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 a_29_47.t5 B1.t2 Y.t0 VNB.t5 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 Y.t2 B1.t3 VPWR.t2 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 a_29_47.t1 A1.t3 VGND.t1 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
R0 A2.n0 A2.t3 212.079
R1 A2.n1 A2.t2 212.079
R2 A2.n0 A2.t0 139.779
R3 A2.n1 A2.t1 139.779
R4 A2 A2.n2 34.319
R5 A2.n2 A2.n0 33.093
R6 A2.n2 A2.n1 19.048
R7 a_29_47.n1 a_29_47.t5 173.697
R8 a_29_47.t0 a_29_47.n3 130.258
R9 a_29_47.n3 a_29_47.n1 56.67
R10 a_29_47.n3 a_29_47.n2 51.655
R11 a_29_47.n1 a_29_47.n0 43.173
R12 a_29_47.n0 a_29_47.t4 25.846
R13 a_29_47.n0 a_29_47.t1 25.846
R14 a_29_47.n2 a_29_47.t3 25.846
R15 a_29_47.n2 a_29_47.t2 25.846
R16 VGND.n2 VGND.n1 118.986
R17 VGND.n2 VGND.n0 118.624
R18 VGND.n0 VGND.t1 36.923
R19 VGND.n0 VGND.t3 35.076
R20 VGND.n1 VGND.t2 25.846
R21 VGND.n1 VGND.t0 25.846
R22 VGND VGND.n2 0.197
R23 VNB VNB.t0 6174.79
R24 VNB.t3 VNB.t1 2610.99
R25 VNB.t4 VNB.t5 2079.12
R26 VNB.t1 VNB.t4 2079.12
R27 VNB.t2 VNB.t3 2079.12
R28 VNB.t0 VNB.t2 2079.12
R29 B1.n2 B1.t1 265.099
R30 B1.n0 B1.t3 263.492
R31 B1.n1 B1.t2 160.666
R32 B1.n0 B1.t0 128.533
R33 B1 B1.n2 99.412
R34 B1.n1 B1.n0 83.468
R35 B1.n2 B1.n1 32.133
R36 Y.n3 Y.n0 304.21
R37 Y.n2 Y.n0 292.5
R38 Y.n5 Y.n4 292.5
R39 Y.n2 Y.n1 145.528
R40 Y Y.n3 30.577
R41 Y.n4 Y.t4 27.58
R42 Y.n4 Y.t5 27.58
R43 Y.n0 Y.t3 27.58
R44 Y.n0 Y.t2 27.58
R45 Y.n1 Y.t0 25.846
R46 Y.n1 Y.t1 25.846
R47 Y Y.n5 22.211
R48 Y Y.n2 9.447
R49 Y.n3 Y 4.902
R50 Y.n5 Y 2.635
R51 VPWR.n1 VPWR.n0 307.239
R52 VPWR.n2 VPWR.t3 252.488
R53 VPWR.n9 VPWR.t1 192.256
R54 VPWR.n0 VPWR.t2 32.505
R55 VPWR.n0 VPWR.t0 30.535
R56 VPWR.n4 VPWR.n3 4.65
R57 VPWR.n6 VPWR.n5 4.65
R58 VPWR.n8 VPWR.n7 4.65
R59 VPWR.n10 VPWR.n9 4.65
R60 VPWR.n2 VPWR.n1 3.815
R61 VPWR.n4 VPWR.n2 0.247
R62 VPWR.n6 VPWR.n4 0.119
R63 VPWR.n8 VPWR.n6 0.119
R64 VPWR.n10 VPWR.n8 0.119
R65 VPWR VPWR.n10 0.023
R66 VPB.t4 VPB.t0 295.95
R67 VPB.t0 VPB.t2 278.193
R68 VPB.t2 VPB.t3 254.517
R69 VPB.t5 VPB.t4 254.517
R70 VPB.t1 VPB.t5 254.517
R71 VPB VPB.t1 204.205
R72 A1.n0 A1.t0 236.179
R73 A1.n1 A1.t2 234.39
R74 A1 A1.n0 175.451
R75 A1.n0 A1.t3 163.879
R76 A1.n1 A1.t1 150.442
R77 A1.n2 A1.n1 76
R78 A1.n2 A1 11.054
R79 A1 A1.n2 2.133
R80 a_112_297.n1 a_112_297.n0 504.326
R81 a_112_297.n1 a_112_297.t2 37.43
R82 a_112_297.t1 a_112_297.n1 31.52
R83 a_112_297.n0 a_112_297.t3 27.58
R84 a_112_297.n0 a_112_297.t0 27.58
C0 VPWR Y 0.28fF
C1 A1 Y 0.22fF
C2 A1 A2 0.37fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__o21ai_4.ext - technology: sky130A

.subckt sky130_fd_sc_hd__o21ai_4 Y B1 A2 A1 VPWR VGND VNB VPB
X0 VPWR.t7 B1.t0 Y.t7 VPB.t11 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_115_297.t3 A1.t0 VPWR.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 a_115_297.t4 A2.t0 Y.t0 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 VPWR.t1 A1.t1 a_115_297.t2 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 VGND.t7 A2.t1 a_32_47.t7 VNB.t7 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 Y.t11 B1.t1 a_32_47.t11 VNB.t11 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 VGND.t3 A1.t2 a_32_47.t3 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 Y.t6 B1.t2 VPWR.t6 VPB.t10 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 a_32_47.t10 B1.t3 Y.t10 VNB.t10 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 Y.t9 B1.t4 a_32_47.t9 VNB.t9 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 Y.t1 A2.t2 a_115_297.t5 VPB.t5 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 a_32_47.t6 A2.t3 VGND.t6 VNB.t6 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 a_32_47.t8 B1.t5 Y.t8 VNB.t8 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 a_32_47.t5 A2.t4 VGND.t5 VNB.t5 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14 a_115_297.t6 A2.t5 Y.t2 VPB.t6 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 a_32_47.t2 A1.t3 VGND.t2 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X16 VPWR.t5 B1.t6 Y.t5 VPB.t9 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17 a_32_47.t1 A1.t4 VGND.t1 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X18 VGND.t4 A2.t6 a_32_47.t4 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X19 Y.t4 B1.t7 VPWR.t4 VPB.t8 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X20 VPWR.t2 A1.t5 a_115_297.t1 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X21 Y.t3 A2.t7 a_115_297.t7 VPB.t7 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X22 VGND.t0 A1.t6 a_32_47.t0 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X23 a_115_297.t0 A1.t7 VPWR.t3 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
R0 B1.n5 B1.t0 212.079
R1 B1.n0 B1.t6 212.079
R2 B1.n2 B1.t2 212.079
R3 B1.n7 B1.t7 212.079
R4 B1.n5 B1.t5 139.779
R5 B1.n0 B1.t3 139.779
R6 B1.n2 B1.t1 139.779
R7 B1.n7 B1.t4 139.779
R8 B1.n4 B1.n1 92.738
R9 B1 B1.n8 86.584
R10 B1.n4 B1.n3 76
R11 B1.n6 B1.n5 76
R12 B1.n1 B1.n0 26.29
R13 B1.n6 B1.n4 16.738
R14 B1.n3 B1.n2 13.145
R15 B1.n8 B1.n7 13.145
R16 B1 B1.n6 6.153
R17 Y.n3 Y.n2 357.252
R18 Y.n3 Y.n1 292.5
R19 Y.n6 Y.n0 149.784
R20 Y.n5 Y.n4 149.405
R21 Y.n9 Y.n8 140.36
R22 Y.n5 Y.n3 100.863
R23 Y.n9 Y.n7 92.5
R24 Y Y.n6 40.834
R25 Y.n0 Y.t5 27.58
R26 Y.n0 Y.t6 27.58
R27 Y.n2 Y.t2 27.58
R28 Y.n2 Y.t1 27.58
R29 Y.n1 Y.t0 27.58
R30 Y.n1 Y.t3 27.58
R31 Y.n4 Y.t7 27.58
R32 Y.n4 Y.t4 27.58
R33 Y.n7 Y.t10 25.846
R34 Y.n7 Y.t11 25.846
R35 Y.n8 Y.t8 25.846
R36 Y.n8 Y.t9 25.846
R37 Y Y.n9 21.683
R38 Y.n6 Y.n5 17.298
R39 VPWR.n6 VPWR.n5 308.957
R40 VPWR.n19 VPWR.n18 307.239
R41 VPWR.n1 VPWR.n0 307.239
R42 VPWR.n2 VPWR.t5 196.104
R43 VPWR.n23 VPWR.t3 194.617
R44 VPWR.n5 VPWR.t4 31.52
R45 VPWR.n5 VPWR.t1 31.52
R46 VPWR.n18 VPWR.t0 27.58
R47 VPWR.n18 VPWR.t2 27.58
R48 VPWR.n0 VPWR.t6 27.58
R49 VPWR.n0 VPWR.t7 27.58
R50 VPWR.n2 VPWR.n1 6.822
R51 VPWR.n4 VPWR.n3 4.65
R52 VPWR.n7 VPWR.n6 4.65
R53 VPWR.n9 VPWR.n8 4.65
R54 VPWR.n11 VPWR.n10 4.65
R55 VPWR.n13 VPWR.n12 4.65
R56 VPWR.n15 VPWR.n14 4.65
R57 VPWR.n17 VPWR.n16 4.65
R58 VPWR.n20 VPWR.n19 4.65
R59 VPWR.n22 VPWR.n21 4.65
R60 VPWR.n24 VPWR.n23 4.65
R61 VPWR.n4 VPWR.n2 0.455
R62 VPWR.n7 VPWR.n4 0.119
R63 VPWR.n9 VPWR.n7 0.119
R64 VPWR.n11 VPWR.n9 0.119
R65 VPWR.n13 VPWR.n11 0.119
R66 VPWR.n15 VPWR.n13 0.119
R67 VPWR.n17 VPWR.n15 0.119
R68 VPWR.n20 VPWR.n17 0.119
R69 VPWR.n22 VPWR.n20 0.119
R70 VPWR.n24 VPWR.n22 0.119
R71 VPWR VPWR.n24 0.022
R72 VPB.t1 VPB.t8 278.193
R73 VPB.t10 VPB.t9 254.517
R74 VPB.t11 VPB.t10 254.517
R75 VPB.t8 VPB.t11 254.517
R76 VPB.t4 VPB.t1 254.517
R77 VPB.t7 VPB.t4 254.517
R78 VPB.t6 VPB.t7 254.517
R79 VPB.t5 VPB.t6 254.517
R80 VPB.t0 VPB.t5 254.517
R81 VPB.t2 VPB.t0 254.517
R82 VPB.t3 VPB.t2 254.517
R83 VPB VPB.t3 210.124
R84 A1.n3 A1.n0 250.009
R85 A1.n0 A1.t1 236.179
R86 A1.n1 A1.t0 212.079
R87 A1.n6 A1.t5 212.079
R88 A1.n4 A1.t7 212.079
R89 A1.n0 A1.t3 163.879
R90 A1.n1 A1.t6 139.779
R91 A1.n6 A1.t4 139.779
R92 A1.n4 A1.t2 139.779
R93 A1.n3 A1.n2 76
R94 A1.n8 A1.n7 76
R95 A1.n8 A1.n5 48.867
R96 A1.n5 A1.n4 10.586
R97 A1.n2 A1.n1 7.303
R98 A1.n7 A1.n6 5.842
R99 A1 A1.n3 4.68
R100 A1 A1.n8 1.814
R101 a_115_297.n4 a_115_297.n0 377.813
R102 a_115_297.n3 a_115_297.n1 350.436
R103 a_115_297.n3 a_115_297.n2 292.5
R104 a_115_297.n5 a_115_297.n4 292.5
R105 a_115_297.n4 a_115_297.n3 57.936
R106 a_115_297.n0 a_115_297.t1 27.58
R107 a_115_297.n0 a_115_297.t0 27.58
R108 a_115_297.n2 a_115_297.t7 27.58
R109 a_115_297.n2 a_115_297.t6 27.58
R110 a_115_297.n1 a_115_297.t2 27.58
R111 a_115_297.n1 a_115_297.t4 27.58
R112 a_115_297.n5 a_115_297.t5 27.58
R113 a_115_297.t3 a_115_297.n5 27.58
R114 A2.n0 A2.t0 212.079
R115 A2.n2 A2.t7 212.079
R116 A2.n5 A2.t5 212.079
R117 A2.n6 A2.t2 212.079
R118 A2.n0 A2.t1 139.779
R119 A2.n2 A2.t3 139.779
R120 A2.n5 A2.t6 139.779
R121 A2.n6 A2.t4 139.779
R122 A2.n4 A2.n1 94.618
R123 A2.n4 A2.n3 76
R124 A2.n8 A2.n7 76
R125 A2.n7 A2.n6 54.042
R126 A2.n8 A2.n4 20.014
R127 A2.n1 A2.n0 13.145
R128 A2.n3 A2.n2 8.763
R129 A2.n7 A2.n5 8.763
R130 A2 A2.n8 8.145
R131 a_32_47.t10 a_32_47.n9 234.646
R132 a_32_47.n4 a_32_47.t3 172.043
R133 a_32_47.n6 a_32_47.n1 92.5
R134 a_32_47.n5 a_32_47.n2 92.5
R135 a_32_47.n4 a_32_47.n3 92.5
R136 a_32_47.n8 a_32_47.n7 92.5
R137 a_32_47.n9 a_32_47.n0 92.5
R138 a_32_47.n9 a_32_47.n8 62.109
R139 a_32_47.n8 a_32_47.n6 57.504
R140 a_32_47.n6 a_32_47.n5 53.697
R141 a_32_47.n5 a_32_47.n4 53.697
R142 a_32_47.n0 a_32_47.t11 25.846
R143 a_32_47.n0 a_32_47.t8 25.846
R144 a_32_47.n7 a_32_47.t9 25.846
R145 a_32_47.n7 a_32_47.t2 25.846
R146 a_32_47.n3 a_32_47.t0 25.846
R147 a_32_47.n3 a_32_47.t1 25.846
R148 a_32_47.n2 a_32_47.t4 25.846
R149 a_32_47.n2 a_32_47.t5 25.846
R150 a_32_47.n1 a_32_47.t7 25.846
R151 a_32_47.n1 a_32_47.t6 25.846
R152 VGND.n3 VGND.n0 109.739
R153 VGND.n2 VGND.n1 106.463
R154 VGND.n7 VGND.n6 106.463
R155 VGND.n12 VGND.n11 106.463
R156 VGND.n0 VGND.t2 33.23
R157 VGND.n0 VGND.t7 25.846
R158 VGND.n1 VGND.t6 25.846
R159 VGND.n1 VGND.t4 25.846
R160 VGND.n6 VGND.t5 25.846
R161 VGND.n6 VGND.t0 25.846
R162 VGND.n11 VGND.t1 25.846
R163 VGND.n11 VGND.t3 25.846
R164 VGND.n5 VGND.n4 4.65
R165 VGND.n8 VGND.n7 4.65
R166 VGND.n10 VGND.n9 4.65
R167 VGND.n13 VGND.n12 3.989
R168 VGND.n3 VGND.n2 3.936
R169 VGND.n5 VGND.n3 0.26
R170 VGND.n13 VGND.n10 0.136
R171 VGND VGND.n13 0.125
R172 VGND.n8 VGND.n5 0.119
R173 VGND.n10 VGND.n8 0.119
R174 VNB VNB.t3 6223.14
R175 VNB.t7 VNB.t2 2272.53
R176 VNB.t11 VNB.t10 2079.12
R177 VNB.t8 VNB.t11 2079.12
R178 VNB.t9 VNB.t8 2079.12
R179 VNB.t2 VNB.t9 2079.12
R180 VNB.t6 VNB.t7 2079.12
R181 VNB.t4 VNB.t6 2079.12
R182 VNB.t5 VNB.t4 2079.12
R183 VNB.t0 VNB.t5 2079.12
R184 VNB.t1 VNB.t0 2079.12
R185 VNB.t3 VNB.t1 2079.12
C0 B1 Y 0.50fF
C1 VPWR Y 0.52fF
C2 A1 Y 0.34fF
C3 A1 A2 0.51fF
C4 VPWR VGND 0.13fF
C5 VPB VPWR 0.12fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__o21ba_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__o21ba_1 B1_N A1 X A2 VGND VPWR VNB VPB
X0 a_222_93.t1 B1_N.t0 VGND.t3 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1 VPWR.t1 A1.t0 a_544_297.t0 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 VGND.t1 a_79_199.t3 X.t1 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 a_222_93.t0 B1_N.t1 VPWR.t3 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 VGND.t2 A2.t0 a_448_47.t1 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 a_448_47.t2 a_222_93.t2 a_79_199.t2 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 a_79_199.t1 a_222_93.t3 VPWR.t2 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 a_544_297.t1 A2.t1 a_79_199.t0 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 a_448_47.t0 A1.t1 VGND.t0 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 VPWR.t0 a_79_199.t4 X.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
R0 B1_N.n0 B1_N.t1 144.547
R1 B1_N.n0 B1_N.t0 128.48
R2 B1_N B1_N.n0 78.715
R3 VGND.n2 VGND.n1 144.432
R4 VGND.n2 VGND.n0 125.505
R5 VGND.n1 VGND.t3 47.142
R6 VGND.n1 VGND.t1 35.428
R7 VGND.n0 VGND.t0 24.923
R8 VGND.n0 VGND.t2 24.923
R9 VGND VGND.n2 0.171
R10 a_222_93.t0 a_222_93.n1 411.161
R11 a_222_93.n0 a_222_93.t3 212.079
R12 a_222_93.n1 a_222_93.t1 184.152
R13 a_222_93.n1 a_222_93.n0 156.333
R14 a_222_93.n0 a_222_93.t2 139.779
R15 VNB VNB.t1 6464.9
R16 VNB.t4 VNB.t3 5463.74
R17 VNB.t1 VNB.t4 2345.05
R18 VNB.t3 VNB.t2 2320.88
R19 VNB.t2 VNB.t0 2030.77
R20 A1.n0 A1.t0 234.801
R21 A1.n0 A1.t1 162.501
R22 A1 A1.n0 91.238
R23 a_544_297.t0 a_544_297.t1 41.37
R24 VPWR.n0 VPWR.t2 515.64
R25 VPWR.n7 VPWR.n6 321.208
R26 VPWR.n1 VPWR.t1 152.253
R27 VPWR.n6 VPWR.t3 114.916
R28 VPWR.n6 VPWR.t0 33.49
R29 VPWR.n3 VPWR.n2 4.65
R30 VPWR.n5 VPWR.n4 4.65
R31 VPWR.n1 VPWR.n0 4.102
R32 VPWR.n8 VPWR.n7 4.05
R33 VPWR.n3 VPWR.n1 0.163
R34 VPWR.n8 VPWR.n5 0.134
R35 VPWR VPWR.n8 0.126
R36 VPWR.n5 VPWR.n3 0.119
R37 VPB.t4 VPB.t3 668.847
R38 VPB.t0 VPB.t4 334.423
R39 VPB.t3 VPB.t2 284.112
R40 VPB.t2 VPB.t1 213.084
R41 VPB VPB.t0 192.367
R42 a_79_199.n0 a_79_199.t4 235.819
R43 a_79_199.n1 a_79_199.t2 190.967
R44 a_79_199.n1 a_79_199.n0 190.267
R45 a_79_199.n0 a_79_199.t3 163.519
R46 a_79_199.n2 a_79_199.n1 97.535
R47 a_79_199.n2 a_79_199.t1 38.415
R48 a_79_199.t0 a_79_199.n2 26.595
R49 X.n0 X.t1 172.272
R50 X.n0 X.t0 121.035
R51 X X.n0 7.611
R52 A2.n0 A2.t1 241.534
R53 A2.n0 A2.t0 169.234
R54 A2 A2.n0 84.533
R55 a_448_47.t0 a_448_47.n0 182.623
R56 a_448_47.n0 a_448_47.t2 36
R57 a_448_47.n0 a_448_47.t1 24.923
.ends

* NGSPICE file created from sky130_fd_sc_hd__o21ba_2.ext - technology: sky130A

.subckt sky130_fd_sc_hd__o21ba_2 B1_N A1 X A2 VGND VPWR VNB VPB
X0 VGND.t1 B1_N.t0 a_27_93.t1 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1 VGND.t0 A2.t0 a_478_47.t1 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 a_478_47.t0 a_27_93.t2 a_174_21.t0 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 a_478_47.t2 A1.t0 VGND.t4 VNB.t5 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 X.t3 a_174_21.t3 VGND.t3 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 VPWR.t4 a_174_21.t4 X.t1 VPB.t5 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 X.t0 a_174_21.t5 VPWR.t3 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 VPWR.t2 A1.t1 a_574_297.t1 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 VGND.t2 a_174_21.t6 X.t2 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 VPWR.t0 B1_N.t1 a_27_93.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10 a_574_297.t0 A2.t1 a_174_21.t2 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 a_174_21.t1 a_27_93.t3 VPWR.t1 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
R0 B1_N.n0 B1_N.t1 148.348
R1 B1_N.n0 B1_N.t0 132.281
R2 B1_N.n1 B1_N.n0 76
R3  B1_N.n1 14.567
R4 B1_N.n1 B1_N 2.011
R5 a_27_93.t0 a_27_93.n1 355.821
R6 a_27_93.n1 a_27_93.n0 318.526
R7 a_27_93.n0 a_27_93.t3 212.079
R8 a_27_93.n1 a_27_93.t1 196.453
R9 a_27_93.n0 a_27_93.t2 139.779
R10 VGND.n1 VGND.t2 189.087
R11 VGND.n6 VGND.n5 139.433
R12 VGND.n2 VGND.n0 120.125
R13 VGND.n5 VGND.t3 41.648
R14 VGND.n5 VGND.t1 38.571
R15 VGND.n0 VGND.t4 24.923
R16 VGND.n0 VGND.t0 24.923
R17 VGND.n4 VGND.n3 4.65
R18 VGND.n7 VGND.n6 4.05
R19 VGND.n2 VGND.n1 3.938
R20 VGND.n4 VGND.n2 0.146
R21 VGND.n7 VGND.n4 0.134
R22 VGND VGND.n7 0.126
R23 VNB VNB.t1 6078.09
R24 VNB.t3 VNB.t2 4593.41
R25 VNB.t2 VNB.t0 2296.7
R26 VNB.t1 VNB.t4 2296.7
R27 VNB.t0 VNB.t5 2030.77
R28 VNB.t4 VNB.t3 2030.77
R29 A2.n0 A2.t1 241.534
R30 A2.n0 A2.t0 169.234
R31 A2 A2.n0 93.676
R32 a_478_47.n0 a_478_47.t2 233.188
R33 a_478_47.t0 a_478_47.n0 35.076
R34 a_478_47.n0 a_478_47.t1 24.923
R35 a_174_21.n2 a_174_21.t4 212.809
R36 a_174_21.n0 a_174_21.t5 212.079
R37 a_174_21.n4 a_174_21.n3 155.917
R38 a_174_21.n0 a_174_21.t3 141.239
R39 a_174_21.n1 a_174_21.t6 139.779
R40 a_174_21.n3 a_174_21.n2 127.818
R41 a_174_21.n3 a_174_21.t0 89.145
R42 a_174_21.n1 a_174_21.n0 59.884
R43 a_174_21.t1 a_174_21.n4 38.415
R44 a_174_21.n4 a_174_21.t2 26.595
R45 a_174_21.n2 a_174_21.n1 0.73
R46 A1.n0 A1.t1 234.801
R47 A1.n0 A1.t0 162.501
R48 A1.n1 A1.n0 76
R49  A1.n1 7.369
R50 A1.n1 A1 1.422
R51 X X.n0 376.28
R52 X X.n1 92.716
R53 X.n0 X.t1 26.595
R54 X.n0 X.t0 26.595
R55 X.n1 X.t2 24.923
R56 X.n1 X.t3 24.923
R57 VPWR.n10 VPWR.n9 308.31
R58 VPWR.n4 VPWR.n3 292.5
R59 VPWR.n1 VPWR.n0 292.5
R60 VPWR.n2 VPWR.t2 196.416
R61 VPWR.n9 VPWR.t0 96.154
R62 VPWR.n0 VPWR.t1 34.475
R63 VPWR.n3 VPWR.t4 30.535
R64 VPWR.n9 VPWR.t3 25.61
R65 VPWR.n6 VPWR.n5 4.65
R66 VPWR.n8 VPWR.n7 4.65
R67 VPWR.n2 VPWR.n1 4.107
R68 VPWR.n11 VPWR.n10 3.941
R69 VPWR.n6 VPWR.n2 0.15
R70 VPWR.n11 VPWR.n8 0.137
R71 VPWR VPWR.n11 0.123
R72 VPWR.n8 VPWR.n6 0.119
R73 VPWR.n5 VPWR.n4 0.106
R74 VPB.t5 VPB.t1 556.386
R75 VPB.t0 VPB.t4 287.071
R76 VPB.t1 VPB.t2 284.112
R77 VPB.t4 VPB.t5 248.598
R78 VPB.t2 VPB.t3 213.084
R79 VPB VPB.t0 192.367
R80 a_574_297.t0 a_574_297.t1 41.37
C0 A2 A1 0.10fF
C1 VGND X 0.17fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__o21ba_4.ext - technology: sky130A

.subckt sky130_fd_sc_hd__o21ba_4 B1_N A1 A2 X VGND VPWR VNB VPB
X0 VPWR.t4 B1_N.t0 a_27_297.t1 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 VPWR.t5 A1.t0 a_743_297.t3 VPB.t7 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 a_743_297.t2 A1.t1 VPWR.t6 VPB.t8 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 a_575_47.t3 a_27_297.t2 a_187_21.t5 VNB.t8 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 a_743_297.t0 A2.t0 a_187_21.t0 VPB.t5 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 VPWR.t8 a_27_297.t3 a_187_21.t3 VPB.t10 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 a_187_21.t1 A2.t1 a_743_297.t1 VPB.t6 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 a_187_21.t2 a_27_297.t4 VPWR.t7 VPB.t9 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 a_187_21.t4 a_27_297.t5 a_575_47.t2 VNB.t7 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 VGND.t4 B1_N.t1 a_27_297.t0 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 VGND.t6 A2.t2 a_575_47.t5 VNB.t10 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 VPWR.t0 a_187_21.t6 X.t3 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 VGND.t8 A1.t2 a_575_47.t1 VNB.t6 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 VGND.t3 a_187_21.t7 X.t7 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14 X.t2 a_187_21.t8 VPWR.t1 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 VPWR.t2 a_187_21.t9 X.t1 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16 a_575_47.t0 A1.t3 VGND.t7 VNB.t5 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X17 a_575_47.t4 A2.t3 VGND.t5 VNB.t9 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X18 X.t0 a_187_21.t10 VPWR.t3 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X19 X.t6 a_187_21.t11 VGND.t2 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X20 X.t5 a_187_21.t12 VGND.t1 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X21 VGND.t0 a_187_21.t13 X.t4 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
R0 B1_N.n0 B1_N.t0 241.534
R1 B1_N.n0 B1_N.t1 169.234
R2 B1_N.n1 B1_N.n0 77.422
R3  B1_N.n1 12.114
R4 B1_N.n1 B1_N 3.428
R5 a_27_297.n3 a_27_297.n2 305.592
R6 a_27_297.n2 a_27_297.t4 252.975
R7 a_27_297.n1 a_27_297.t3 212.079
R8 a_27_297.n0 a_27_297.t2 201.124
R9 a_27_297.n3 a_27_297.t0 144.687
R10 a_27_297.n0 a_27_297.t5 139.779
R11 a_27_297.t1 a_27_297.n3 128.643
R12 a_27_297.n2 a_27_297.n1 20.448
R13 a_27_297.n1 a_27_297.n0 14.606
R14 VPWR.n0 VPWR.t8 552.677
R15 VPWR.n6 VPWR.n5 308.79
R16 VPWR.n11 VPWR.n10 308.79
R17 VPWR.n16 VPWR.n15 308.79
R18 VPWR.n2 VPWR.n1 168.628
R19 VPWR.n1 VPWR.t6 26.595
R20 VPWR.n1 VPWR.t5 26.595
R21 VPWR.n5 VPWR.t7 26.595
R22 VPWR.n5 VPWR.t0 26.595
R23 VPWR.n10 VPWR.t1 26.595
R24 VPWR.n10 VPWR.t2 26.595
R25 VPWR.n15 VPWR.t3 26.595
R26 VPWR.n15 VPWR.t4 26.595
R27 VPWR.n4 VPWR.n3 4.65
R28 VPWR.n7 VPWR.n6 4.65
R29 VPWR.n9 VPWR.n8 4.65
R30 VPWR.n12 VPWR.n11 4.65
R31 VPWR.n14 VPWR.n13 4.65
R32 VPWR.n2 VPWR.n0 4.138
R33 VPWR.n17 VPWR.n16 4.095
R34 VPWR.n4 VPWR.n2 0.136
R35 VPWR.n17 VPWR.n14 0.133
R36 VPWR VPWR.n17 0.127
R37 VPWR.n7 VPWR.n4 0.119
R38 VPWR.n9 VPWR.n7 0.119
R39 VPWR.n12 VPWR.n9 0.119
R40 VPWR.n14 VPWR.n12 0.119
R41 VPB.t10 VPB.t6 556.386
R42 VPB VPB.t4 263.395
R43 VPB.t7 VPB.t8 248.598
R44 VPB.t5 VPB.t7 248.598
R45 VPB.t6 VPB.t5 248.598
R46 VPB.t9 VPB.t10 248.598
R47 VPB.t0 VPB.t9 248.598
R48 VPB.t1 VPB.t0 248.598
R49 VPB.t2 VPB.t1 248.598
R50 VPB.t3 VPB.t2 248.598
R51 VPB.t4 VPB.t3 248.598
R52 A1.n0 A1.t1 212.079
R53 A1.n1 A1.t0 212.079
R54 A1.n0 A1.t3 139.779
R55 A1.n1 A1.t2 139.779
R56 A1 A1.n2 76.777
R57 A1.n2 A1.n1 38.706
R58 A1.n2 A1.n0 22.639
R59 a_743_297.n1 a_743_297.t1 613.707
R60 a_743_297.t2 a_743_297.n1 202.763
R61 a_743_297.n1 a_743_297.n0 87.816
R62 a_743_297.n0 a_743_297.t3 26.595
R63 a_743_297.n0 a_743_297.t0 26.595
R64 a_187_21.n6 a_187_21.t6 212.079
R65 a_187_21.n2 a_187_21.t8 212.079
R66 a_187_21.n4 a_187_21.t9 212.079
R67 a_187_21.n3 a_187_21.t10 212.079
R68 a_187_21.n10 a_187_21.n0 192.066
R69 a_187_21.n11 a_187_21.n10 189.567
R70 a_187_21.n6 a_187_21.t13 139.779
R71 a_187_21.n2 a_187_21.t12 139.779
R72 a_187_21.n4 a_187_21.t7 139.779
R73 a_187_21.n3 a_187_21.t11 139.779
R74 a_187_21.n9 a_187_21.n8 101.631
R75 a_187_21.n8 a_187_21.n5 97.76
R76 a_187_21.n9 a_187_21.n1 92.5
R77 a_187_21.n8 a_187_21.n7 76
R78 a_187_21.n10 a_187_21.n9 69.941
R79 a_187_21.n4 a_187_21.n3 61.345
R80 a_187_21.n5 a_187_21.n4 54.042
R81 a_187_21.n0 a_187_21.t0 26.595
R82 a_187_21.n0 a_187_21.t1 26.595
R83 a_187_21.t3 a_187_21.n11 26.595
R84 a_187_21.n11 a_187_21.t2 26.595
R85 a_187_21.n1 a_187_21.t5 24.923
R86 a_187_21.n1 a_187_21.t4 24.923
R87 a_187_21.n7 a_187_21.n6 18.987
R88 a_187_21.n5 a_187_21.n2 7.303
R89 a_575_47.n2 a_575_47.t2 224.124
R90 a_575_47.n1 a_575_47.t0 124.965
R91 a_575_47.n1 a_575_47.n0 52.624
R92 a_575_47.n2 a_575_47.n1 48.575
R93 a_575_47.n3 a_575_47.n2 42.273
R94 a_575_47.n0 a_575_47.t1 24.923
R95 a_575_47.n0 a_575_47.t4 24.923
R96 a_575_47.n3 a_575_47.t5 24.923
R97 a_575_47.t3 a_575_47.n3 24.923
R98 VNB VNB.t4 6658.31
R99 VNB.t0 VNB.t7 4545.05
R100 VNB.t6 VNB.t5 2030.77
R101 VNB.t9 VNB.t6 2030.77
R102 VNB.t10 VNB.t9 2030.77
R103 VNB.t8 VNB.t10 2030.77
R104 VNB.t7 VNB.t8 2030.77
R105 VNB.t1 VNB.t0 2030.77
R106 VNB.t3 VNB.t1 2030.77
R107 VNB.t2 VNB.t3 2030.77
R108 VNB.t4 VNB.t2 2030.77
R109 A2.n0 A2.t0 212.079
R110 A2.n1 A2.t1 212.079
R111 A2.n0 A2.t3 139.779
R112 A2.n1 A2.t2 139.779
R113 A2 A2.n2 76.676
R114 A2.n2 A2.n0 30.672
R115 A2.n2 A2.n1 30.672
R116 VGND.n10 VGND.t0 193.925
R117 VGND.n3 VGND.n0 125.915
R118 VGND.n2 VGND.n1 115.464
R119 VGND.n16 VGND.n15 115.464
R120 VGND.n22 VGND.n21 74.837
R121 VGND.n0 VGND.t7 24.923
R122 VGND.n0 VGND.t8 24.923
R123 VGND.n1 VGND.t5 24.923
R124 VGND.n1 VGND.t6 24.923
R125 VGND.n15 VGND.t1 24.923
R126 VGND.n15 VGND.t3 24.923
R127 VGND.n21 VGND.t2 24.923
R128 VGND.n21 VGND.t4 24.923
R129 VGND.n23 VGND.n22 12.429
R130 VGND.n3 VGND.n2 12.212
R131 VGND.n5 VGND.n4 4.65
R132 VGND.n7 VGND.n6 4.65
R133 VGND.n9 VGND.n8 4.65
R134 VGND.n12 VGND.n11 4.65
R135 VGND.n14 VGND.n13 4.65
R136 VGND.n18 VGND.n17 4.65
R137 VGND.n20 VGND.n19 4.65
R138 VGND.n11 VGND.n10 3.764
R139 VGND.n17 VGND.n16 2.258
R140 VGND.n5 VGND.n3 0.344
R141 VGND.n23 VGND.n20 0.132
R142 VGND VGND.n23 0.129
R143 VGND.n7 VGND.n5 0.119
R144 VGND.n9 VGND.n7 0.119
R145 VGND.n12 VGND.n9 0.119
R146 VGND.n14 VGND.n12 0.119
R147 VGND.n18 VGND.n14 0.119
R148 VGND.n20 VGND.n18 0.119
R149 X.n2 X.n0 322.284
R150 X.n2 X.n1 293.94
R151 X X.n6 93.857
R152 X.n4 X.n3 52.041
R153 X.n5 X.n4 34.584
R154 X.n1 X.t1 26.595
R155 X.n1 X.t0 26.595
R156 X.n0 X.t3 26.595
R157 X.n0 X.t2 26.595
R158 X.n6 X.t4 24.923
R159 X.n6 X.t5 24.923
R160 X.n3 X.t7 24.923
R161 X.n3 X.t6 24.923
R162 X.n4 X.n2 24.32
R163 X X.n5 11.83
C0 VPWR VGND 0.13fF
C1 VPB VPWR 0.12fF
C2 X VGND 0.43fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__o21bai_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__o21bai_1 A1 Y B1_N A2 VPWR VGND VNB VPB
X0 a_388_297.t1 A2.t0 Y.t2 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_105_352.t0 B1_N.t0 VGND.t1 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 a_297_47.t0 a_105_352.t2 Y.t0 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 a_297_47.t1 A1.t0 VGND.t0 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 VPWR.t1 A1.t1 a_388_297.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 VGND.t2 A2.t1 a_297_47.t2 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 VPWR.t2 B1_N.t1 a_105_352.t1 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7 Y.t1 a_105_352.t3 VPWR.t0 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
R0 A2.n0 A2.t0 241.534
R1 A2.n0 A2.t1 169.234
R2 A2 A2.n0 95.809
R3 Y.n1 Y.t0 210.836
R4 Y.n1 Y.n0 93.995
R5 Y.n0 Y.t1 33.49
R6 Y.n0 Y.t2 26.595
R7 Y Y.n1 8.576
R8 a_388_297.t0 a_388_297.t1 50.235
R9 VPB VPB.t3 423.208
R10 VPB.t3 VPB.t1 325.545
R11 VPB.t1 VPB.t2 269.314
R12 VPB.t2 VPB.t0 239.719
R13 B1_N.n0 B1_N.t1 300.981
R14 B1_N.n0 B1_N.t0 132.281
R15 B1_N B1_N.n0 89.151
R16 VGND.n1 VGND.t1 165.782
R17 VGND.n1 VGND.n0 120.252
R18 VGND.n0 VGND.t0 24.923
R19 VGND.n0 VGND.t2 24.923
R20 VGND VGND.n1 0.042
R21 a_105_352.n1 a_105_352.t1 399.396
R22 a_105_352.n0 a_105_352.t3 212.079
R23 a_105_352.t0 a_105_352.n1 157.842
R24 a_105_352.n1 a_105_352.n0 146.109
R25 a_105_352.n0 a_105_352.t2 139.779
R26 VNB VNB.t2 6078.09
R27 VNB.t2 VNB.t0 4545.05
R28 VNB.t0 VNB.t3 2224.18
R29 VNB.t3 VNB.t1 2030.77
R30 a_297_47.n0 a_297_47.t1 194.913
R31 a_297_47.t0 a_297_47.n0 31.384
R32 a_297_47.n0 a_297_47.t2 25.846
R33 A1.n0 A1.t1 234.801
R34 A1.n0 A1.t0 162.501
R35 A1 A1.n0 79.961
R36 VPWR.n1 VPWR.n0 182.12
R37 VPWR.n1 VPWR.t1 148.696
R38 VPWR.n0 VPWR.t2 101.11
R39 VPWR.n0 VPWR.t0 43.55
R40 VPWR VPWR.n1 0.272
C0 Y VPWR 0.24fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__o21bai_2.ext - technology: sky130A

.subckt sky130_fd_sc_hd__o21bai_2 B1_N Y A2 A1 VGND VPWR VNB VPB
X0 a_397_297.t3 A2.t0 Y.t3 VPB.t5 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 VPWR.t0 B1_N.t0 a_28_297.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 Y.t2 A2.t1 a_397_297.t2 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 VGND.t4 A2.t2 a_229_47.t5 VNB.t6 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 VGND.t2 A1.t0 a_229_47.t3 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 a_28_297.t1 B1_N.t1 VGND.t0 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 Y.t4 a_28_297.t2 a_229_47.t1 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 VPWR.t2 a_28_297.t3 Y.t5 VPB.t6 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 a_397_297.t0 A1.t1 VPWR.t3 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 a_229_47.t0 a_28_297.t4 Y.t0 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 Y.t1 a_28_297.t5 VPWR.t1 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 a_229_47.t4 A2.t3 VGND.t3 VNB.t5 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 a_229_47.t2 A1.t2 VGND.t1 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 VPWR.t4 A1.t3 a_397_297.t1 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
R0 A2.n0 A2.t0 212.079
R1 A2.n1 A2.t1 212.079
R2 A2.n0 A2.t3 139.779
R3 A2.n1 A2.t2 139.779
R4 A2 A2.n2 81.44
R5 A2.n2 A2.n0 30.672
R6 A2.n2 A2.n1 30.672
R7 Y.n2 Y.n1 202.321
R8 Y.n2 Y.n0 137.758
R9 Y Y.n3 126.392
R10 Y.n1 Y.t3 26.595
R11 Y.n1 Y.t2 26.595
R12 Y.n0 Y.t5 26.595
R13 Y.n0 Y.t1 26.595
R14 Y.n3 Y.t0 24.923
R15 Y.n3 Y.t4 24.923
R16 Y Y.n2 4.266
R17 a_397_297.t2 a_397_297.n1 256.512
R18 a_397_297.n1 a_397_297.t0 202.763
R19 a_397_297.n1 a_397_297.n0 87.815
R20 a_397_297.n0 a_397_297.t1 26.595
R21 a_397_297.n0 a_397_297.t3 26.595
R22 VPB.t6 VPB.t4 556.386
R23 VPB.t0 VPB.t1 287.071
R24 VPB.t3 VPB.t2 248.598
R25 VPB.t5 VPB.t3 248.598
R26 VPB.t4 VPB.t5 248.598
R27 VPB.t1 VPB.t6 248.598
R28 VPB VPB.t0 195.327
R29 B1_N.n0 B1_N.t0 140.101
R30 B1_N.n0 B1_N.t1 124.034
R31 B1_N B1_N.n0 84.145
R32 a_28_297.t0 a_28_297.n3 417.937
R33 a_28_297.n2 a_28_297.t5 242.751
R34 a_28_297.n1 a_28_297.t3 212.079
R35 a_28_297.n0 a_28_297.t4 201.124
R36 a_28_297.n3 a_28_297.t1 157.863
R37 a_28_297.n0 a_28_297.t2 139.779
R38 a_28_297.n3 a_28_297.n2 105.364
R39 a_28_297.n2 a_28_297.n1 30.672
R40 a_28_297.n1 a_28_297.n0 14.606
R41 VPWR.n0 VPWR.t2 198.576
R42 VPWR.n2 VPWR.n1 168.03
R43 VPWR.n6 VPWR.n5 167.463
R44 VPWR.n5 VPWR.t0 96.154
R45 VPWR.n1 VPWR.t3 26.595
R46 VPWR.n1 VPWR.t4 26.595
R47 VPWR.n5 VPWR.t1 25.61
R48 VPWR.n4 VPWR.n3 4.65
R49 VPWR.n7 VPWR.n6 4.037
R50 VPWR.n2 VPWR.n0 4.019
R51 VPWR.n4 VPWR.n2 0.138
R52 VPWR.n7 VPWR.n4 0.135
R53 VPWR VPWR.n7 0.126
R54 a_229_47.t1 a_229_47.n3 138.557
R55 a_229_47.n1 a_229_47.t2 124.965
R56 a_229_47.n1 a_229_47.n0 52.624
R57 a_229_47.n3 a_229_47.n1 48.574
R58 a_229_47.n3 a_229_47.n2 42.273
R59 a_229_47.n2 a_229_47.t5 24.923
R60 a_229_47.n2 a_229_47.t0 24.923
R61 a_229_47.n0 a_229_47.t3 24.923
R62 a_229_47.n0 a_229_47.t4 24.923
R63 VGND.n12 VGND.t0 174.365
R64 VGND.n3 VGND.n0 123.286
R65 VGND.n2 VGND.n1 115.464
R66 VGND.n1 VGND.t3 24.923
R67 VGND.n1 VGND.t4 24.923
R68 VGND.n0 VGND.t1 24.923
R69 VGND.n0 VGND.t2 24.923
R70 VGND.n13 VGND.n12 7.285
R71 VGND.n5 VGND.n4 4.65
R72 VGND.n7 VGND.n6 4.65
R73 VGND.n9 VGND.n8 4.65
R74 VGND.n11 VGND.n10 4.65
R75 VGND.n3 VGND.n2 4.024
R76 VGND.n5 VGND.n3 0.25
R77 VGND.n7 VGND.n5 0.119
R78 VGND.n9 VGND.n7 0.119
R79 VGND.n11 VGND.n9 0.119
R80 VGND.n13 VGND.n11 0.119
R81 VGND VGND.n13 0.022
R82 VNB VNB.t0 6102.26
R83 VNB.t0 VNB.t2 4859.34
R84 VNB.t4 VNB.t3 2030.77
R85 VNB.t5 VNB.t4 2030.77
R86 VNB.t6 VNB.t5 2030.77
R87 VNB.t1 VNB.t6 2030.77
R88 VNB.t2 VNB.t1 2030.77
R89 A1.n0 A1.t1 212.079
R90 A1.n1 A1.t3 212.079
R91 A1.n0 A1.t2 139.779
R92 A1.n1 A1.t0 139.779
R93 A1 A1.n2 79.84
R94 A1.n2 A1.n1 38.706
R95 A1.n2 A1.n0 22.639
C0 VPWR Y 0.29fF
C1 A2 Y 0.15fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__o21bai_4.ext - technology: sky130A

.subckt sky130_fd_sc_hd__o21bai_4 Y B1_N A1 A2 VGND VPWR VNB VPB
X0 Y.t3 a_33_297.t2 VPWR.t3 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_225_47.t3 a_33_297.t3 Y.t7 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 VPWR.t2 a_33_297.t4 Y.t2 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 a_33_297.t0 B1_N.t0 VGND.t0 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 Y.t1 a_33_297.t5 VPWR.t1 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 Y.t11 A2.t0 a_561_297.t3 VPB.t10 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 Y.t6 a_33_297.t6 a_225_47.t2 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 Y.t5 a_33_297.t7 a_225_47.t1 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 VGND.t6 A2.t1 a_225_47.t9 VNB.t10 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 VGND.t1 A2.t2 a_225_47.t4 VNB.t5 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 a_561_297.t4 A1.t0 VPWR.t5 VPB.t8 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 a_225_47.t0 a_33_297.t8 Y.t4 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 VPWR.t6 A1.t1 a_561_297.t5 VPB.t9 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13 a_225_47.t7 A1.t2 VGND.t4 VNB.t8 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14 a_225_47.t8 A1.t3 VGND.t5 VNB.t9 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X15 a_225_47.t5 A2.t3 VGND.t2 VNB.t6 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X16 a_225_47.t6 A2.t4 VGND.t3 VNB.t7 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X17 VPWR.t7 A1.t4 a_561_297.t6 VPB.t11 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X18 a_561_297.t7 A1.t5 VPWR.t8 VPB.t12 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X19 VPWR.t4 B1_N.t1 a_33_297.t1 VPB.t7 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X20 a_561_297.t2 A2.t5 Y.t8 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X21 VGND.t7 A1.t6 a_225_47.t10 VNB.t11 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X22 Y.t9 A2.t6 a_561_297.t1 VPB.t5 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X23 VGND.t8 A1.t7 a_225_47.t11 VNB.t12 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X24 a_561_297.t0 A2.t7 Y.t10 VPB.t6 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X25 VPWR.t0 a_33_297.t9 Y.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
R0 a_33_297.n11 a_33_297.t5 225.224
R1 a_33_297.n1 a_33_297.t9 212.079
R2 a_33_297.n4 a_33_297.t2 212.079
R3 a_33_297.n8 a_33_297.t4 212.079
R4 a_33_297.n0 a_33_297.t8 201.124
R5 a_33_297.t1 a_33_297.n13 172.254
R6 a_33_297.n7 a_33_297.t6 139.779
R7 a_33_297.n3 a_33_297.t3 139.779
R8 a_33_297.n0 a_33_297.t7 139.779
R9 a_33_297.n13 a_33_297.t0 108.608
R10 a_33_297.n6 a_33_297.n2 96.723
R11 a_33_297.n12 a_33_297.n11 76
R12 a_33_297.n6 a_33_297.n5 76
R13 a_33_297.n10 a_33_297.n9 76
R14 a_33_297.n2 a_33_297.n1 21.909
R15 a_33_297.n10 a_33_297.n6 20.723
R16 a_33_297.n12 a_33_297.n10 20.723
R17 a_33_297.n1 a_33_297.n0 14.606
R18 a_33_297.n4 a_33_297.n3 14.606
R19 a_33_297.n13 a_33_297.n12 13.409
R20 a_33_297.n9 a_33_297.n7 13.145
R21 a_33_297.n5 a_33_297.n4 10.224
R22 a_33_297.n9 a_33_297.n8 1.46
R23 VPWR.n14 VPWR.t0 198.576
R24 VPWR.n24 VPWR.n23 176.855
R25 VPWR.n1 VPWR.n0 175.109
R26 VPWR.n3 VPWR.n2 171.981
R27 VPWR.n19 VPWR.n18 171.981
R28 VPWR.n0 VPWR.t5 26.595
R29 VPWR.n0 VPWR.t6 26.595
R30 VPWR.n2 VPWR.t8 26.595
R31 VPWR.n2 VPWR.t7 26.595
R32 VPWR.n18 VPWR.t3 26.595
R33 VPWR.n18 VPWR.t2 26.595
R34 VPWR.n23 VPWR.t1 26.595
R35 VPWR.n23 VPWR.t4 26.595
R36 VPWR.n4 VPWR.n3 5.647
R37 VPWR.n5 VPWR.n4 4.65
R38 VPWR.n7 VPWR.n6 4.65
R39 VPWR.n9 VPWR.n8 4.65
R40 VPWR.n11 VPWR.n10 4.65
R41 VPWR.n13 VPWR.n12 4.65
R42 VPWR.n15 VPWR.n14 4.65
R43 VPWR.n17 VPWR.n16 4.65
R44 VPWR.n20 VPWR.n19 4.65
R45 VPWR.n22 VPWR.n21 4.65
R46 VPWR.n25 VPWR.n24 4.105
R47 VPWR.n5 VPWR.n1 0.544
R48 VPWR.n25 VPWR.n22 0.133
R49 VPWR VPWR.n25 0.128
R50 VPWR.n7 VPWR.n5 0.119
R51 VPWR.n9 VPWR.n7 0.119
R52 VPWR.n11 VPWR.n9 0.119
R53 VPWR.n13 VPWR.n11 0.119
R54 VPWR.n15 VPWR.n13 0.119
R55 VPWR.n17 VPWR.n15 0.119
R56 VPWR.n20 VPWR.n17 0.119
R57 VPWR.n22 VPWR.n20 0.119
R58 Y.n2 Y.n0 196.784
R59 Y.n5 Y.n3 157.601
R60 Y.n2 Y.n1 154.829
R61 Y.n9 Y.n7 150.852
R62 Y.n5 Y.n4 110.76
R63 Y.n9 Y.n8 92.5
R64 Y Y.n9 29.724
R65 Y.n3 Y.t2 26.595
R66 Y.n3 Y.t1 26.595
R67 Y.n4 Y.t0 26.595
R68 Y.n4 Y.t3 26.595
R69 Y.n0 Y.t8 26.595
R70 Y.n0 Y.t9 26.595
R71 Y.n1 Y.t10 26.595
R72 Y.n1 Y.t11 26.595
R73 Y.n6 Y.n5 24.989
R74 Y.n7 Y.t7 24.923
R75 Y.n7 Y.t6 24.923
R76 Y.n8 Y.t4 24.923
R77 Y.n8 Y.t5 24.923
R78 Y.n6 Y.n2 23.466
R79 Y Y.n6 2.56
R80 VPB.t0 VPB.t10 556.386
R81 VPB.t9 VPB.t8 248.598
R82 VPB.t12 VPB.t9 248.598
R83 VPB.t11 VPB.t12 248.598
R84 VPB.t4 VPB.t11 248.598
R85 VPB.t5 VPB.t4 248.598
R86 VPB.t6 VPB.t5 248.598
R87 VPB.t10 VPB.t6 248.598
R88 VPB.t3 VPB.t0 248.598
R89 VPB.t2 VPB.t3 248.598
R90 VPB.t1 VPB.t2 248.598
R91 VPB.t7 VPB.t1 248.598
R92 VPB VPB.t7 221.962
R93 a_225_47.n8 a_225_47.t2 234.208
R94 a_225_47.n1 a_225_47.t8 128.218
R95 a_225_47.n9 a_225_47.n8 92.5
R96 a_225_47.n8 a_225_47.n7 64.803
R97 a_225_47.n1 a_225_47.n0 52.624
R98 a_225_47.n3 a_225_47.n2 52.624
R99 a_225_47.n5 a_225_47.n4 52.624
R100 a_225_47.n7 a_225_47.n5 48.574
R101 a_225_47.n7 a_225_47.n6 42.273
R102 a_225_47.n3 a_225_47.n1 36.266
R103 a_225_47.n5 a_225_47.n3 36.266
R104 a_225_47.n6 a_225_47.t9 24.923
R105 a_225_47.n6 a_225_47.t0 24.923
R106 a_225_47.n0 a_225_47.t10 24.923
R107 a_225_47.n0 a_225_47.t7 24.923
R108 a_225_47.n2 a_225_47.t11 24.923
R109 a_225_47.n2 a_225_47.t6 24.923
R110 a_225_47.n4 a_225_47.t4 24.923
R111 a_225_47.n4 a_225_47.t5 24.923
R112 a_225_47.n9 a_225_47.t1 24.923
R113 a_225_47.t3 a_225_47.n9 24.923
R114 VNB VNB.t4 6319.84
R115 VNB.t4 VNB.t2 4545.05
R116 VNB.t11 VNB.t9 2030.77
R117 VNB.t8 VNB.t11 2030.77
R118 VNB.t12 VNB.t8 2030.77
R119 VNB.t7 VNB.t12 2030.77
R120 VNB.t5 VNB.t7 2030.77
R121 VNB.t6 VNB.t5 2030.77
R122 VNB.t10 VNB.t6 2030.77
R123 VNB.t0 VNB.t10 2030.77
R124 VNB.t1 VNB.t0 2030.77
R125 VNB.t3 VNB.t1 2030.77
R126 VNB.t2 VNB.t3 2030.77
R127 B1_N.n0 B1_N.t1 232.736
R128 B1_N.n0 B1_N.t0 160.436
R129 B1_N B1_N.n0 90.933
R130 VGND.n1 VGND.n0 124.367
R131 VGND.n3 VGND.n2 115.464
R132 VGND.n7 VGND.n6 115.464
R133 VGND.n13 VGND.n12 115.464
R134 VGND.n28 VGND.t0 111.584
R135 VGND.n0 VGND.t5 24.923
R136 VGND.n0 VGND.t7 24.923
R137 VGND.n2 VGND.t4 24.923
R138 VGND.n2 VGND.t8 24.923
R139 VGND.n6 VGND.t3 24.923
R140 VGND.n6 VGND.t1 24.923
R141 VGND.n12 VGND.t2 24.923
R142 VGND.n12 VGND.t6 24.923
R143 VGND.n4 VGND.n3 15.058
R144 VGND.n8 VGND.n7 13.552
R145 VGND.n29 VGND.n28 10.673
R146 VGND.n14 VGND.n13 7.529
R147 VGND.n5 VGND.n4 4.65
R148 VGND.n9 VGND.n8 4.65
R149 VGND.n11 VGND.n10 4.65
R150 VGND.n15 VGND.n14 4.65
R151 VGND.n17 VGND.n16 4.65
R152 VGND.n19 VGND.n18 4.65
R153 VGND.n21 VGND.n20 4.65
R154 VGND.n23 VGND.n22 4.65
R155 VGND.n25 VGND.n24 4.65
R156 VGND.n27 VGND.n26 4.65
R157 VGND.n5 VGND.n1 0.473
R158 VGND.n9 VGND.n5 0.119
R159 VGND.n11 VGND.n9 0.119
R160 VGND.n15 VGND.n11 0.119
R161 VGND.n17 VGND.n15 0.119
R162 VGND.n19 VGND.n17 0.119
R163 VGND.n21 VGND.n19 0.119
R164 VGND.n23 VGND.n21 0.119
R165 VGND.n25 VGND.n23 0.119
R166 VGND.n27 VGND.n25 0.119
R167 VGND.n29 VGND.n27 0.119
R168 VGND VGND.n29 0.022
R169 A2.n0 A2.t5 212.079
R170 A2.n2 A2.t6 212.079
R171 A2.n7 A2.t7 212.079
R172 A2.n5 A2.t0 212.079
R173 A2.n0 A2.t4 139.779
R174 A2.n2 A2.t2 139.779
R175 A2.n7 A2.t3 139.779
R176 A2.n5 A2.t1 139.779
R177 A2.n9 A2.n6 97.76
R178 A2.n4 A2.n1 97.76
R179 A2.n4 A2.n3 76
R180 A2.n9 A2.n8 76
R181 A2.n1 A2.n0 21.909
R182 A2 A2.n9 16.32
R183 A2.n6 A2.n5 13.145
R184 A2.n3 A2.n2 10.224
R185 A2 A2.n4 5.44
R186 A2.n8 A2.n7 1.46
R187 a_561_297.t3 a_561_297.n5 224.71
R188 a_561_297.n1 a_561_297.t4 181.779
R189 a_561_297.n5 a_561_297.n4 154.573
R190 a_561_297.n1 a_561_297.n0 110.76
R191 a_561_297.n3 a_561_297.n2 90.234
R192 a_561_297.n5 a_561_297.n3 64.95
R193 a_561_297.n3 a_561_297.n1 64.95
R194 a_561_297.n2 a_561_297.t6 26.595
R195 a_561_297.n2 a_561_297.t2 26.595
R196 a_561_297.n0 a_561_297.t5 26.595
R197 a_561_297.n0 a_561_297.t7 26.595
R198 a_561_297.n4 a_561_297.t1 26.595
R199 a_561_297.n4 a_561_297.t0 26.595
R200 A1.n0 A1.t0 212.079
R201 A1.n1 A1.t1 212.079
R202 A1.n3 A1.t5 212.079
R203 A1.n4 A1.t4 212.079
R204 A1.n0 A1.t3 139.779
R205 A1.n1 A1.t6 139.779
R206 A1.n3 A1.t2 139.779
R207 A1.n4 A1.t7 139.779
R208 A1.n5 A1 95.809
R209 A1.n10 A1.n2 76
R210 A1.n9 A1.n8 76
R211 A1.n7 A1.n6 76
R212 A1.n6 A1.n5 49.66
R213 A1.n2 A1.n1 35.054
R214 A1.n2 A1.n0 26.29
R215 A1.n10 A1.n9 20.723
R216 A1.n9 A1.n7 20.723
R217  A1.n10 13.714
R218 A1.n5 A1.n4 8.763
R219 A1.n6 A1.n3 2.921
R220 A1.n7 A1 0.914
C0 VPWR VGND 0.15fF
C1 A2 Y 0.26fF
C2 VPB VPWR 0.14fF
C3 VPWR Y 0.66fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__o22a_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__o22a_1 A2 X B1 A1 B2 VGND VPWR VNB VPB
X0 a_78_199.t2 B1.t0 a_215_47.t2 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 VPWR.t1 A1.t0 a_493_297.t0 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 a_493_297.t1 A2.t0 a_78_199.t3 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 VPWR.t0 a_78_199.t4 X.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 VGND.t2 A2.t1 a_215_47.t0 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 a_78_199.t0 B2.t0 a_292_297.t0 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 a_215_47.t3 A1.t1 VGND.t1 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 a_215_47.t1 B2.t1 a_78_199.t1 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 a_292_297.t1 B1.t1 VPWR.t2 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 VGND.t0 a_78_199.t5 X.t1 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
R0 B1.n0 B1.t1 1578.82
R1 B1.n0 B1.t0 157.452
R2 B1 B1.n0 81.376
R3 a_215_47.n0 a_215_47.t2 230.998
R4 a_215_47.n0 a_215_47.t3 136.943
R5 a_215_47.n1 a_215_47.n0 43.173
R6 a_215_47.n1 a_215_47.t1 39.692
R7 a_215_47.t0 a_215_47.n1 24.923
R8 a_78_199.n0 a_78_199.t4 230.361
R9 a_78_199.n3 a_78_199.n2 181.088
R10 a_78_199.n2 a_78_199.n1 162.64
R11 a_78_199.n0 a_78_199.t5 158.061
R12 a_78_199.n2 a_78_199.n0 76
R13 a_78_199.n3 a_78_199.t3 65.995
R14 a_78_199.t0 a_78_199.n3 26.595
R15 a_78_199.n1 a_78_199.t1 24.923
R16 a_78_199.n1 a_78_199.t2 24.923
R17 VNB VNB.t1 6078.09
R18 VNB.t1 VNB.t3 4545.05
R19 VNB.t2 VNB.t0 2417.58
R20 VNB.t0 VNB.t4 2030.77
R21 VNB.t3 VNB.t2 2030.77
R22 A1.n0 A1.t0 235.47
R23 A1.n0 A1.t1 163.17
R24 A1 A1.n0 80.48
R25 a_493_297.t0 a_493_297.t1 41.37
R26 VPWR.n0 VPWR.t1 150.774
R27 VPWR.n6 VPWR.n5 146.25
R28 VPWR.n2 VPWR.n1 146.25
R29 VPWR.n5 VPWR.t0 30.535
R30 VPWR.n1 VPWR.t2 26.595
R31 VPWR.n4 VPWR.n3 4.65
R32 VPWR.n7 VPWR.n6 4.442
R33 VPWR.n3 VPWR.n2 0.344
R34 VPWR.n4 VPWR.n0 0.142
R35 VPWR.n7 VPWR.n4 0.135
R36 VPWR VPWR.n7 0.126
R37 VPB.t0 VPB.t3 529.75
R38 VPB.t2 VPB.t4 366.978
R39 VPB.t3 VPB.t2 227.881
R40 VPB.t4 VPB.t1 213.084
R41 VPB VPB.t0 204.205
R42 A2.n0 A2.t0 239.503
R43 A2.n0 A2.t1 167.203
R44 A2 A2.n0 108.406
R45 X.n0 X.t1 176.551
R46 X.n0 X.t0 120.053
R47 X X.n0 9.914
R48 VGND.n1 VGND.t0 202.114
R49 VGND.n1 VGND.n0 118.013
R50 VGND.n0 VGND.t1 24.923
R51 VGND.n0 VGND.t2 24.923
R52 VGND VGND.n1 0.141
R53 B2.n0 B2.t0 241.534
R54 B2.n0 B2.t1 169.234
R55 B2 B2.n0 90.336
R56 a_292_297.t0 a_292_297.t1 46.295
C0 X VPWR 0.14fF
C1 A2 VPWR 0.18fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__o22a_2.ext - technology: sky130A

.subckt sky130_fd_sc_hd__o22a_2 A2 X B1 A1 B2 VGND VPWR VNB VPB
X0 a_301_47.t2 B2.t0 a_81_21.t2 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 VGND.t0 A2.t0 a_301_47.t1 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 a_383_297.t0 B1.t0 VPWR.t2 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 VPWR.t1 a_81_21.t4 X.t1 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 a_301_47.t3 A1.t0 VGND.t3 VNB.t5 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 VGND.t2 a_81_21.t5 X.t3 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 X.t2 a_81_21.t6 VGND.t1 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 X.t0 a_81_21.t7 VPWR.t0 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 VPWR.t3 A1.t1 a_579_297.t1 VPB.t5 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 a_81_21.t0 B1.t1 a_301_47.t0 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 a_579_297.t0 A2.t1 a_81_21.t1 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 a_81_21.t3 B2.t1 a_383_297.t1 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
R0 B2.n0 B2.t1 241.534
R1 B2.n0 B2.t0 169.234
R2 B2 B2.n0 90.336
R3 a_81_21.n2 a_81_21.t4 212.079
R4 a_81_21.n0 a_81_21.t7 212.079
R5 a_81_21.n5 a_81_21.n4 181.332
R6 a_81_21.n4 a_81_21.n3 161.279
R7 a_81_21.n0 a_81_21.t6 141.239
R8 a_81_21.n1 a_81_21.t5 139.779
R9 a_81_21.n4 a_81_21.n2 108.863
R10 a_81_21.t1 a_81_21.n5 65.995
R11 a_81_21.n1 a_81_21.n0 59.884
R12 a_81_21.n5 a_81_21.t3 26.595
R13 a_81_21.n3 a_81_21.t2 24.923
R14 a_81_21.n3 a_81_21.t0 24.923
R15 a_81_21.n2 a_81_21.n1 1.46
R16 a_301_47.t0 a_301_47.n1 231.004
R17 a_301_47.n1 a_301_47.t3 153.014
R18 a_301_47.n1 a_301_47.n0 46.251
R19 a_301_47.n0 a_301_47.t2 40.615
R20 a_301_47.n0 a_301_47.t1 29.538
R21 VNB VNB.t0 6198.96
R22 VNB.t1 VNB.t2 4545.05
R23 VNB.t4 VNB.t3 2562.64
R24 VNB.t3 VNB.t5 2030.77
R25 VNB.t2 VNB.t4 2030.77
R26 VNB.t0 VNB.t1 2030.77
R27 A2.n0 A2.t1 239.503
R28 A2.n0 A2.t0 167.203
R29 A2 A2.n0 107.942
R30 VGND.n1 VGND.t2 202.598
R31 VGND.n2 VGND.n0 117.996
R32 VGND.n5 VGND.t1 113.91
R33 VGND.n0 VGND.t3 24.923
R34 VGND.n0 VGND.t0 24.923
R35 VGND.n6 VGND.n5 7.661
R36 VGND.n4 VGND.n3 4.65
R37 VGND.n2 VGND.n1 4.086
R38 VGND.n4 VGND.n2 0.136
R39 VGND.n6 VGND.n4 0.119
R40 VGND VGND.n6 0.026
R41 B1.n0 B1.t0 230.791
R42 B1.n0 B1.t1 158.491
R43 B1 B1.n0 81.376
R44 VPWR.n0 VPWR.t3 197.193
R45 VPWR.n11 VPWR.t0 154.763
R46 VPWR.n6 VPWR.n5 146.25
R47 VPWR.n2 VPWR.n1 146.25
R48 VPWR.n5 VPWR.t1 34.475
R49 VPWR.n1 VPWR.t2 26.595
R50 VPWR.n4 VPWR.n3 4.65
R51 VPWR.n8 VPWR.n7 4.65
R52 VPWR.n10 VPWR.n9 4.65
R53 VPWR.n12 VPWR.n11 4.65
R54 VPWR.n3 VPWR.n2 0.275
R55 VPWR.n4 VPWR.n0 0.142
R56 VPWR.n7 VPWR.n6 0.137
R57 VPWR.n8 VPWR.n4 0.119
R58 VPWR.n10 VPWR.n8 0.119
R59 VPWR.n12 VPWR.n10 0.119
R60 VPWR VPWR.n12 0.026
R61 a_383_297.t0 a_383_297.t1 41.37
R62 VPB.t2 VPB.t3 550.467
R63 VPB.t4 VPB.t0 366.978
R64 VPB.t1 VPB.t2 248.598
R65 VPB.t0 VPB.t5 213.084
R66 VPB.t3 VPB.t4 213.084
R67 VPB VPB.t1 213.084
R68 X.n2 X.n0 169.28
R69 X.n2 X.n1 92.309
R70 X.n1 X.t1 26.595
R71 X.n1 X.t0 26.595
R72 X.n0 X.t3 24.923
R73 X.n0 X.t2 24.923
R74 X X.n2 12.803
R75 A1.n0 A1.t1 235.47
R76 A1.n0 A1.t0 163.17
R77 A1.n1 A1.n0 76
R78  A1.n1 11.4
R79 A1.n1 A1 2.2
R80 a_579_297.t0 a_579_297.t1 41.37
C0 VPWR VGND 0.11fF
C1 B1 B2 0.11fF
C2 A2 A1 0.14fF
C3 VPWR X 0.25fF
C4 A2 VPWR 0.14fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__o22a_4.ext - technology: sky130A

.subckt sky130_fd_sc_hd__o22a_4 B2 B1 X A1 A2 VGND VPWR VNB VPB
X0 VPWR.t7 B1.t0 a_566_297.t3 VPB.t9 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_484_47.t5 B1.t1 a_96_21.t5 VNB.t9 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 X.t3 a_96_21.t8 VGND.t3 VNB.t5 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 VPWR.t0 a_96_21.t9 X.t7 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 X.t6 a_96_21.t10 VPWR.t1 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 a_566_297.t0 B2.t0 a_96_21.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 VPWR.t2 a_96_21.t11 X.t5 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 X.t2 a_96_21.t12 VGND.t2 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 VGND.t1 a_96_21.t13 X.t1 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 a_96_21.t1 B2.t1 a_566_297.t1 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 VPWR.t4 A1.t0 a_918_297.t3 VPB.t6 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 a_484_47.t2 A1.t1 VGND.t4 VNB.t6 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 a_566_297.t2 B1.t2 VPWR.t6 VPB.t8 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13 a_484_47.t0 B2.t2 a_96_21.t2 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14 a_96_21.t6 A2.t0 a_918_297.t0 VPB.t10 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 a_918_297.t1 A2.t1 a_96_21.t7 VPB.t11 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16 a_484_47.t7 A2.t2 VGND.t7 VNB.t11 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X17 a_918_297.t2 A1.t2 VPWR.t5 VPB.t7 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X18 a_96_21.t4 B1.t3 a_484_47.t4 VNB.t8 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X19 VGND.t6 A2.t3 a_484_47.t6 VNB.t10 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X20 a_96_21.t3 B2.t3 a_484_47.t1 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X21 VGND.t5 A1.t3 a_484_47.t3 VNB.t7 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X22 X.t4 a_96_21.t14 VPWR.t3 VPB.t5 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X23 VGND.t0 a_96_21.t15 X.t0 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
R0 B1.n1 B1.t2 241.534
R1 B1.n0 B1.t0 241.534
R2 B1.n1 B1.t3 169.234
R3 B1.n0 B1.t1 169.234
R4 B1.n2 B1.n0 162.479
R5 B1.n2 B1.n1 76
R6 B1 B1.n2 6.874
R7 a_566_297.n1 a_566_297.n0 638.833
R8 a_566_297.n0 a_566_297.t1 26.595
R9 a_566_297.n0 a_566_297.t2 26.595
R10 a_566_297.n1 a_566_297.t3 26.595
R11 a_566_297.t0 a_566_297.n1 26.595
R12 VPWR.n1 VPWR.n0 308.79
R13 VPWR.n14 VPWR.n13 292.5
R14 VPWR.n10 VPWR.n9 292.5
R15 VPWR.n24 VPWR.t3 197.04
R16 VPWR.n20 VPWR.n19 170.445
R17 VPWR.n2 VPWR.t4 169.602
R18 VPWR.n0 VPWR.t5 42.355
R19 VPWR.n9 VPWR.t6 26.595
R20 VPWR.n13 VPWR.t0 26.595
R21 VPWR.n19 VPWR.t1 26.595
R22 VPWR.n19 VPWR.t2 26.595
R23 VPWR.n0 VPWR.t7 26.595
R24 VPWR.n4 VPWR.n3 4.65
R25 VPWR.n6 VPWR.n5 4.65
R26 VPWR.n8 VPWR.n7 4.65
R27 VPWR.n12 VPWR.n11 4.65
R28 VPWR.n16 VPWR.n15 4.65
R29 VPWR.n18 VPWR.n17 4.65
R30 VPWR.n21 VPWR.n20 4.65
R31 VPWR.n23 VPWR.n22 4.65
R32 VPWR.n25 VPWR.n24 4.65
R33 VPWR.n2 VPWR.n1 4.078
R34 VPWR.n15 VPWR.n14 0.847
R35 VPWR.n11 VPWR.n10 0.282
R36 VPWR.n4 VPWR.n2 0.138
R37 VPWR.n6 VPWR.n4 0.119
R38 VPWR.n8 VPWR.n6 0.119
R39 VPWR.n12 VPWR.n8 0.119
R40 VPWR.n16 VPWR.n12 0.119
R41 VPWR.n18 VPWR.n16 0.119
R42 VPWR.n21 VPWR.n18 0.119
R43 VPWR.n23 VPWR.n21 0.119
R44 VPWR.n25 VPWR.n23 0.119
R45 VPWR VPWR.n25 0.022
R46 VPB.t2 VPB.t8 556.386
R47 VPB.t9 VPB.t7 295.95
R48 VPB.t11 VPB.t6 248.598
R49 VPB.t10 VPB.t11 248.598
R50 VPB.t7 VPB.t10 248.598
R51 VPB.t0 VPB.t9 248.598
R52 VPB.t1 VPB.t0 248.598
R53 VPB.t8 VPB.t1 248.598
R54 VPB.t3 VPB.t2 248.598
R55 VPB.t4 VPB.t3 248.598
R56 VPB.t5 VPB.t4 248.598
R57 VPB VPB.t5 242.679
R58 a_96_21.n16 a_96_21.n0 415.604
R59 a_96_21.n17 a_96_21.n16 292.5
R60 a_96_21.n9 a_96_21.t9 212.079
R61 a_96_21.n6 a_96_21.t10 212.079
R62 a_96_21.n3 a_96_21.t11 212.079
R63 a_96_21.n1 a_96_21.t14 212.079
R64 a_96_21.n9 a_96_21.t13 139.779
R65 a_96_21.n6 a_96_21.t8 139.779
R66 a_96_21.n3 a_96_21.t15 139.779
R67 a_96_21.n1 a_96_21.t12 139.779
R68 a_96_21.n14 a_96_21.n12 133.853
R69 a_96_21.n16 a_96_21.n15 109.214
R70 a_96_21.n5 a_96_21.n2 97.76
R71 a_96_21.n14 a_96_21.n13 92.5
R72 a_96_21.n8 a_96_21.n7 76
R73 a_96_21.n5 a_96_21.n4 76
R74 a_96_21.n11 a_96_21.n10 76
R75 a_96_21.n15 a_96_21.n14 56.138
R76 a_96_21.n0 a_96_21.t7 26.595
R77 a_96_21.n0 a_96_21.t6 26.595
R78 a_96_21.t0 a_96_21.n17 26.595
R79 a_96_21.n17 a_96_21.t1 26.595
R80 a_96_21.n12 a_96_21.t5 24.923
R81 a_96_21.n12 a_96_21.t3 24.923
R82 a_96_21.n13 a_96_21.t2 24.923
R83 a_96_21.n13 a_96_21.t4 24.923
R84 a_96_21.n2 a_96_21.n1 21.909
R85 a_96_21.n11 a_96_21.n8 21.76
R86 a_96_21.n8 a_96_21.n5 21.76
R87 a_96_21.n10 a_96_21.n9 13.145
R88 a_96_21.n15 a_96_21.n11 11.2
R89 a_96_21.n4 a_96_21.n3 10.224
R90 a_96_21.n7 a_96_21.n6 1.46
R91 a_484_47.n3 a_484_47.t4 219.833
R92 a_484_47.n1 a_484_47.t2 128.218
R93 a_484_47.n3 a_484_47.n2 92.5
R94 a_484_47.n1 a_484_47.n0 52.624
R95 a_484_47.n4 a_484_47.n3 51.052
R96 a_484_47.n4 a_484_47.n1 48.239
R97 a_484_47.n5 a_484_47.n4 43.173
R98 a_484_47.t5 a_484_47.n5 33.23
R99 a_484_47.n5 a_484_47.t3 31.384
R100 a_484_47.n2 a_484_47.t1 24.923
R101 a_484_47.n2 a_484_47.t0 24.923
R102 a_484_47.n0 a_484_47.t6 24.923
R103 a_484_47.n0 a_484_47.t7 24.923
R104 VNB VNB.t4 6489.08
R105 VNB.t3 VNB.t8 4545.05
R106 VNB.t9 VNB.t7 2417.58
R107 VNB.t10 VNB.t6 2030.77
R108 VNB.t11 VNB.t10 2030.77
R109 VNB.t7 VNB.t11 2030.77
R110 VNB.t1 VNB.t9 2030.77
R111 VNB.t0 VNB.t1 2030.77
R112 VNB.t8 VNB.t0 2030.77
R113 VNB.t5 VNB.t3 2030.77
R114 VNB.t2 VNB.t5 2030.77
R115 VNB.t4 VNB.t2 2030.77
R116 VGND.n14 VGND.t1 193.925
R117 VGND.n25 VGND.t2 188.321
R118 VGND.n3 VGND.n0 125.865
R119 VGND.n2 VGND.n1 115.464
R120 VGND.n20 VGND.n19 115.464
R121 VGND.n0 VGND.t4 24.923
R122 VGND.n0 VGND.t6 24.923
R123 VGND.n1 VGND.t7 24.923
R124 VGND.n1 VGND.t5 24.923
R125 VGND.n19 VGND.t3 24.923
R126 VGND.n19 VGND.t0 24.923
R127 VGND.n26 VGND.n25 13.308
R128 VGND.n3 VGND.n2 11.839
R129 VGND.n5 VGND.n4 4.65
R130 VGND.n7 VGND.n6 4.65
R131 VGND.n9 VGND.n8 4.65
R132 VGND.n11 VGND.n10 4.65
R133 VGND.n13 VGND.n12 4.65
R134 VGND.n16 VGND.n15 4.65
R135 VGND.n18 VGND.n17 4.65
R136 VGND.n22 VGND.n21 4.65
R137 VGND.n24 VGND.n23 4.65
R138 VGND.n15 VGND.n14 3.388
R139 VGND.n21 VGND.n20 2.635
R140 VGND.n5 VGND.n3 0.34
R141 VGND.n7 VGND.n5 0.119
R142 VGND.n9 VGND.n7 0.119
R143 VGND.n11 VGND.n9 0.119
R144 VGND.n13 VGND.n11 0.119
R145 VGND.n16 VGND.n13 0.119
R146 VGND.n18 VGND.n16 0.119
R147 VGND.n22 VGND.n18 0.119
R148 VGND.n24 VGND.n22 0.119
R149 VGND.n26 VGND.n24 0.119
R150 VGND VGND.n26 0.022
R151 X.n2 X.n0 155.695
R152 X.n2 X.n1 111.273
R153 X.n5 X.n3 88.89
R154 X.n5 X.n4 52.624
R155 X X.n2 39.416
R156 X X.n5 29.379
R157 X.n0 X.t7 26.595
R158 X.n0 X.t6 26.595
R159 X.n1 X.t5 26.595
R160 X.n1 X.t4 26.595
R161 X.n3 X.t1 24.923
R162 X.n3 X.t3 24.923
R163 X.n4 X.t0 24.923
R164 X.n4 X.t2 24.923
R165 B2.n0 B2.t0 212.079
R166 B2.n1 B2.t1 212.079
R167 B2.n0 B2.t3 139.779
R168 B2.n1 B2.t2 139.779
R169 B2 B2.n2 77.268
R170 B2.n2 B2.n0 30.672
R171 B2.n2 B2.n1 30.672
R172 A1.n0 A1.t0 241.534
R173 A1.n1 A1.t2 241.534
R174 A1.n2 A1.n1 184.186
R175 A1.n0 A1.t1 169.234
R176 A1.n1 A1.t3 169.234
R177 A1.n2 A1.n0 76
R178 A1 A1.n2 23.68
R179 a_918_297.n1 a_918_297.n0 496.201
R180 a_918_297.n0 a_918_297.t3 26.595
R181 a_918_297.n0 a_918_297.t1 26.595
R182 a_918_297.n1 a_918_297.t0 26.595
R183 a_918_297.t2 a_918_297.n1 26.595
R184 A2.n0 A2.t1 212.079
R185 A2.n1 A2.t0 212.079
R186 A2.n0 A2.t3 139.779
R187 A2.n1 A2.t2 139.779
R188 A2 A2.n2 81.12
R189 A2.n2 A2.n0 30.672
R190 A2.n2 A2.n1 30.672
C0 A1 A2 0.31fF
C1 X VGND 0.43fF
C2 B1 A1 0.14fF
C3 A1 VPWR 0.10fF
C4 VPB VPWR 0.13fF
C5 VPWR VGND 0.14fF
C6 VPWR X 0.52fF
C7 B1 B2 0.33fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__o22ai_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__o22ai_1 A2 B1 Y A1 B2 VGND VPWR VNB VPB
X0 VGND.t1 A2.t0 a_27_47.t1 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 a_27_47.t3 B2.t0 Y.t1 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 VPWR.t1 A1.t0 a_307_297.t1 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 a_307_297.t0 A2.t1 Y.t2 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 a_27_47.t0 A1.t1 VGND.t0 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 Y.t0 B2.t1 a_109_297.t1 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 a_109_297.t0 B1.t0 VPWR.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 Y.t3 B1.t1 a_27_47.t2 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
R0 A2.n0 A2.t1 241.534
R1 A2.n0 A2.t0 169.234
R2 A2 A2.n0 114.322
R3 a_27_47.n1 a_27_47.t2 230.648
R4 a_27_47.t0 a_27_47.n1 154.354
R5 a_27_47.n1 a_27_47.n0 46.251
R6 a_27_47.n0 a_27_47.t3 36.923
R7 a_27_47.n0 a_27_47.t1 28.615
R8 VGND VGND.n0 117.915
R9 VGND.n0 VGND.t0 24.923
R10 VGND.n0 VGND.t1 24.923
R11 VNB VNB.t2 6078.09
R12 VNB.t3 VNB.t1 2441.76
R13 VNB.t2 VNB.t3 2103.3
R14 VNB.t1 VNB.t0 2030.77
R15 B2.n0 B2.t1 239.984
R16 B2.n0 B2.t0 167.684
R17 B2 B2.n0 102.624
R18 Y.n2 Y.n0 193.794
R19 Y.n2 Y.n1 146.314
R20 Y.n1 Y.t2 65.01
R21 Y.n0 Y.t1 27.692
R22 Y.n1 Y.t0 26.595
R23 Y.n0 Y.t3 24.923
R24 Y Y.n2 2.113
R25 A1.n0 A1.t0 236.179
R26 A1.n0 A1.t1 163.879
R27 A1 A1.n0 80.16
R28 a_307_297.t0 a_307_297.t1 41.37
R29 VPWR.n0 VPWR.t0 588.653
R30 VPWR.n0 VPWR.t1 151.695
R31 VPWR VPWR.n0 0.041
R32 VPB.t1 VPB.t2 364.018
R33 VPB.t0 VPB.t1 221.962
R34 VPB.t2 VPB.t3 213.084
R35 VPB VPB.t0 192.367
R36 a_109_297.t0 a_109_297.t1 44.325
R37 B1.n0 B1.t0 230.154
R38 B1.n0 B1.t1 157.854
R39 B1 B1.n0 97.066
C0 VPWR Y 0.12fF
C1 VPWR A2 0.18fF
C2 Y B2 0.22fF
C3 B2 A2 0.12fF
C4 Y B1 0.16fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__o22ai_2.ext - technology: sky130A

.subckt sky130_fd_sc_hd__o22ai_2 B2 B1 Y A1 A2 VGND VPWR VNB VPB
X0 Y.t5 B2.t0 a_27_297.t3 VPB.t7 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 Y.t7 B2.t1 a_27_47.t7 VNB.t7 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 a_27_297.t1 B1.t0 VPWR.t1 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 a_475_297.t3 A1.t0 VPWR.t2 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 a_27_47.t0 A2.t0 VGND.t1 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 VPWR.t3 A1.t1 a_475_297.t2 VPB.t5 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 a_27_47.t4 A1.t2 VGND.t3 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 a_27_47.t2 B1.t1 Y.t2 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 Y.t3 B1.t2 a_27_47.t3 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 a_27_47.t6 B2.t2 Y.t6 VNB.t6 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 VGND.t2 A1.t3 a_27_47.t5 VNB.t5 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 VPWR.t0 B1.t3 a_27_297.t0 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 a_475_297.t0 A2.t1 Y.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13 Y.t1 A2.t2 a_475_297.t1 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14 a_27_297.t2 B2.t3 Y.t4 VPB.t6 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 VGND.t0 A2.t3 a_27_47.t1 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
R0 B2.n0 B2.t3 212.079
R1 B2.n1 B2.t0 212.079
R2 B2.n0 B2.t2 139.779
R3 B2.n1 B2.t1 139.779
R4 B2 B2.n2 34.262
R5 B2.n2 B2.n1 31.06
R6 B2.n2 B2.n0 19.887
R7 a_27_297.n1 a_27_297.t2 246.118
R8 a_27_297.t0 a_27_297.n1 202.055
R9 a_27_297.n1 a_27_297.n0 90.234
R10 a_27_297.n0 a_27_297.t3 26.595
R11 a_27_297.n0 a_27_297.t1 26.595
R12 Y.n2 Y.n0 188.606
R13 Y Y.n1 177.94
R14 Y.n5 Y.n4 145.012
R15 Y.n5 Y.n3 92.5
R16 Y Y.n5 68.77
R17 Y.n1 Y.t4 26.595
R18 Y.n1 Y.t5 26.595
R19 Y.n0 Y.t0 26.595
R20 Y.n0 Y.t1 26.595
R21 Y.n3 Y.t6 24.923
R22 Y.n3 Y.t7 24.923
R23 Y.n4 Y.t2 24.923
R24 Y.n4 Y.t3 24.923
R25 Y.n2 Y 7.466
R26 Y Y.n2 4.702
R27 VPB.t6 VPB.t1 580.062
R28 VPB.t5 VPB.t4 248.598
R29 VPB.t0 VPB.t5 248.598
R30 VPB.t1 VPB.t0 248.598
R31 VPB.t7 VPB.t6 248.598
R32 VPB.t3 VPB.t7 248.598
R33 VPB.t2 VPB.t3 248.598
R34 VPB VPB.t2 201.246
R35 a_27_47.n5 a_27_47.t3 143.301
R36 a_27_47.n2 a_27_47.t4 128.218
R37 a_27_47.n7 a_27_47.n0 102.461
R38 a_27_47.n5 a_27_47.n4 92.5
R39 a_27_47.n7 a_27_47.n6 92.5
R40 a_27_47.n3 a_27_47.n2 67.512
R41 a_27_47.n6 a_27_47.n5 63.247
R42 a_27_47.n2 a_27_47.n1 52.624
R43 a_27_47.n6 a_27_47.n3 41.788
R44 a_27_47.n0 a_27_47.t1 25.846
R45 a_27_47.n4 a_27_47.t7 24.923
R46 a_27_47.n4 a_27_47.t2 24.923
R47 a_27_47.n1 a_27_47.t5 24.923
R48 a_27_47.n1 a_27_47.t0 24.923
R49 a_27_47.t6 a_27_47.n7 24.923
R50 VNB VNB.t3 6150.61
R51 VNB.t6 VNB.t1 4738.46
R52 VNB.t5 VNB.t4 2030.77
R53 VNB.t0 VNB.t5 2030.77
R54 VNB.t1 VNB.t0 2030.77
R55 VNB.t7 VNB.t6 2030.77
R56 VNB.t2 VNB.t7 2030.77
R57 VNB.t3 VNB.t2 2030.77
R58 B1.n0 B1.t0 212.079
R59 B1.n1 B1.t3 212.079
R60 B1.n0 B1.t1 139.779
R61 B1.n1 B1.t2 139.779
R62 B1 B1.n2 34.095
R63 B1.n2 B1.n0 32.392
R64 B1.n2 B1.n1 18.507
R65 VPWR.n2 VPWR.n0 176.458
R66 VPWR.n2 VPWR.n1 175.493
R67 VPWR.n0 VPWR.t2 26.595
R68 VPWR.n0 VPWR.t3 26.595
R69 VPWR.n1 VPWR.t1 26.595
R70 VPWR.n1 VPWR.t0 26.595
R71 VPWR VPWR.n2 0.142
R72 A1.n0 A1.t0 212.079
R73 A1.n1 A1.t1 212.079
R74 A1.n0 A1.t2 139.779
R75 A1.n1 A1.t3 139.779
R76 A1 A1.n2 34.107
R77 A1.n2 A1.n1 32.128
R78 A1.n2 A1.n0 18.771
R79 a_475_297.n0 a_475_297.t1 246.12
R80 a_475_297.n0 a_475_297.t3 202.055
R81 a_475_297.n1 a_475_297.n0 90.234
R82 a_475_297.t2 a_475_297.n1 26.595
R83 a_475_297.n1 a_475_297.t0 26.595
R84 A2.n0 A2.t1 212.079
R85 A2.n1 A2.t2 212.079
R86 A2.n0 A2.t0 139.779
R87 A2.n1 A2.t3 139.779
R88 A2 A2.n2 34.307
R89 A2.n2 A2.n0 31.337
R90 A2.n2 A2.n1 19.611
R91 VGND.n2 VGND.n0 124.932
R92 VGND.n2 VGND.n1 121.761
R93 VGND.n0 VGND.t3 24.923
R94 VGND.n0 VGND.t2 24.923
R95 VGND.n1 VGND.t1 24.923
R96 VGND.n1 VGND.t0 24.923
R97 VGND VGND.n2 0.854
C0 B2 Y 0.26fF
C1 A2 Y 0.12fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__o22ai_4.ext - technology: sky130A

.subckt sky130_fd_sc_hd__o22ai_4 A1 Y A2 B1 B2 VGND VPWR VNB VPB
X0 a_33_47.t3 B2.t0 Y.t5 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 VGND.t3 A1.t0 a_33_47.t5 VNB.t5 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 VGND.t5 A2.t0 a_33_47.t13 VNB.t13 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 a_33_47.t9 B1.t0 Y.t10 VNB.t9 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 a_797_297.t7 B2.t1 Y.t7 VPB.t11 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 Y.t14 A2.t1 a_115_297.t7 VPB.t15 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 a_797_297.t3 B1.t1 VPWR.t7 VPB.t7 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 Y.t6 B2.t2 a_797_297.t6 VPB.t10 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 a_115_297.t6 A2.t2 Y.t15 VPB.t14 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 VPWR.t6 B1.t2 a_797_297.t2 VPB.t6 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 a_33_47.t6 A1.t1 VGND.t2 VNB.t6 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 VGND.t1 A1.t2 a_33_47.t7 VNB.t7 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 a_33_47.t14 A2.t3 VGND.t6 VNB.t14 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 a_33_47.t15 A2.t4 VGND.t7 VNB.t15 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14 Y.t8 A2.t5 a_115_297.t5 VPB.t13 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 a_33_47.t8 A1.t3 VGND.t0 VNB.t8 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X16 a_797_297.t1 B1.t3 VPWR.t5 VPB.t5 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17 a_115_297.t3 A1.t4 VPWR.t3 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X18 VPWR.t2 A1.t5 a_115_297.t2 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X19 VPWR.t4 B1.t4 a_797_297.t0 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X20 VGND.t4 A2.t6 a_33_47.t4 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X21 a_33_47.t10 B1.t5 Y.t11 VNB.t10 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X22 a_797_297.t5 B2.t3 Y.t1 VPB.t9 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X23 VPWR.t1 A1.t6 a_115_297.t1 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X24 Y.t4 B2.t4 a_33_47.t2 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X25 Y.t0 B2.t5 a_797_297.t4 VPB.t8 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X26 Y.t12 B1.t6 a_33_47.t11 VNB.t11 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X27 Y.t3 B2.t6 a_33_47.t1 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X28 a_115_297.t4 A2.t7 Y.t9 VPB.t12 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X29 Y.t13 B1.t7 a_33_47.t12 VNB.t12 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X30 a_33_47.t0 B2.t7 Y.t2 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X31 a_115_297.t0 A1.t7 VPWR.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
R0 B2.n0 B2.t3 212.079
R1 B2.n7 B2.t5 212.079
R2 B2.n4 B2.t1 212.079
R3 B2.n2 B2.t2 212.079
R4 B2.n0 B2.t6 139.779
R5 B2.n7 B2.t0 139.779
R6 B2.n4 B2.t4 139.779
R7 B2.n2 B2.t7 139.779
R8 B2.n6 B2.n3 97.76
R9 B2 B2.n1 86.88
R10 B2.n9 B2.n8 76
R11 B2.n6 B2.n5 76
R12 B2.n9 B2.n6 21.76
R13 B2.n1 B2.n0 19.718
R14 B2.n3 B2.n2 15.336
R15 B2 B2.n9 10.88
R16 B2.n8 B2.n7 8.033
R17 B2.n5 B2.n4 3.651
R18 Y.n13 Y.n12 346.333
R19 Y.n2 Y.n1 346.333
R20 Y.n2 Y.n0 292.5
R21 Y.n13 Y.n11 292.5
R22 Y.n4 Y.n2 181.214
R23 Y.n14 Y.n10 148.908
R24 Y.n10 Y.n9 92.5
R25 Y.n8 Y.n7 92.5
R26 Y.n6 Y.n5 92.5
R27 Y.n4 Y.n3 92.5
R28 Y.n6 Y.n4 61.44
R29 Y.n8 Y.n6 61.44
R30 Y.n10 Y.n8 61.44
R31 Y.n11 Y.t9 26.595
R32 Y.n11 Y.t14 26.595
R33 Y.n12 Y.t15 26.595
R34 Y.n12 Y.t8 26.595
R35 Y.n0 Y.t1 26.595
R36 Y.n0 Y.t0 26.595
R37 Y.n1 Y.t7 26.595
R38 Y.n1 Y.t6 26.595
R39 Y.n3 Y.t10 24.923
R40 Y.n3 Y.t3 24.923
R41 Y.n5 Y.t5 24.923
R42 Y.n5 Y.t4 24.923
R43 Y.n7 Y.t2 24.923
R44 Y.n7 Y.t13 24.923
R45 Y.n9 Y.t11 24.923
R46 Y.n9 Y.t12 24.923
R47 Y Y.n13 3.576
R48 Y Y.n14 2.258
R49 Y.n14 Y 1.129
R50 a_33_47.n12 a_33_47.t9 219.833
R51 a_33_47.n3 a_33_47.t7 128.218
R52 a_33_47.n11 a_33_47.n0 92.5
R53 a_33_47.n10 a_33_47.n1 92.5
R54 a_33_47.n13 a_33_47.n12 92.5
R55 a_33_47.n3 a_33_47.n2 52.624
R56 a_33_47.n5 a_33_47.n4 52.624
R57 a_33_47.n7 a_33_47.n6 52.624
R58 a_33_47.n10 a_33_47.n9 51.719
R59 a_33_47.n9 a_33_47.n7 49.159
R60 a_33_47.n12 a_33_47.n11 48.872
R61 a_33_47.n11 a_33_47.n10 48.872
R62 a_33_47.n9 a_33_47.n8 42.888
R63 a_33_47.n5 a_33_47.n3 38.786
R64 a_33_47.n7 a_33_47.n5 36.266
R65 a_33_47.n8 a_33_47.t11 34.153
R66 a_33_47.n1 a_33_47.t12 24.923
R67 a_33_47.n1 a_33_47.t10 24.923
R68 a_33_47.n0 a_33_47.t2 24.923
R69 a_33_47.n0 a_33_47.t0 24.923
R70 a_33_47.n8 a_33_47.t8 24.923
R71 a_33_47.n6 a_33_47.t4 24.923
R72 a_33_47.n6 a_33_47.t15 24.923
R73 a_33_47.n4 a_33_47.t13 24.923
R74 a_33_47.n4 a_33_47.t14 24.923
R75 a_33_47.n2 a_33_47.t5 24.923
R76 a_33_47.n2 a_33_47.t6 24.923
R77 a_33_47.n13 a_33_47.t1 24.923
R78 a_33_47.t3 a_33_47.n13 24.923
R79 VNB VNB.t7 6223.14
R80 VNB.t8 VNB.t11 2272.53
R81 VNB.t1 VNB.t9 2030.77
R82 VNB.t3 VNB.t1 2030.77
R83 VNB.t2 VNB.t3 2030.77
R84 VNB.t0 VNB.t2 2030.77
R85 VNB.t12 VNB.t0 2030.77
R86 VNB.t10 VNB.t12 2030.77
R87 VNB.t11 VNB.t10 2030.77
R88 VNB.t4 VNB.t8 2030.77
R89 VNB.t15 VNB.t4 2030.77
R90 VNB.t13 VNB.t15 2030.77
R91 VNB.t14 VNB.t13 2030.77
R92 VNB.t5 VNB.t14 2030.77
R93 VNB.t6 VNB.t5 2030.77
R94 VNB.t7 VNB.t6 2030.77
R95 A1.n1 A1.n0 248.98
R96 A1.n0 A1.t6 241.534
R97 A1.n2 A1.t4 212.079
R98 A1.n5 A1.t5 212.079
R99 A1.n3 A1.t7 212.079
R100 A1.n0 A1.t3 169.234
R101 A1.n2 A1.t0 139.779
R102 A1.n5 A1.t1 139.779
R103 A1.n3 A1.t2 139.779
R104 A1.n7 A1.n6 76
R105 A1.n6 A1.n5 48.2
R106 A1.n4 A1 43.175
R107 A1.n4 A1.n3 31.954
R108 A1.n5 A1.n4 18.353
R109 A1.n6 A1.n2 13.145
R110 A1 A1.n1 5.44
R111 A1 A1.n7 2.656
R112 A1.n7 A1.n1 0.724
R113 VGND.n3 VGND.n0 126.078
R114 VGND.n2 VGND.n1 115.464
R115 VGND.n7 VGND.n6 115.464
R116 VGND.n13 VGND.n12 115.464
R117 VGND.n0 VGND.t0 24.923
R118 VGND.n0 VGND.t4 24.923
R119 VGND.n1 VGND.t7 24.923
R120 VGND.n1 VGND.t5 24.923
R121 VGND.n6 VGND.t6 24.923
R122 VGND.n6 VGND.t3 24.923
R123 VGND.n12 VGND.t2 24.923
R124 VGND.n12 VGND.t1 24.923
R125 VGND.n3 VGND.n2 14.445
R126 VGND.n14 VGND.n13 5.652
R127 VGND.n5 VGND.n4 4.65
R128 VGND.n9 VGND.n8 4.65
R129 VGND.n11 VGND.n10 4.65
R130 VGND.n8 VGND.n7 4.517
R131 VGND.n5 VGND.n3 0.37
R132 VGND.n14 VGND.n11 0.132
R133 VGND VGND.n14 0.129
R134 VGND.n9 VGND.n5 0.119
R135 VGND.n11 VGND.n9 0.119
R136 A2.n0 A2.t7 212.079
R137 A2.n2 A2.t1 212.079
R138 A2.n7 A2.t2 212.079
R139 A2.n5 A2.t5 212.079
R140 A2.n0 A2.t6 139.779
R141 A2.n2 A2.t4 139.779
R142 A2.n7 A2.t0 139.779
R143 A2.n5 A2.t3 139.779
R144 A2.n9 A2.n6 97.76
R145 A2.n4 A2.n1 97.76
R146 A2.n4 A2.n3 76
R147 A2.n9 A2.n8 76
R148 A2.n6 A2.n5 21.909
R149 A2.n1 A2.n0 13.145
R150 A2 A2.n9 12.48
R151 A2.n8 A2.n7 10.224
R152 A2 A2.n4 9.28
R153 A2.n3 A2.n2 1.46
R154 B1.n0 B1.t4 238.589
R155 B1 B1.n0 235.199
R156 B1.n1 B1.t1 212.079
R157 B1.n3 B1.t2 212.079
R158 B1.n2 B1.t3 212.079
R159 B1.n0 B1.t0 166.289
R160 B1.n1 B1.t7 139.779
R161 B1.n3 B1.t5 139.779
R162 B1.n2 B1.t6 139.779
R163 B1.n3 B1.n2 61.345
R164 B1 B1.n4 30.752
R165 B1.n4 B1.n3 27.06
R166 B1.n4 B1.n1 22.468
R167 a_797_297.n4 a_797_297.n3 375.897
R168 a_797_297.n2 a_797_297.n0 346.476
R169 a_797_297.n2 a_797_297.n1 292.5
R170 a_797_297.n5 a_797_297.n4 142.024
R171 a_797_297.n4 a_797_297.n2 61.678
R172 a_797_297.n3 a_797_297.t2 26.595
R173 a_797_297.n3 a_797_297.t1 26.595
R174 a_797_297.n1 a_797_297.t4 26.595
R175 a_797_297.n1 a_797_297.t7 26.595
R176 a_797_297.n0 a_797_297.t0 26.595
R177 a_797_297.n0 a_797_297.t5 26.595
R178 a_797_297.t6 a_797_297.n5 26.595
R179 a_797_297.n5 a_797_297.t3 26.595
R180 VPB.t1 VPB.t5 278.193
R181 VPB.t9 VPB.t4 248.598
R182 VPB.t8 VPB.t9 248.598
R183 VPB.t11 VPB.t8 248.598
R184 VPB.t10 VPB.t11 248.598
R185 VPB.t7 VPB.t10 248.598
R186 VPB.t6 VPB.t7 248.598
R187 VPB.t5 VPB.t6 248.598
R188 VPB.t12 VPB.t1 248.598
R189 VPB.t15 VPB.t12 248.598
R190 VPB.t14 VPB.t15 248.598
R191 VPB.t13 VPB.t14 248.598
R192 VPB.t3 VPB.t13 248.598
R193 VPB.t2 VPB.t3 248.598
R194 VPB.t0 VPB.t2 248.598
R195 VPB VPB.t0 210.124
R196 a_115_297.n4 a_115_297.n0 346.333
R197 a_115_297.n5 a_115_297.n4 292.5
R198 a_115_297.n3 a_115_297.n1 160.328
R199 a_115_297.n3 a_115_297.n2 142.024
R200 a_115_297.n4 a_115_297.n3 61.677
R201 a_115_297.n2 a_115_297.t5 26.595
R202 a_115_297.n2 a_115_297.t3 26.595
R203 a_115_297.n1 a_115_297.t2 26.595
R204 a_115_297.n1 a_115_297.t0 26.595
R205 a_115_297.n0 a_115_297.t1 26.595
R206 a_115_297.n0 a_115_297.t4 26.595
R207 a_115_297.n5 a_115_297.t7 26.595
R208 a_115_297.t6 a_115_297.n5 26.595
R209 VPWR.n0 VPWR.t4 554.815
R210 VPWR.n8 VPWR.n7 316.936
R211 VPWR.n2 VPWR.n1 314.9
R212 VPWR.n20 VPWR.n19 314.004
R213 VPWR.n24 VPWR.t0 154.764
R214 VPWR.n7 VPWR.t1 34.475
R215 VPWR.n7 VPWR.t5 28.565
R216 VPWR.n19 VPWR.t3 26.595
R217 VPWR.n19 VPWR.t2 26.595
R218 VPWR.n1 VPWR.t7 26.595
R219 VPWR.n1 VPWR.t6 26.595
R220 VPWR.n9 VPWR.n8 8.658
R221 VPWR.n4 VPWR.n3 4.65
R222 VPWR.n6 VPWR.n5 4.65
R223 VPWR.n10 VPWR.n9 4.65
R224 VPWR.n12 VPWR.n11 4.65
R225 VPWR.n14 VPWR.n13 4.65
R226 VPWR.n16 VPWR.n15 4.65
R227 VPWR.n18 VPWR.n17 4.65
R228 VPWR.n21 VPWR.n20 4.65
R229 VPWR.n23 VPWR.n22 4.65
R230 VPWR.n25 VPWR.n24 4.65
R231 VPWR.n3 VPWR.n2 4.141
R232 VPWR.n4 VPWR.n0 0.134
R233 VPWR.n6 VPWR.n4 0.119
R234 VPWR.n10 VPWR.n6 0.119
R235 VPWR.n12 VPWR.n10 0.119
R236 VPWR.n14 VPWR.n12 0.119
R237 VPWR.n16 VPWR.n14 0.119
R238 VPWR.n18 VPWR.n16 0.119
R239 VPWR.n21 VPWR.n18 0.119
R240 VPWR.n23 VPWR.n21 0.119
R241 VPWR.n25 VPWR.n23 0.119
R242 VPWR VPWR.n25 0.022
C0 VPWR Y 0.18fF
C1 VPB VPWR 0.14fF
C2 VPWR VGND 0.15fF
C3 B1 Y 0.70fF
C4 A1 A2 0.53fF
C5 B2 Y 0.18fF
C6 B1 B2 0.52fF
C7 A1 Y 0.35fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__o31a_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__o31a_1 X A2 B1 A1 A3 VGND VPWR VNB VPB
X0 a_103_199.t2 B1.t0 a_253_47.t3 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 VPWR.t1 a_103_199.t3 X.t0 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 a_337_297.t1 A2.t0 a_253_297.t0 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 a_103_199.t0 A3.t0 a_337_297.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 a_253_297.t1 A1.t0 VPWR.t2 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 VPWR.t0 B1.t1 a_103_199.t1 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 VGND.t3 a_103_199.t4 X.t1 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 a_253_47.t0 A1.t1 VGND.t1 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 a_253_47.t2 A3.t1 VGND.t0 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 VGND.t2 A2.t1 a_253_47.t1 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
R0 B1.n0 B1.t1 238.154
R1 B1.n0 B1.t0 165.854
R2 B1 B1.n0 80.848
R3 a_253_47.n1 a_253_47.n0 265.792
R4 a_253_47.n0 a_253_47.t3 30.461
R5 a_253_47.n0 a_253_47.t2 30.461
R6 a_253_47.n1 a_253_47.t1 24.923
R7 a_253_47.t0 a_253_47.n1 24.923
R8 a_103_199.n1 a_103_199.n0 297.399
R9 a_103_199.n0 a_103_199.t3 241.534
R10 a_103_199.n1 a_103_199.t2 184.907
R11 a_103_199.n0 a_103_199.t4 169.234
R12 a_103_199.n2 a_103_199.n1 138.493
R13 a_103_199.t0 a_103_199.n2 56.145
R14 a_103_199.n2 a_103_199.t1 27.58
R15 VNB VNB.t4 6948.42
R16 VNB.t4 VNB.t0 2610.99
R17 VNB.t2 VNB.t3 2320.88
R18 VNB.t1 VNB.t2 2320.88
R19 VNB.t0 VNB.t1 2030.77
R20 X.n0 X.t0 188.677
R21 X X.n2 94.39
R22 X.n3 X.n2 92.5
R23 X.n2 X.t1 39.692
R24 X X.n4 11.561
R25 X.n3 X 8
R26 X.n1 X.n0 5.997
R27 X.n4 X 2.477
R28 X.n0 X 2.402
R29 X X.n1 2.064
R30 X X.n3 1.89
R31 X.n4 X 1.745
R32 X.n1 X 1.454
R33 VPWR.n1 VPWR.t0 213.54
R34 VPWR.n1 VPWR.n0 170.313
R35 VPWR.n0 VPWR.t2 38.415
R36 VPWR.n0 VPWR.t1 38.415
R37 VPWR VPWR.n1 0.167
R38 VPB.t0 VPB.t2 340.342
R39 VPB.t3 VPB.t4 319.626
R40 VPB VPB.t3 298.909
R41 VPB.t1 VPB.t0 284.112
R42 VPB.t4 VPB.t1 248.598
R43 A2.n0 A2.t0 241.534
R44 A2.n0 A2.t1 169.234
R45 A2.n1 A2.n0 76
R46 A2 A2.n1 16.3
R47 A2.n1 A2 2.873
R48 a_253_297.t0 a_253_297.t1 53.19
R49 a_337_297.t0 a_337_297.t1 65.01
R50 A3.n0 A3.t0 241.534
R51 A3.n0 A3.t1 169.234
R52 A3 A3.n0 77.189
R53 A1.n0 A1.t0 241.534
R54 A1.n0 A1.t1 169.234
R55 A1 A1.n0 78.971
R56 VGND.n2 VGND.n1 97.749
R57 VGND.n2 VGND.n0 60.907
R58 VGND.n0 VGND.t1 36
R59 VGND.n0 VGND.t3 36
R60 VGND.n1 VGND.t0 30.461
R61 VGND.n1 VGND.t2 30.461
R62 VGND VGND.n2 0.306
C0 A2 A3 0.16fF
C1 X VGND 0.17fF
C2 A1 A2 0.10fF
C3 X VPWR 0.19fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__o31a_2.ext - technology: sky130A

.subckt sky130_fd_sc_hd__o31a_2 X A1 A2 B1 A3 VGND VPWR VNB VPB
X0 a_108_21.t1 B1.t0 a_346_47.t1 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 a_346_47.t3 A3.t0 VGND.t4 VNB.t5 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 X.t3 a_108_21.t3 VGND.t3 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 a_108_21.t2 A3.t1 a_430_297.t1 VPB.t5 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 a_430_297.t0 A2.t0 a_346_297.t1 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 VPWR.t3 a_108_21.t4 X.t1 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 a_346_297.t0 A1.t0 VPWR.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 VGND.t1 A2.t1 a_346_47.t2 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 X.t0 a_108_21.t5 VPWR.t2 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 VPWR.t1 B1.t1 a_108_21.t0 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 VGND.t2 a_108_21.t6 X.t2 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 a_346_47.t0 A1.t1 VGND.t0 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
R0 B1.n0 B1.t1 238.154
R1 B1.n0 B1.t0 165.854
R2 B1 B1.n0 80.848
R3 a_346_47.n1 a_346_47.n0 265.792
R4 a_346_47.n0 a_346_47.t1 30.461
R5 a_346_47.n0 a_346_47.t3 30.461
R6 a_346_47.n1 a_346_47.t2 24.923
R7 a_346_47.t0 a_346_47.n1 24.923
R8 a_108_21.n2 a_108_21.n1 297.399
R9 a_108_21.n1 a_108_21.t4 212.079
R10 a_108_21.n0 a_108_21.t5 212.079
R11 a_108_21.n2 a_108_21.t1 184.585
R12 a_108_21.n1 a_108_21.t6 139.779
R13 a_108_21.n0 a_108_21.t3 139.779
R14 a_108_21.n3 a_108_21.n2 138.493
R15 a_108_21.n1 a_108_21.n0 73.03
R16 a_108_21.n3 a_108_21.t2 56.145
R17 a_108_21.t0 a_108_21.n3 27.58
R18 VNB VNB.t4 6755.01
R19 VNB.t3 VNB.t0 2610.99
R20 VNB.t4 VNB.t3 2417.58
R21 VNB.t5 VNB.t1 2320.88
R22 VNB.t2 VNB.t5 2320.88
R23 VNB.t0 VNB.t2 2030.77
R24 A3.n0 A3.t1 241.534
R25 A3.n0 A3.t0 169.234
R26 A3 A3.n0 77.189
R27 VGND.n8 VGND.t3 118.032
R28 VGND.n3 VGND.n2 97.618
R29 VGND.n1 VGND.n0 58.789
R30 VGND.n0 VGND.t0 36
R31 VGND.n0 VGND.t2 36
R32 VGND.n2 VGND.t4 30.461
R33 VGND.n2 VGND.t1 30.461
R34 VGND.n9 VGND.n8 4.65
R35 VGND.n5 VGND.n4 4.65
R36 VGND.n7 VGND.n6 4.65
R37 VGND.n3 VGND.n1 3.927
R38 VGND.n5 VGND.n3 0.341
R39 VGND.n7 VGND.n5 0.119
R40 VGND.n9 VGND.n7 0.119
R41 VGND VGND.n9 0.02
R42 X.n1 X.n0 146.322
R43 X X.n3 94.39
R44 X.n4 X.n3 92.5
R45 X.n0 X.t1 42.355
R46 X.n3 X.t2 39.692
R47 X.n0 X.t0 26.595
R48 X.n3 X.t3 24.923
R49 X.n6 X 23.272
R50 X X.n5 11.561
R51 X X.n6 10.735
R52 X.n4 X 8
R53 X.n2 X.n1 5.997
R54 X.n6 X 3.303
R55 X.n5 X 2.477
R56 X.n1 X 2.402
R57 X X.n2 2.064
R58 X X.n4 1.89
R59 X.n5 X 1.745
R60 X.n2 X 1.454
R61 a_430_297.t0 a_430_297.t1 65.01
R62 VPB.t5 VPB.t1 340.342
R63 VPB.t4 VPB.t0 319.626
R64 VPB.t3 VPB.t4 295.95
R65 VPB.t2 VPB.t5 284.112
R66 VPB VPB.t3 275.233
R67 VPB.t0 VPB.t2 248.598
R68 A2.n0 A2.t0 241.534
R69 A2.n0 A2.t1 169.234
R70 A2.n1 A2.n0 76
R71 A2 A2.n1 16.3
R72 A2.n1 A2 2.873
R73 a_346_297.t0 a_346_297.t1 53.19
R74 VPWR.n0 VPWR.t1 212.152
R75 VPWR.n7 VPWR.t2 177.307
R76 VPWR.n2 VPWR.n1 166.691
R77 VPWR.n1 VPWR.t0 38.415
R78 VPWR.n1 VPWR.t3 38.415
R79 VPWR.n4 VPWR.n3 4.65
R80 VPWR.n6 VPWR.n5 4.65
R81 VPWR.n8 VPWR.n7 4.65
R82 VPWR.n3 VPWR.n2 1.129
R83 VPWR.n4 VPWR.n0 0.135
R84 VPWR.n6 VPWR.n4 0.119
R85 VPWR.n8 VPWR.n6 0.119
R86 VPWR VPWR.n8 0.02
R87 A1.n0 A1.t0 241.534
R88 A1.n0 A1.t1 169.234
R89 A1 A1.n0 78.971
C0 VPWR X 0.34fF
C1 A2 A3 0.16fF
C2 A1 A2 0.10fF
C3 X VGND 0.29fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__o31a_4.ext - technology: sky130A

.subckt sky130_fd_sc_hd__o31a_4 X B1 A3 A2 A1 VGND VPWR VNB VPB
X0 VPWR.t3 A1.t0 a_926_297.t3 VPB.t5 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 VGND.t4 A1.t1 a_496_47.t6 VNB.t6 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 a_926_297.t2 A1.t2 VPWR.t2 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 VGND.t0 A3.t0 a_496_47.t0 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 VGND.t6 a_102_21.t6 X.t7 VNB.t8 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 VGND.t1 A2.t0 a_496_47.t3 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 a_926_297.t0 A2.t1 a_672_297.t3 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 a_102_21.t0 B1.t0 VPWR.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 a_496_47.t4 A2.t2 VGND.t2 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 X.t6 a_102_21.t7 VGND.t7 VNB.t9 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 a_102_21.t1 B1.t1 a_496_47.t1 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 VPWR.t4 a_102_21.t8 X.t3 VPB.t8 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 X.t5 a_102_21.t9 VGND.t8 VNB.t10 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 X.t2 a_102_21.t10 VPWR.t5 VPB.t9 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14 VPWR.t6 a_102_21.t11 X.t1 VPB.t10 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 a_672_297.t1 A3.t1 a_102_21.t5 VPB.t7 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16 a_496_47.t2 B1.t2 a_102_21.t2 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X17 a_102_21.t4 A3.t2 a_672_297.t0 VPB.t6 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X18 VGND.t9 a_102_21.t12 X.t4 VNB.t11 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X19 X.t0 a_102_21.t13 VPWR.t7 VPB.t11 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X20 a_496_47.t7 A3.t3 VGND.t5 VNB.t7 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X21 VPWR.t1 B1.t3 a_102_21.t3 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X22 a_496_47.t5 A1.t3 VGND.t3 VNB.t5 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X23 a_672_297.t2 A2.t3 a_926_297.t1 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
R0 A1.n0 A1.t2 221.719
R1 A1.n1 A1.t0 221.719
R2 A1.n0 A1.t1 149.419
R3 A1.n1 A1.t3 149.419
R4 A1 A1.n2 80.196
R5 A1.n2 A1.n1 58.911
R6 A1.n2 A1.n0 16.066
R7 a_926_297.n1 a_926_297.n0 638.76
R8 a_926_297.n0 a_926_297.t1 26.595
R9 a_926_297.n0 a_926_297.t2 26.595
R10 a_926_297.n1 a_926_297.t3 26.595
R11 a_926_297.t0 a_926_297.n1 26.595
R12 VPWR.n1 VPWR.t1 570.302
R13 VPWR.n2 VPWR.n0 310.351
R14 VPWR.n15 VPWR.t7 186.806
R15 VPWR.n11 VPWR.n10 163.438
R16 VPWR.n6 VPWR.n5 118.495
R17 VPWR.n10 VPWR.t5 29.55
R18 VPWR.n10 VPWR.t6 29.55
R19 VPWR.n5 VPWR.t0 26.595
R20 VPWR.n5 VPWR.t4 26.595
R21 VPWR.n0 VPWR.t2 26.595
R22 VPWR.n0 VPWR.t3 26.595
R23 VPWR.n4 VPWR.n3 4.65
R24 VPWR.n7 VPWR.n6 4.65
R25 VPWR.n9 VPWR.n8 4.65
R26 VPWR.n12 VPWR.n11 4.65
R27 VPWR.n14 VPWR.n13 4.65
R28 VPWR.n16 VPWR.n15 4.65
R29 VPWR.n2 VPWR.n1 4.006
R30 VPWR.n4 VPWR.n2 0.138
R31 VPWR.n7 VPWR.n4 0.119
R32 VPWR.n9 VPWR.n7 0.119
R33 VPWR.n12 VPWR.n9 0.119
R34 VPWR.n14 VPWR.n12 0.119
R35 VPWR.n16 VPWR.n14 0.119
R36 VPWR VPWR.n16 0.027
R37 VPB.t1 VPB.t6 580.062
R38 VPB VPB.t11 272.274
R39 VPB.t10 VPB.t9 266.355
R40 VPB.t0 VPB.t1 260.436
R41 VPB.t4 VPB.t3 248.598
R42 VPB.t5 VPB.t4 248.598
R43 VPB.t2 VPB.t5 248.598
R44 VPB.t7 VPB.t2 248.598
R45 VPB.t6 VPB.t7 248.598
R46 VPB.t8 VPB.t0 248.598
R47 VPB.t9 VPB.t8 248.598
R48 VPB.t11 VPB.t10 248.598
R49 a_496_47.n4 a_496_47.t1 236.423
R50 a_496_47.n2 a_496_47.t4 162.247
R51 a_496_47.n3 a_496_47.n0 98.147
R52 a_496_47.n2 a_496_47.n1 98.147
R53 a_496_47.n5 a_496_47.n4 92.5
R54 a_496_47.n4 a_496_47.n3 49.596
R55 a_496_47.n3 a_496_47.n2 43.008
R56 a_496_47.t0 a_496_47.n5 30.461
R57 a_496_47.n5 a_496_47.t2 26.769
R58 a_496_47.n0 a_496_47.t3 24.923
R59 a_496_47.n0 a_496_47.t7 24.923
R60 a_496_47.n1 a_496_47.t6 24.923
R61 a_496_47.n1 a_496_47.t5 24.923
R62 VGND.n24 VGND.t8 175.576
R63 VGND.n3 VGND.n0 109.768
R64 VGND.n2 VGND.n1 106.463
R65 VGND.n7 VGND.n6 106.463
R66 VGND.n20 VGND.n19 106.463
R67 VGND.n15 VGND.t6 104.361
R68 VGND.n19 VGND.t7 27.692
R69 VGND.n19 VGND.t9 27.692
R70 VGND.n0 VGND.t2 24.923
R71 VGND.n0 VGND.t4 24.923
R72 VGND.n1 VGND.t3 24.923
R73 VGND.n1 VGND.t1 24.923
R74 VGND.n6 VGND.t5 24.923
R75 VGND.n6 VGND.t0 24.923
R76 VGND.n25 VGND.n24 7.596
R77 VGND.n5 VGND.n4 4.65
R78 VGND.n8 VGND.n7 4.65
R79 VGND.n10 VGND.n9 4.65
R80 VGND.n12 VGND.n11 4.65
R81 VGND.n14 VGND.n13 4.65
R82 VGND.n16 VGND.n15 4.65
R83 VGND.n18 VGND.n17 4.65
R84 VGND.n21 VGND.n20 4.65
R85 VGND.n23 VGND.n22 4.65
R86 VGND.n3 VGND.n2 3.896
R87 VGND.n5 VGND.n3 0.264
R88 VGND.n8 VGND.n5 0.119
R89 VGND.n10 VGND.n8 0.119
R90 VGND.n12 VGND.n10 0.119
R91 VGND.n14 VGND.n12 0.119
R92 VGND.n16 VGND.n14 0.119
R93 VGND.n18 VGND.n16 0.119
R94 VGND.n21 VGND.n18 0.119
R95 VGND.n23 VGND.n21 0.119
R96 VGND.n25 VGND.n23 0.119
R97 VGND VGND.n25 0.027
R98 VNB VNB.t10 6730.83
R99 VNB.t8 VNB.t1 4641.76
R100 VNB.t2 VNB.t0 2224.18
R101 VNB.t11 VNB.t9 2175.82
R102 VNB.t6 VNB.t4 2030.77
R103 VNB.t5 VNB.t6 2030.77
R104 VNB.t3 VNB.t5 2030.77
R105 VNB.t7 VNB.t3 2030.77
R106 VNB.t0 VNB.t7 2030.77
R107 VNB.t1 VNB.t2 2030.77
R108 VNB.t9 VNB.t8 2030.77
R109 VNB.t10 VNB.t11 2030.77
R110 A3.n0 A3.t1 221.719
R111 A3.n1 A3.t2 221.719
R112 A3.n0 A3.t3 149.419
R113 A3.n1 A3.t0 149.419
R114 A3 A3.n2 80.406
R115 A3.n2 A3.n1 38.381
R116 A3.n2 A3.n0 36.596
R117 a_102_21.n10 a_102_21.n9 232.533
R118 a_102_21.n5 a_102_21.t8 221.719
R119 a_102_21.n3 a_102_21.t10 221.719
R120 a_102_21.n2 a_102_21.t11 221.719
R121 a_102_21.n1 a_102_21.t13 221.719
R122 a_102_21.n5 a_102_21.t6 149.419
R123 a_102_21.n3 a_102_21.t7 149.419
R124 a_102_21.n2 a_102_21.t12 149.419
R125 a_102_21.n1 a_102_21.t9 149.419
R126 a_102_21.n11 a_102_21.n10 146.805
R127 a_102_21.n8 a_102_21.n0 131.924
R128 a_102_21.n7 a_102_21.n6 76
R129 a_102_21.n2 a_102_21.n1 74.977
R130 a_102_21.n7 a_102_21.n4 49.588
R131 a_102_21.n4 a_102_21.n2 42.664
R132 a_102_21.n10 a_102_21.n8 41.563
R133 a_102_21.n8 a_102_21.n7 40.306
R134 a_102_21.t0 a_102_21.n11 30.535
R135 a_102_21.n9 a_102_21.t5 26.595
R136 a_102_21.n9 a_102_21.t4 26.595
R137 a_102_21.n11 a_102_21.t3 26.595
R138 a_102_21.n0 a_102_21.t2 24.923
R139 a_102_21.n0 a_102_21.t1 24.923
R140 a_102_21.n4 a_102_21.n3 21.736
R141 a_102_21.n6 a_102_21.n5 16.066
R142 X.n8 X.n5 209.736
R143 X.n8 X.n6 166.323
R144 X.n3 X.n2 139.804
R145 X.n1 X.n0 92.5
R146 X X.n3 88.145
R147 X.n9 X.n4 73.309
R148 X.n5 X.t3 26.595
R149 X.n5 X.t2 26.595
R150 X.n6 X.t1 26.595
R151 X.n6 X.t0 26.595
R152 X.n2 X.t7 24.923
R153 X.n2 X.t6 24.923
R154 X.n0 X.t4 24.923
R155 X.n0 X.t5 24.923
R156 X X.n9 6.884
R157 X.n8 X.n7 5.953
R158 X.n9 X 4.654
R159 X.n7 X 3.49
R160 X.n4 X.n1 3.339
R161 X X.n8 2.473
R162 X.n4 X 1.163
R163 X.n3 X.n1 1.113
R164 X.n7 X 0.893
R165 X.n9 X 0.43
R166 A2.n0 A2.t1 241.534
R167 A2.n2 A2.t3 241.437
R168 A2.n0 A2.t0 169.234
R169 A2.n2 A2.t2 169.137
R170 A2.n1 A2.n0 76
R171 A2.n3 A2.n2 76
R172 A2.n1 A2 11.331
R173 A2 A2.n1 7.973
R174 A2 A2.n3 5.102
R175 A2.n3 A2 0.984
R176 a_672_297.n0 a_672_297.t0 627.643
R177 a_672_297.n1 a_672_297.t2 434.219
R178 a_672_297.n2 a_672_297.t3 24.625
R179 a_672_297.n4 a_672_297.n3 14.775
R180 a_672_297.t1 a_672_297.n4 11.82
R181 a_672_297.n1 a_672_297.n0 10.528
R182 a_672_297.n2 a_672_297.n1 9.3
R183 a_672_297.n3 a_672_297.n2 1.97
R184 B1.n0 B1.t0 300.267
R185 B1.n0 B1.t3 221.719
R186 B1.n2 B1.t2 172.626
R187 B1.n1 B1.t1 149.419
R188 B1.n3 B1.n2 76
R189 B1.n2 B1.n1 51.77
R190 B1.n1 B1.n0 17.851
R191 B1.n4 B1 8.32
R192 B1 B1.n4 8.302
R193 B1.n3 B1 1.902
R194 B1.n4 B1.n3 1.556
C0 X VGND 0.45fF
C1 A2 A1 0.31fF
C2 VPWR X 0.62fF
C3 A3 A2 0.11fF
C4 VPB VPWR 0.13fF
C5 VPWR VGND 0.11fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__o31ai_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__o31ai_1 Y A2 A1 A3 B1 VPWR VGND VNB VPB
X0 Y.t1 B1.t0 a_109_47.t1 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 Y.t0 A3.t0 a_193_297.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 a_193_297.t1 A2.t0 a_109_297.t0 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 VGND.t0 A2.t1 a_109_47.t0 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 VPWR.t0 B1.t1 Y.t2 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 a_109_47.t3 A3.t1 VGND.t1 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 a_109_297.t1 A1.t0 VPWR.t1 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 a_109_47.t2 A1.t1 VGND.t2 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
R0 B1.n0 B1.t1 212.079
R1 B1.n0 B1.t0 165.339
R2 B1 B1.n0 117.615
R3 a_109_47.n1 a_109_47.n0 144.391
R4 a_109_47.n0 a_109_47.t1 84.923
R5 a_109_47.n0 a_109_47.t3 27.692
R6 a_109_47.t0 a_109_47.n1 24.923
R7 a_109_47.n1 a_109_47.t2 24.923
R8 Y.n0 Y 302.918
R9 Y.n3 Y.n0 292.5
R10 Y.n0 Y.t0 127.065
R11 Y.n1 Y.t1 82.25
R12 Y.n0 Y.t2 27.58
R13 Y Y.n2 16.669
R14 Y.n3 Y 11.311
R15 Y Y.n3 8.93
R16 Y.n2 Y.n1 6.569
R17 Y.n2 Y 3.572
R18 Y.n1 Y 2.492
R19 Y.n2 Y 1.359
R20 VNB VNB.t2 6053.91
R21 VNB.t3 VNB.t1 3674.73
R22 VNB.t0 VNB.t3 2030.77
R23 VNB.t2 VNB.t0 2030.77
R24 A3.n0 A3.t0 232.471
R25 A3.n0 A3.t1 160.171
R26 A3 A3.n0 77.482
R27 a_193_297.t0 a_193_297.t1 53.19
R28 VPB.t0 VPB.t1 553.426
R29 VPB.t3 VPB.t0 248.598
R30 VPB.t2 VPB.t3 248.598
R31 VPB VPB.t2 189.408
R32 A2.n0 A2.t0 241.534
R33 A2.n0 A2.t1 169.234
R34 A2.n1 A2.n0 76
R35 A2 A2.n1 8.197
R36 A2.n1 A2 1.582
R37 a_109_297.t0 a_109_297.t1 53.19
R38 VGND.n1 VGND.n0 122.715
R39 VGND.n1 VGND.t2 120.431
R40 VGND.n0 VGND.t1 24.923
R41 VGND.n0 VGND.t0 24.923
R42 VGND VGND.n1 0.176
R43 VPWR.n0 VPWR.t0 157.235
R44 VPWR.n0 VPWR.t1 148.487
R45 VPWR VPWR.n0 0.043
R46 A1.n0 A1.t0 230.361
R47 A1.n0 A1.t1 158.061
R48 A1 A1.n0 81.376
C0 VPWR Y 0.20fF
C1 A2 A3 0.18fF
C2 A3 Y 0.15fF
C3 A1 A2 0.10fF
C4 Y VGND 0.13fF
C5 B1 Y 0.13fF
C6 A2 VPWR 0.17fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__o31ai_2.ext - technology: sky130A

.subckt sky130_fd_sc_hd__o31ai_2 A1 Y B1 A3 A2 VGND VPWR VNB VPB
X0 a_281_297.t3 A3.t0 Y.t5 VPB.t7 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_281_297.t0 A2.t0 a_27_297.t1 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 VGND.t1 A2.t1 a_27_47.t1 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 a_27_297.t2 A1.t0 VPWR.t1 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 a_27_47.t2 A1.t1 VGND.t2 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 VGND.t3 A1.t2 a_27_47.t3 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 a_27_47.t7 A3.t1 VGND.t5 VNB.t7 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 VPWR.t2 B1.t0 Y.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 VPWR.t0 A1.t3 a_27_297.t3 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 a_27_47.t4 B1.t1 Y.t1 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 a_27_47.t0 A2.t2 VGND.t0 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 VGND.t4 A3.t2 a_27_47.t6 VNB.t6 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 Y.t2 B1.t2 a_27_47.t5 VNB.t5 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 Y.t4 A3.t3 a_281_297.t2 VPB.t6 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14 Y.t3 B1.t3 VPWR.t3 VPB.t5 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 a_27_297.t0 A2.t3 a_281_297.t1 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
R0 A3.n0 A3.t3 221.719
R1 A3.n2 A3.t0 221.719
R2 A3.n3 A3.t2 161.915
R3 A3.n0 A3.t1 149.419
R4 A3.n1 A3 82.162
R5 A3.n4 A3.n3 76
R6 A3.n2 A3.n1 58.911
R7 A3.n1 A3.n0 16.066
R8 A3 A3.n4 11.851
R9 A3.n4 A3 9.955
R10 A3.n3 A3.n2 1.785
R11 Y.n5 Y.n4 292.5
R12 Y.n4 Y.n3 292.5
R13 Y.n0 Y.t5 174.078
R14 Y.n2 Y.n1 108.41
R15 Y Y.n7 92.887
R16 Y.n2 Y.n0 44.27
R17 Y.n7 Y.t2 39.692
R18 Y.n7 Y.t1 32.307
R19 Y.n4 Y.t3 26.595
R20 Y.n1 Y.t0 26.595
R21 Y.n1 Y.t4 26.595
R22 Y.n6 Y.n5 19.764
R23 Y.n6 Y.n2 12.8
R24 Y.n3 Y 12.047
R25 Y Y.n6 5.236
R26 Y.n0 Y 2.054
R27 Y.n3 Y 0.752
R28 Y.n5 Y 0.752
R29 a_281_297.n1 a_281_297.n0 712.999
R30 a_281_297.n0 a_281_297.t1 26.595
R31 a_281_297.n0 a_281_297.t0 26.595
R32 a_281_297.t2 a_281_297.n1 26.595
R33 a_281_297.n1 a_281_297.t3 26.595
R34 VPB.t4 VPB.t7 568.224
R35 VPB.t0 VPB.t5 319.626
R36 VPB.t6 VPB.t0 248.598
R37 VPB.t7 VPB.t6 248.598
R38 VPB.t3 VPB.t4 248.598
R39 VPB.t1 VPB.t3 248.598
R40 VPB.t2 VPB.t1 248.598
R41 VPB VPB.t2 201.246
R42 A2.n2 A2.t3 221.719
R43 A2.n3 A2.t0 221.719
R44 A2.n0 A2.t2 180.659
R45 A2.n3 A2.t1 149.419
R46 A2.n1 A2.n0 76
R47 A2.n5 A2.n4 76
R48 A2.n4 A2.n3 43.737
R49 A2.n4 A2.n2 31.24
R50 A2.n5 A2.n1 16.118
R51 A2.n1 A2 3.555
R52 A2 A2.n5 2.133
R53 a_27_297.n0 a_27_297.t0 218.348
R54 a_27_297.n0 a_27_297.t3 172.656
R55 a_27_297.n1 a_27_297.n0 108.41
R56 a_27_297.t1 a_27_297.n1 26.595
R57 a_27_297.n1 a_27_297.t2 26.595
R58 a_27_47.n3 a_27_47.t4 219.34
R59 a_27_47.n1 a_27_47.t3 126.698
R60 a_27_47.n4 a_27_47.n1 67.011
R61 a_27_47.n4 a_27_47.n3 60.48
R62 a_27_47.n1 a_27_47.n0 53.206
R63 a_27_47.n5 a_27_47.n4 53.205
R64 a_27_47.n3 a_27_47.n2 43.173
R65 a_27_47.n5 a_27_47.t6 39.692
R66 a_27_47.t0 a_27_47.n5 32.307
R67 a_27_47.n2 a_27_47.t5 24.923
R68 a_27_47.n2 a_27_47.t7 24.923
R69 a_27_47.n0 a_27_47.t1 24.923
R70 a_27_47.n0 a_27_47.t2 24.923
R71 VGND.n11 VGND.n10 114.711
R72 VGND.n1 VGND.n0 109.779
R73 VGND.n3 VGND.n2 92.5
R74 VGND.n5 VGND.n4 92.5
R75 VGND.n0 VGND.t5 39.692
R76 VGND.n2 VGND.t0 24.923
R77 VGND.n4 VGND.t1 24.923
R78 VGND.n0 VGND.t4 24.923
R79 VGND.n10 VGND.t2 24.923
R80 VGND.n10 VGND.t3 24.923
R81 VGND.n6 VGND.n3 5.485
R82 VGND.n12 VGND.n11 4.899
R83 VGND.n7 VGND.n6 4.65
R84 VGND.n9 VGND.n8 4.65
R85 VGND.n6 VGND.n5 1.422
R86 VGND.n7 VGND.n1 0.241
R87 VGND.n12 VGND.n9 0.132
R88 VGND VGND.n12 0.127
R89 VGND.n9 VGND.n7 0.119
R90 VNB VNB.t3 6150.61
R91 VNB.t1 VNB.t0 3674.73
R92 VNB.t5 VNB.t4 2610.99
R93 VNB.t0 VNB.t6 2610.99
R94 VNB.t6 VNB.t7 2417.58
R95 VNB.t7 VNB.t5 2030.77
R96 VNB.t2 VNB.t1 2030.77
R97 VNB.t3 VNB.t2 2030.77
R98 A1.n0 A1.t0 221.719
R99 A1.n2 A1.t3 221.719
R100 A1.n0 A1.t1 149.419
R101 A1.n2 A1.t2 149.419
R102 A1.n3 A1.n2 77.785
R103 A1.n4 A1.n1 76
R104 A1.n2 A1.n1 58.911
R105 A1.n1 A1.n0 16.066
R106 A1.n3 A1 15.644
R107 A1 A1.n4 11.851
R108 A1.n4 A1 9.955
R109 A1 A1.n3 6.162
R110 VPWR.n2 VPWR.n1 178.919
R111 VPWR.n2 VPWR.n0 167.645
R112 VPWR.n0 VPWR.t2 42.355
R113 VPWR.n0 VPWR.t3 34.475
R114 VPWR.n1 VPWR.t1 26.595
R115 VPWR.n1 VPWR.t0 26.595
R116 VPWR VPWR.n2 0.145
R117 B1.n1 B1.t3 212.079
R118 B1.n0 B1.t0 212.079
R119 B1.n1 B1.t1 139.779
R120 B1.n0 B1.t2 139.779
R121 B1 B1.n1 117.506
R122 B1.n1 B1.n0 78.872
C0 VPWR Y 0.40fF
C1 A3 Y 0.22fF
C2 B1 Y 0.16fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__o31ai_4.ext - technology: sky130A

.subckt sky130_fd_sc_hd__o31ai_4 A3 A2 A1 Y B1 VGND VPWR VNB VPB
X0 Y.t11 A3.t0 a_449_297.t7 VPB.t15 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 VPWR.t3 A1.t0 a_27_297.t7 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 a_449_297.t6 A3.t1 Y.t10 VPB.t14 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 Y.t9 A3.t2 a_449_297.t5 VPB.t13 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 VGND.t7 A1.t1 a_31_47.t8 VNB.t8 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 a_27_297.t6 A1.t2 VPWR.t2 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 Y.t0 B1.t0 a_31_47.t0 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 a_449_297.t4 A3.t3 Y.t8 VPB.t12 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 Y.t1 B1.t1 a_31_47.t9 VNB.t9 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 a_31_47.t7 A1.t3 VGND.t6 VNB.t7 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 a_27_297.t0 A2.t0 a_449_297.t0 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 VGND.t5 A1.t4 a_31_47.t6 VNB.t6 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 a_31_47.t5 A1.t5 VGND.t4 VNB.t5 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 Y.t2 B1.t2 VPWR.t4 VPB.t8 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14 a_31_47.t1 A2.t1 VGND.t0 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X15 a_31_47.t2 A2.t2 VGND.t1 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X16 a_449_297.t1 A2.t3 a_27_297.t1 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17 VPWR.t5 B1.t3 Y.t3 VPB.t9 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X18 Y.t4 B1.t4 VPWR.t6 VPB.t10 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X19 VPWR.t1 A1.t6 a_27_297.t5 VPB.t6 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X20 VGND.t2 A2.t4 a_31_47.t3 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X21 VPWR.t7 B1.t5 Y.t5 VPB.t11 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X22 VGND.t3 A2.t5 a_31_47.t4 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X23 VGND.t11 A3.t4 a_31_47.t15 VNB.t15 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X24 a_31_47.t14 A3.t5 VGND.t10 VNB.t14 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X25 a_27_297.t2 A2.t6 a_449_297.t2 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X26 VGND.t9 A3.t6 a_31_47.t13 VNB.t13 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X27 a_31_47.t12 A3.t7 VGND.t8 VNB.t12 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X28 a_449_297.t3 A2.t7 a_27_297.t3 VPB.t5 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X29 a_31_47.t10 B1.t6 Y.t6 VNB.t10 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X30 a_27_297.t4 A1.t7 VPWR.t0 VPB.t7 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X31 a_31_47.t11 B1.t7 Y.t7 VNB.t11 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
R0 A3.n0 A3.t0 221.719
R1 A3.n2 A3.t1 221.719
R2 A3.n12 A3.t2 221.719
R3 A3.n4 A3.t3 221.719
R4 A3.n6 A3.t4 165.485
R5 A3.n0 A3.t7 149.419
R6 A3.n11 A3.t5 149.419
R7 A3.n3 A3.t6 149.419
R8 A3.n15 A3.n1 76
R9 A3.n14 A3.n13 76
R10 A3.n10 A3.n9 76
R11 A3.n8 A3.n7 76
R12 A3.n1 A3.n0 61.588
R13 A3.n7 A3.n6 60.696
R14 A3.n10 A3.n4 41.951
R15 A3.n13 A3.n12 27.67
R16 A3.n13 A3.n3 25.885
R17 A3.n3 A3.n2 21.422
R18 A3.n12 A3.n11 21.422
R19 A3 A3.n15 21.236
R20 A3.n8 A3.n5 19.781
R21 A3.n9 A3 19.49
R22 A3.n7 A3.n4 18.744
R23 A3 A3.n14 14.254
R24 A3.n2 A3.n1 13.388
R25 A3.n14 A3 12.509
R26 A3.n11 A3.n10 11.603
R27 A3.n9 A3 7.272
R28 A3.n5 A3 6.4
R29 A3.n15 A3 5.527
R30 A3 A3.n8 0.29
R31 a_449_297.n4 a_449_297.n3 351.819
R32 a_449_297.n5 a_449_297.n4 292.5
R33 a_449_297.n2 a_449_297.n0 164.17
R34 a_449_297.n2 a_449_297.n1 146.25
R35 a_449_297.n4 a_449_297.n2 57.95
R36 a_449_297.n3 a_449_297.t2 26.595
R37 a_449_297.n3 a_449_297.t3 26.595
R38 a_449_297.n1 a_449_297.t5 26.595
R39 a_449_297.n1 a_449_297.t4 26.595
R40 a_449_297.n0 a_449_297.t7 26.595
R41 a_449_297.n0 a_449_297.t6 26.595
R42 a_449_297.t0 a_449_297.n5 26.595
R43 a_449_297.n5 a_449_297.t1 26.595
R44 Y.n13 Y.t8 473.37
R45 Y.n5 Y.n4 292.5
R46 Y.n6 Y.n5 292.5
R47 Y.n14 Y.n12 292.5
R48 Y.n2 Y.n0 137.3
R49 Y.n9 Y.n8 108.145
R50 Y.n15 Y.n11 108.145
R51 Y.n2 Y.n1 92.5
R52 Y.n12 Y.t10 26.595
R53 Y.n12 Y.t9 26.595
R54 Y.n11 Y.t5 26.595
R55 Y.n11 Y.t11 26.595
R56 Y.n8 Y.t3 26.595
R57 Y.n8 Y.t4 26.595
R58 Y.n5 Y.t2 26.595
R59 Y.n0 Y.t7 24.923
R60 Y.n0 Y.t1 24.923
R61 Y.n1 Y.t6 24.923
R62 Y.n1 Y.t0 24.923
R63 Y.n10 Y 23.524
R64 Y Y.n7 20.736
R65 Y.n10 Y 19.712
R66 Y.n9 Y 17.92
R67 Y.n13 Y 17.664
R68 Y Y.n3 15.221
R69 Y Y.n15 13.824
R70 Y.n14 Y 13.824
R71 Y.n4 Y 11.003
R72 Y.n15 Y 9.728
R73 Y Y.n14 9.728
R74 Y.n3 Y 8.302
R75 Y Y.n9 5.632
R76 Y Y.n13 5.632
R77 Y.n7 Y 5.614
R78 Y.n7 Y.n6 5.389
R79 Y.n4 Y 4.266
R80 Y.n6 Y 4.266
R81 Y.n3 Y.n2 4
R82 Y.n3 Y 4
R83 Y Y.n10 3.84
R84 VPB.t2 VPB.t12 565.264
R85 VPB.t9 VPB.t8 248.598
R86 VPB.t10 VPB.t9 248.598
R87 VPB.t11 VPB.t10 248.598
R88 VPB.t15 VPB.t11 248.598
R89 VPB.t14 VPB.t15 248.598
R90 VPB.t13 VPB.t14 248.598
R91 VPB.t12 VPB.t13 248.598
R92 VPB.t3 VPB.t2 248.598
R93 VPB.t4 VPB.t3 248.598
R94 VPB.t5 VPB.t4 248.598
R95 VPB.t7 VPB.t5 248.598
R96 VPB.t1 VPB.t7 248.598
R97 VPB.t0 VPB.t1 248.598
R98 VPB.t6 VPB.t0 248.598
R99 VPB VPB.t6 204.205
R100 A1.n1 A1.t7 221.719
R101 A1.n2 A1.t0 221.719
R102 A1.n7 A1.t2 221.719
R103 A1.n8 A1.t6 221.719
R104 A1.n1 A1.t5 149.419
R105 A1.n2 A1.t1 149.419
R106 A1.n7 A1.t3 149.419
R107 A1.n8 A1.t4 149.419
R108 A1 A1.n3 78.94
R109 A1.n4 A1.n0 76
R110 A1.n6 A1.n5 76
R111 A1.n10 A1.n9 76
R112 A1.n6 A1.n0 60.696
R113 A1.n9 A1.n7 56.233
R114 A1.n3 A1.n2 50.877
R115 A1.n3 A1.n1 24.1
R116 A1.n9 A1.n8 18.744
R117 A1 A1.n10 15.394
R118 A1.n5 A1 11.243
R119 A1.n2 A1.n0 9.818
R120 A1.n4 A1 8.821
R121 A1 A1.n4 7.091
R122 A1.n5 A1 4.67
R123 A1.n7 A1.n6 4.462
R124 A1.n10 A1 0.518
R125 a_27_297.n6 a_27_297.n5 360.908
R126 a_27_297.n6 a_27_297.t0 178.88
R127 a_27_297.n2 a_27_297.t5 151.723
R128 a_27_297.n5 a_27_297.n4 149.494
R129 a_27_297.n2 a_27_297.n1 103.798
R130 a_27_297.n3 a_27_297.n0 93.013
R131 a_27_297.n5 a_27_297.n3 36.349
R132 a_27_297.n3 a_27_297.n2 32.547
R133 a_27_297.n0 a_27_297.t3 26.595
R134 a_27_297.n0 a_27_297.t4 26.595
R135 a_27_297.n1 a_27_297.t7 26.595
R136 a_27_297.n1 a_27_297.t6 26.595
R137 a_27_297.n4 a_27_297.t1 26.595
R138 a_27_297.n4 a_27_297.t2 26.595
R139 VPWR.n29 VPWR.n28 314.711
R140 VPWR.n23 VPWR.n22 314.711
R141 VPWR.n3 VPWR.n2 166.945
R142 VPWR.n1 VPWR.n0 163.438
R143 VPWR.n2 VPWR.t4 26.595
R144 VPWR.n2 VPWR.t5 26.595
R145 VPWR.n0 VPWR.t6 26.595
R146 VPWR.n0 VPWR.t7 26.595
R147 VPWR.n28 VPWR.t2 26.595
R148 VPWR.n28 VPWR.t1 26.595
R149 VPWR.n22 VPWR.t0 26.595
R150 VPWR.n22 VPWR.t3 26.595
R151 VPWR.n24 VPWR.n23 5.27
R152 VPWR.n30 VPWR.n29 4.899
R153 VPWR.n5 VPWR.n4 4.65
R154 VPWR.n7 VPWR.n6 4.65
R155 VPWR.n9 VPWR.n8 4.65
R156 VPWR.n11 VPWR.n10 4.65
R157 VPWR.n13 VPWR.n12 4.65
R158 VPWR.n15 VPWR.n14 4.65
R159 VPWR.n17 VPWR.n16 4.65
R160 VPWR.n19 VPWR.n18 4.65
R161 VPWR.n21 VPWR.n20 4.65
R162 VPWR.n25 VPWR.n24 4.65
R163 VPWR.n27 VPWR.n26 4.65
R164 VPWR.n3 VPWR.n1 3.683
R165 VPWR.n5 VPWR.n3 0.255
R166 VPWR.n30 VPWR.n27 0.132
R167 VPWR VPWR.n30 0.129
R168 VPWR.n7 VPWR.n5 0.119
R169 VPWR.n9 VPWR.n7 0.119
R170 VPWR.n11 VPWR.n9 0.119
R171 VPWR.n13 VPWR.n11 0.119
R172 VPWR.n15 VPWR.n13 0.119
R173 VPWR.n17 VPWR.n15 0.119
R174 VPWR.n19 VPWR.n17 0.119
R175 VPWR.n21 VPWR.n19 0.119
R176 VPWR.n25 VPWR.n21 0.119
R177 VPWR.n27 VPWR.n25 0.119
R178 a_31_47.n11 a_31_47.t11 133.874
R179 a_31_47.n2 a_31_47.t6 129.504
R180 a_31_47.n9 a_31_47.n0 104.17
R181 a_31_47.n11 a_31_47.n10 92.5
R182 a_31_47.n13 a_31_47.n12 92.5
R183 a_31_47.n12 a_31_47.n9 83.952
R184 a_31_47.n9 a_31_47.n8 82.07
R185 a_31_47.n12 a_31_47.n11 55.272
R186 a_31_47.n2 a_31_47.n1 53.206
R187 a_31_47.n4 a_31_47.n3 53.206
R188 a_31_47.n6 a_31_47.n5 53.206
R189 a_31_47.n8 a_31_47.n7 53.206
R190 a_31_47.n4 a_31_47.n2 38.4
R191 a_31_47.n6 a_31_47.n4 38.4
R192 a_31_47.n8 a_31_47.n6 38.4
R193 a_31_47.n1 a_31_47.t8 24.923
R194 a_31_47.n1 a_31_47.t7 24.923
R195 a_31_47.n3 a_31_47.t3 24.923
R196 a_31_47.n3 a_31_47.t5 24.923
R197 a_31_47.n5 a_31_47.t4 24.923
R198 a_31_47.n5 a_31_47.t1 24.923
R199 a_31_47.n7 a_31_47.t15 24.923
R200 a_31_47.n7 a_31_47.t2 24.923
R201 a_31_47.n0 a_31_47.t13 24.923
R202 a_31_47.n0 a_31_47.t14 24.923
R203 a_31_47.n10 a_31_47.t9 24.923
R204 a_31_47.n10 a_31_47.t10 24.923
R205 a_31_47.t0 a_31_47.n13 24.923
R206 a_31_47.n13 a_31_47.t12 24.923
R207 VGND.n13 VGND.n12 114.711
R208 VGND.n17 VGND.n16 114.711
R209 VGND.n23 VGND.n22 114.711
R210 VGND.n29 VGND.n28 114.711
R211 VGND.n1 VGND.n0 96.612
R212 VGND.n3 VGND.n2 92.5
R213 VGND.n5 VGND.n4 92.5
R214 VGND.n4 VGND.t11 38.769
R215 VGND.n0 VGND.t8 36
R216 VGND.n0 VGND.t9 36
R217 VGND.n2 VGND.t10 24.923
R218 VGND.n12 VGND.t1 24.923
R219 VGND.n12 VGND.t3 24.923
R220 VGND.n16 VGND.t0 24.923
R221 VGND.n16 VGND.t2 24.923
R222 VGND.n22 VGND.t4 24.923
R223 VGND.n22 VGND.t7 24.923
R224 VGND.n28 VGND.t6 24.923
R225 VGND.n28 VGND.t5 24.923
R226 VGND.n14 VGND.n13 17.317
R227 VGND.n18 VGND.n17 11.294
R228 VGND.n24 VGND.n23 5.27
R229 VGND.n30 VGND.n29 4.899
R230 VGND.n6 VGND.n5 4.774
R231 VGND.n7 VGND.n6 4.65
R232 VGND.n9 VGND.n8 4.65
R233 VGND.n11 VGND.n10 4.65
R234 VGND.n15 VGND.n14 4.65
R235 VGND.n19 VGND.n18 4.65
R236 VGND.n21 VGND.n20 4.65
R237 VGND.n25 VGND.n24 4.65
R238 VGND.n27 VGND.n26 4.65
R239 VGND.n6 VGND.n3 2.133
R240 VGND.n7 VGND.n1 0.597
R241 VGND.n30 VGND.n27 0.132
R242 VGND VGND.n30 0.129
R243 VGND.n9 VGND.n7 0.119
R244 VGND.n11 VGND.n9 0.119
R245 VGND.n15 VGND.n11 0.119
R246 VGND.n19 VGND.n15 0.119
R247 VGND.n21 VGND.n19 0.119
R248 VGND.n25 VGND.n21 0.119
R249 VGND.n27 VGND.n25 0.119
R250 VNB VNB.t6 6174.79
R251 VNB.t15 VNB.t14 4037.36
R252 VNB.t13 VNB.t12 2610.99
R253 VNB.t9 VNB.t11 2030.77
R254 VNB.t10 VNB.t9 2030.77
R255 VNB.t0 VNB.t10 2030.77
R256 VNB.t12 VNB.t0 2030.77
R257 VNB.t14 VNB.t13 2030.77
R258 VNB.t2 VNB.t15 2030.77
R259 VNB.t4 VNB.t2 2030.77
R260 VNB.t1 VNB.t4 2030.77
R261 VNB.t3 VNB.t1 2030.77
R262 VNB.t5 VNB.t3 2030.77
R263 VNB.t8 VNB.t5 2030.77
R264 VNB.t7 VNB.t8 2030.77
R265 VNB.t6 VNB.t7 2030.77
R266 B1.n0 B1.t2 221.719
R267 B1.n3 B1.t3 221.719
R268 B1.n7 B1.t4 221.719
R269 B1.n6 B1.t5 221.719
R270 B1.n0 B1.t7 149.419
R271 B1.n3 B1.t1 149.419
R272 B1.n7 B1.t6 149.419
R273 B1.n6 B1.t0 149.419
R274 B1.n2 B1.n1 76
R275 B1.n5 B1.n4 76
R276 B1.n9 B1.n8 76
R277 B1.n7 B1.n6 74.977
R278 B1.n4 B1.n2 60.696
R279 B1.n8 B1.n7 25.885
R280 B1.n9 B1.n5 19.781
R281 B1.n1 B1 15.418
R282 B1.n4 B1.n3 11.603
R283 B1.n1 B1 11.345
R284 B1.n5 B1 4.363
R285 B1.n2 B1.n0 2.677
R286 B1 B1.n9 2.618
R287 A2.n0 A2.t0 221.719
R288 A2.n2 A2.t3 221.719
R289 A2.n8 A2.t6 221.719
R290 A2.n9 A2.t7 221.719
R291 A2.n0 A2.t2 149.419
R292 A2.n2 A2.t5 149.419
R293 A2.n8 A2.t1 149.419
R294 A2.n9 A2.t4 149.419
R295 A2.n5 A2.n3 76
R296 A2.n7 A2.n6 76
R297 A2.n11 A2.n10 76
R298 A2.n7 A2.n3 60.696
R299 A2.n10 A2.n8 58.911
R300 A2.n2 A2.n1 48.2
R301 A2.n1 A2.n0 26.777
R302 A2.n10 A2.n9 16.066
R303 A2.n3 A2.n2 12.496
R304 A2.n5 A2.n4 11.762
R305 A2.n6 A2 10.724
R306 A2 A2.n11 9.34
R307 A2.n11 A2 6.572
R308 A2.n6 A2 5.189
R309 A2.n4 A2 3.113
R310 A2.n8 A2.n7 1.785
R311 A2 A2.n5 1.037
C0 VPB VPWR 0.15fF
C1 VPWR VGND 0.16fF
C2 A3 Y 0.40fF
C3 A1 A2 0.12fF
C4 B1 Y 0.42fF
C5 VPWR Y 0.60fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__o32a_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__o32a_1 X A3 A1 A2 B1 B2 VPWR VGND VNB VPB
X0 a_77_199.t1 B2.t0 a_227_47.t3 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 a_323_297.t0 A2.t0 a_227_297.t0 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 a_227_297.t1 A1.t0 VPWR.t1 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 a_227_47.t2 B1.t0 a_77_199.t0 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 VGND.t1 a_77_199.t4 X.t1 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 VPWR.t2 B1.t1 a_539_297.t0 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 a_227_47.t0 A3.t0 VGND.t0 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 VPWR.t0 a_77_199.t5 X.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 a_77_199.t3 A3.t1 a_323_297.t1 VPB.t5 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 VGND.t2 A2.t1 a_227_47.t1 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 a_227_47.t4 A1.t1 VGND.t3 VNB.t5 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 a_539_297.t1 B2.t1 a_77_199.t2 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
R0 B2.n0 B2.t1 236.179
R1 B2.n0 B2.t0 163.879
R2 B2.n1 B2.n0 76
R3 B2.n1 B2 10.276
R4 B2 B2.n1 1.983
R5 a_227_47.n1 a_227_47.t2 222.807
R6 a_227_47.n1 a_227_47.n0 112.751
R7 a_227_47.n2 a_227_47.n1 43.173
R8 a_227_47.t0 a_227_47.n2 40.615
R9 a_227_47.n0 a_227_47.t4 31.384
R10 a_227_47.n2 a_227_47.t3 31.384
R11 a_227_47.n0 a_227_47.t1 29.538
R12 a_77_199.n2 a_77_199.n0 259.573
R13 a_77_199.n0 a_77_199.t5 236.179
R14 a_77_199.n2 a_77_199.n1 215.984
R15 a_77_199.n0 a_77_199.t4 163.879
R16 a_77_199.n3 a_77_199.n2 143.027
R17 a_77_199.n1 a_77_199.t0 42.461
R18 a_77_199.t2 a_77_199.n3 39.4
R19 a_77_199.n3 a_77_199.t3 37.43
R20 a_77_199.n1 a_77_199.t1 33.23
R21 VNB VNB.t1 6985.92
R22 VNB.t4 VNB.t3 2707.69
R23 VNB.t0 VNB.t4 2610.99
R24 VNB.t2 VNB.t0 2610.99
R25 VNB.t5 VNB.t2 2320.88
R26 VNB.t1 VNB.t5 2030.77
R27 A2.n0 A2.t0 236.179
R28 A2.n0 A2.t1 163.879
R29 A2.n1 A2.n0 76
R30 A2 A2.n1 10.847
R31 A2.n1 A2 2.04
R32 a_227_297.t0 a_227_297.t1 65.01
R33 a_323_297.t0 a_323_297.t1 76.83
R34 VPB.t3 VPB.t4 331.464
R35 VPB.t5 VPB.t3 319.626
R36 VPB.t1 VPB.t5 319.626
R37 VPB VPB.t0 295.95
R38 VPB.t2 VPB.t1 284.112
R39 VPB.t0 VPB.t2 248.598
R40 A1.n0 A1.t0 236.179
R41 A1.n0 A1.t1 163.879
R42 A1 A1.n0 78.816
R43 VPWR.n1 VPWR.n0 170.001
R44 VPWR.n1 VPWR.t2 153.481
R45 VPWR.n0 VPWR.t1 26.595
R46 VPWR.n0 VPWR.t0 26.595
R47 VPWR VPWR.n1 0.158
R48 B1.n0 B1.t1 229.182
R49 B1.n0 B1.t0 156.882
R50 B1 B1.n0 78.56
R51 X.t0 X 477.343
R52 X.n1 X.t0 424.813
R53 X.n0 X.t1 83.875
R54 X.n1 X.n0 63.964
R55 X.n0 X 3.733
R56 X X.n1 0.831
R57 VGND.n2 VGND.n0 124.645
R58 VGND.n2 VGND.n1 111.563
R59 VGND.n1 VGND.t0 36
R60 VGND.n1 VGND.t2 36
R61 VGND.n0 VGND.t3 24.923
R62 VGND.n0 VGND.t1 24.923
R63 VGND VGND.n2 0.301
R64 a_539_297.t0 a_539_297.t1 80.77
R65 A3.n0 A3.t1 236.179
R66 A3.n0 A3.t0 163.879
R67 A3.n1 A3.n0 76
R68 A3.n1 A3 13.265
R69 A3 A3.n1 2.56
C0 X VPWR 0.14fF
C1 A3 B2 0.15fF
C2 VGND X 0.15fF
C3 A2 A3 0.13fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__o32a_2.ext - technology: sky130A

.subckt sky130_fd_sc_hd__o32a_2 B1 B2 A3 A2 A1 X VGND VPWR VNB VPB
X0 a_429_297.t1 A2.t0 a_345_297.t1 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 VGND.t3 A2.t1 a_345_47.t3 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 VPWR.t3 a_79_21.t4 X.t3 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 VGND.t0 a_79_21.t5 X.t1 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 a_345_47.t0 A3.t0 VGND.t1 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 a_345_297.t0 A1.t0 VPWR.t0 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 a_629_297.t0 B2.t0 a_79_21.t2 VPB.t5 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 VPWR.t1 B1.t0 a_629_297.t1 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 a_79_21.t3 B2.t1 a_345_47.t4 VNB.t5 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 a_345_47.t2 B1.t1 a_79_21.t1 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 a_79_21.t0 A3.t1 a_429_297.t0 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 X.t2 a_79_21.t6 VPWR.t2 VPB.t6 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 X.t0 a_79_21.t7 VGND.t4 VNB.t6 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 a_345_47.t1 A1.t1 VGND.t2 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
R0 A2.n0 A2.t0 241.534
R1 A2.n0 A2.t1 169.234
R2 A2 A2.n0 77.651
R3 a_345_297.t0 a_345_297.t1 53.19
R4 a_429_297.t0 a_429_297.t1 84.71
R5 VPB.t0 VPB.t2 449.844
R6 VPB.t4 VPB.t1 343.302
R7 VPB.t5 VPB.t3 313.707
R8 VPB.t1 VPB.t5 248.598
R9 VPB.t2 VPB.t4 248.598
R10 VPB.t6 VPB.t0 248.598
R11 VPB VPB.t6 189.408
R12 a_345_47.n1 a_345_47.t2 139.74
R13 a_345_47.n1 a_345_47.n0 107.481
R14 a_345_47.n2 a_345_47.n1 43.173
R15 a_345_47.n0 a_345_47.t3 24.923
R16 a_345_47.n0 a_345_47.t1 24.923
R17 a_345_47.n2 a_345_47.t4 24.923
R18 a_345_47.t0 a_345_47.n2 24.923
R19 VGND.n3 VGND.n2 110.882
R20 VGND.n6 VGND.t4 108.334
R21 VGND.n1 VGND.n0 64.067
R22 VGND.n0 VGND.t2 58.153
R23 VGND.n0 VGND.t0 54.461
R24 VGND.n2 VGND.t1 39.692
R25 VGND.n2 VGND.t3 39.692
R26 VGND.n7 VGND.n6 4.65
R27 VGND.n5 VGND.n4 4.65
R28 VGND.n3 VGND.n1 3.652
R29 VGND.n5 VGND.n3 0.172
R30 VGND.n7 VGND.n5 0.119
R31 VGND VGND.n7 0.02
R32 VNB VNB.t6 6053.91
R33 VNB.t0 VNB.t2 3674.73
R34 VNB.t4 VNB.t1 2804.4
R35 VNB.t5 VNB.t3 2562.64
R36 VNB.t1 VNB.t5 2030.77
R37 VNB.t2 VNB.t4 2030.77
R38 VNB.t6 VNB.t0 2030.77
R39 a_79_21.n3 a_79_21.n1 239.14
R40 a_79_21.n1 a_79_21.t4 212.079
R41 a_79_21.n0 a_79_21.t6 212.079
R42 a_79_21.n3 a_79_21.n2 186.04
R43 a_79_21.n4 a_79_21.n3 154.518
R44 a_79_21.n1 a_79_21.t5 139.779
R45 a_79_21.n0 a_79_21.t7 139.779
R46 a_79_21.n1 a_79_21.n0 61.345
R47 a_79_21.n2 a_79_21.t3 39.692
R48 a_79_21.n2 a_79_21.t1 30.461
R49 a_79_21.n4 a_79_21.t2 26.595
R50 a_79_21.t0 a_79_21.n4 26.595
R51 X.n3 X.n2 292.5
R52 X.n4 X.n3 147.104
R53 X X.n0 94.245
R54 X.n1 X.n0 92.5
R55 X.n3 X.t3 26.595
R56 X.n3 X.t2 26.595
R57 X.n0 X.t1 24.923
R58 X.n0 X.t0 24.923
R59 X.n1 X 11.442
R60 X.n4 X 10.71
R61 X.n2 X 8.339
R62 X.n2 X 4.848
R63 X X.n4 2.439
R64 X X.n1 1.745
R65 VPWR.n4 VPWR.n3 292.5
R66 VPWR.n2 VPWR.n1 292.5
R67 VPWR.n9 VPWR.t2 151.631
R68 VPWR.n0 VPWR.t1 148.473
R69 VPWR.n1 VPWR.t0 26.595
R70 VPWR.n3 VPWR.t3 26.595
R71 VPWR.n5 VPWR.n2 5.458
R72 VPWR.n6 VPWR.n5 4.65
R73 VPWR.n8 VPWR.n7 4.65
R74 VPWR.n10 VPWR.n9 4.65
R75 VPWR.n5 VPWR.n4 0.941
R76 VPWR.n6 VPWR.n0 0.134
R77 VPWR.n8 VPWR.n6 0.119
R78 VPWR.n10 VPWR.n8 0.119
R79 VPWR VPWR.n10 0.02
R80 A3.n0 A3.t1 237.733
R81 A3.n0 A3.t0 165.433
R82 A3 A3.n0 78.064
R83 A1.n0 A1.t0 240.482
R84 A1.n0 A1.t1 168.182
R85 A1 A1.n0 79.2
R86 B2.n0 B2.t0 241.534
R87 B2.n0 B2.t1 169.234
R88 B2 B2.n0 79.303
R89 a_629_297.t0 a_629_297.t1 74.86
R90 B1.n0 B1.t0 232.209
R91 B1.n0 B1.t1 159.909
R92 B1 B1.n0 77.536
C0 A2 A3 0.12fF
C1 VPWR X 0.26fF
C2 A1 A2 0.12fF
C3 VPWR VGND 0.11fF
C4 X VGND 0.23fF
C5 A3 B2 0.12fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__o32a_4.ext - technology: sky130A

.subckt sky130_fd_sc_hd__o32a_4 X B2 A1 A2 A3 B1 VGND VPWR VNB VPB
X0 a_27_47.t5 B2.t0 a_549_297.t5 VNB.t9 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 VGND.t3 a_549_297.t8 X.t7 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 VPWR.t3 a_549_297.t9 X.t3 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 a_27_297.t2 A2.t0 a_277_297.t3 VPB.t8 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 a_277_297.t2 A2.t1 a_27_297.t1 VPB.t12 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 a_549_297.t7 B2.t1 a_739_297.t3 VPB.t10 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 a_27_47.t2 A3.t0 VGND.t4 VNB.t6 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 a_27_297.t0 A1.t0 VPWR.t6 VPB.t11 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 a_739_297.t2 B2.t2 a_549_297.t6 VPB.t9 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 a_739_297.t0 B1.t0 VPWR.t4 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 a_27_47.t8 A1.t1 VGND.t8 VNB.t12 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 a_27_47.t6 A2.t2 VGND.t6 VNB.t10 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 a_549_297.t4 B2.t3 a_27_47.t4 VNB.t8 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 a_277_297.t0 A3.t1 a_549_297.t2 VPB.t6 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14 VPWR.t5 B1.t1 a_739_297.t1 VPB.t5 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 X.t2 a_549_297.t10 VPWR.t2 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16 a_27_47.t0 B1.t2 a_549_297.t0 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X17 a_549_297.t3 A3.t2 a_277_297.t1 VPB.t7 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X18 VGND.t5 A3.t3 a_27_47.t3 VNB.t7 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X19 VPWR.t1 a_549_297.t11 X.t1 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X20 VGND.t2 a_549_297.t12 X.t6 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X21 VGND.t7 A2.t3 a_27_47.t7 VNB.t11 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X22 X.t0 a_549_297.t13 VPWR.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X23 a_549_297.t1 B1.t3 a_27_47.t1 VNB.t5 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X24 X.t5 a_549_297.t14 VGND.t1 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X25 X.t4 a_549_297.t15 VGND.t0 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X26 VPWR.t7 A1.t2 a_27_297.t3 VPB.t13 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X27 VGND.t9 A1.t3 a_27_47.t9 VNB.t13 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
R0 B2.n0 B2.t2 221.719
R1 B2.n1 B2.t1 221.719
R2 B2.n0 B2.t3 149.419
R3 B2.n1 B2.t0 149.419
R4 B2 B2.n2 95.52
R5 B2.n2 B2.n0 40.166
R6 B2.n2 B2.n1 40.166
R7 a_549_297.n16 a_549_297.n15 425.056
R8 a_549_297.n14 a_549_297.n13 401.744
R9 a_549_297.n0 a_549_297.t9 221.719
R10 a_549_297.n2 a_549_297.t10 221.719
R11 a_549_297.n5 a_549_297.t11 221.719
R12 a_549_297.n8 a_549_297.t13 221.719
R13 a_549_297.n15 a_549_297.t0 166.346
R14 a_549_297.n10 a_549_297.t4 166.346
R15 a_549_297.n0 a_549_297.t8 149.419
R16 a_549_297.n2 a_549_297.t15 149.419
R17 a_549_297.n5 a_549_297.t12 149.419
R18 a_549_297.n8 a_549_297.t14 149.419
R19 a_549_297.n9 a_549_297.n8 112.596
R20 a_549_297.n4 a_549_297.n1 107.623
R21 a_549_297.n12 a_549_297.n11 92.5
R22 a_549_297.n4 a_549_297.n3 76
R23 a_549_297.n7 a_549_297.n6 76
R24 a_549_297.n12 a_549_297.n10 64.752
R25 a_549_297.n15 a_549_297.n14 43.67
R26 a_549_297.n10 a_549_297.n9 41.451
R27 a_549_297.n1 a_549_297.n0 37.488
R28 a_549_297.n3 a_549_297.n2 37.488
R29 a_549_297.n6 a_549_297.n5 37.488
R30 a_549_297.n13 a_549_297.t7 32.505
R31 a_549_297.n7 a_549_297.n4 31.623
R32 a_549_297.n9 a_549_297.n7 30.612
R33 a_549_297.n13 a_549_297.t6 26.595
R34 a_549_297.t2 a_549_297.n16 26.595
R35 a_549_297.n16 a_549_297.t3 26.595
R36 a_549_297.n11 a_549_297.t5 24.923
R37 a_549_297.n11 a_549_297.t1 24.923
R38 a_549_297.n14 a_549_297.n12 3.011
R39 a_27_47.n3 a_27_47.t9 168.632
R40 a_27_47.n7 a_27_47.n6 145.528
R41 a_27_47.n5 a_27_47.t2 117.423
R42 a_27_47.n4 a_27_47.n1 92.5
R43 a_27_47.n3 a_27_47.n2 92.5
R44 a_27_47.n6 a_27_47.n0 92.5
R45 a_27_47.n6 a_27_47.n5 85.138
R46 a_27_47.n5 a_27_47.n4 51.712
R47 a_27_47.n4 a_27_47.n3 44.032
R48 a_27_47.t5 a_27_47.n7 30.461
R49 a_27_47.n1 a_27_47.t6 28.615
R50 a_27_47.n0 a_27_47.t1 24.923
R51 a_27_47.n0 a_27_47.t0 24.923
R52 a_27_47.n2 a_27_47.t7 24.923
R53 a_27_47.n2 a_27_47.t8 24.923
R54 a_27_47.n1 a_27_47.t3 24.923
R55 a_27_47.n7 a_27_47.t4 24.923
R56 VNB.t6 VNB.t4 6962.64
R57 VNB VNB.t13 6053.91
R58 VNB.t8 VNB.t1 4545.05
R59 VNB.t9 VNB.t8 2175.82
R60 VNB.t10 VNB.t7 2127.47
R61 VNB.t0 VNB.t3 2030.77
R62 VNB.t2 VNB.t0 2030.77
R63 VNB.t1 VNB.t2 2030.77
R64 VNB.t5 VNB.t9 2030.77
R65 VNB.t4 VNB.t5 2030.77
R66 VNB.t7 VNB.t6 2030.77
R67 VNB.t11 VNB.t10 2030.77
R68 VNB.t12 VNB.t11 2030.77
R69 VNB.t13 VNB.t12 2030.77
R70 X.n5 X.n3 146.035
R71 X.n5 X.n4 107.635
R72 X.n2 X.n0 87.175
R73 X.n2 X.n1 52.818
R74 X.n3 X.t1 26.595
R75 X.n3 X.t0 26.595
R76 X.n4 X.t3 26.595
R77 X.n4 X.t2 26.595
R78 X.n0 X.t6 24.923
R79 X.n0 X.t5 24.923
R80 X.n1 X.t7 24.923
R81 X.n1 X.t4 24.923
R82 X X.n5 16.326
R83 X.n6 X.n2 11.452
R84 X.n6 X 7.706
R85 X X.n6 1.175
R86 VGND.n0 VGND.t3 199.891
R87 VGND.n2 VGND.n1 114.711
R88 VGND.n5 VGND.t1 113.911
R89 VGND.n23 VGND.n22 92.5
R90 VGND.n29 VGND.n28 92.5
R91 VGND.n35 VGND.n34 92.5
R92 VGND.n34 VGND.t8 24.923
R93 VGND.n34 VGND.t9 24.923
R94 VGND.n28 VGND.t6 24.923
R95 VGND.n28 VGND.t7 24.923
R96 VGND.n22 VGND.t4 24.923
R97 VGND.n22 VGND.t5 24.923
R98 VGND.n1 VGND.t0 24.923
R99 VGND.n1 VGND.t2 24.923
R100 VGND.n3 VGND.n2 16.564
R101 VGND.n6 VGND.n5 12.047
R102 VGND.n37 VGND.n36 4.65
R103 VGND.n27 VGND.n26 4.65
R104 VGND.n31 VGND.n30 4.65
R105 VGND.n33 VGND.n32 4.65
R106 VGND.n4 VGND.n3 4.65
R107 VGND.n7 VGND.n6 4.65
R108 VGND.n9 VGND.n8 4.65
R109 VGND.n11 VGND.n10 4.65
R110 VGND.n13 VGND.n12 4.65
R111 VGND.n15 VGND.n14 4.65
R112 VGND.n17 VGND.n16 4.65
R113 VGND.n19 VGND.n18 4.65
R114 VGND.n21 VGND.n20 4.65
R115 VGND.n25 VGND.n24 4.65
R116 VGND.n24 VGND.n23 3.49
R117 VGND.n30 VGND.n29 2.094
R118 VGND.n4 VGND.n0 0.456
R119 VGND.n36 VGND.n35 0.232
R120 VGND.n7 VGND.n4 0.119
R121 VGND.n9 VGND.n7 0.119
R122 VGND.n11 VGND.n9 0.119
R123 VGND.n13 VGND.n11 0.119
R124 VGND.n15 VGND.n13 0.119
R125 VGND.n17 VGND.n15 0.119
R126 VGND.n19 VGND.n17 0.119
R127 VGND.n21 VGND.n19 0.119
R128 VGND.n25 VGND.n21 0.119
R129 VGND.n27 VGND.n25 0.119
R130 VGND.n31 VGND.n27 0.119
R131 VGND.n33 VGND.n31 0.119
R132 VGND.n37 VGND.n33 0.119
R133 VGND.n38 VGND.n37 0.119
R134 VGND VGND.n38 0.02
R135 VPWR.n15 VPWR.n14 318.476
R136 VPWR.n0 VPWR.t3 201.307
R137 VPWR.n5 VPWR.t0 201.189
R138 VPWR.n33 VPWR.n32 174.594
R139 VPWR.n2 VPWR.n1 174.594
R140 VPWR.n32 VPWR.t6 26.595
R141 VPWR.n32 VPWR.t7 26.595
R142 VPWR.n14 VPWR.t4 26.595
R143 VPWR.n14 VPWR.t5 26.595
R144 VPWR.n1 VPWR.t2 26.595
R145 VPWR.n1 VPWR.t1 26.595
R146 VPWR.n3 VPWR.n2 16.564
R147 VPWR.n6 VPWR.n5 12.047
R148 VPWR.n16 VPWR.n15 9.788
R149 VPWR.n35 VPWR.n34 4.65
R150 VPWR.n4 VPWR.n3 4.65
R151 VPWR.n7 VPWR.n6 4.65
R152 VPWR.n9 VPWR.n8 4.65
R153 VPWR.n11 VPWR.n10 4.65
R154 VPWR.n13 VPWR.n12 4.65
R155 VPWR.n17 VPWR.n16 4.65
R156 VPWR.n19 VPWR.n18 4.65
R157 VPWR.n21 VPWR.n20 4.65
R158 VPWR.n23 VPWR.n22 4.65
R159 VPWR.n25 VPWR.n24 4.65
R160 VPWR.n27 VPWR.n26 4.65
R161 VPWR.n29 VPWR.n28 4.65
R162 VPWR.n31 VPWR.n30 4.65
R163 VPWR.n34 VPWR.n33 0.752
R164 VPWR.n4 VPWR.n0 0.456
R165 VPWR.n7 VPWR.n4 0.119
R166 VPWR.n9 VPWR.n7 0.119
R167 VPWR.n11 VPWR.n9 0.119
R168 VPWR.n13 VPWR.n11 0.119
R169 VPWR.n17 VPWR.n13 0.119
R170 VPWR.n19 VPWR.n17 0.119
R171 VPWR.n21 VPWR.n19 0.119
R172 VPWR.n23 VPWR.n21 0.119
R173 VPWR.n25 VPWR.n23 0.119
R174 VPWR.n27 VPWR.n25 0.119
R175 VPWR.n29 VPWR.n27 0.119
R176 VPWR.n31 VPWR.n29 0.119
R177 VPWR.n35 VPWR.n31 0.119
R178 VPWR.n36 VPWR.n35 0.119
R179 VPWR VPWR.n36 0.02
R180 VPB.t9 VPB.t0 556.386
R181 VPB.t6 VPB.t5 556.386
R182 VPB.t8 VPB.t7 556.386
R183 VPB.t10 VPB.t9 266.355
R184 VPB.t2 VPB.t3 248.598
R185 VPB.t1 VPB.t2 248.598
R186 VPB.t0 VPB.t1 248.598
R187 VPB.t4 VPB.t10 248.598
R188 VPB.t5 VPB.t4 248.598
R189 VPB.t7 VPB.t6 248.598
R190 VPB.t12 VPB.t8 248.598
R191 VPB.t11 VPB.t12 248.598
R192 VPB.t13 VPB.t11 248.598
R193 VPB VPB.t13 189.408
R194 A2.n0 A2.t0 221.719
R195 A2.n1 A2.t1 221.719
R196 A2.n0 A2.t2 149.419
R197 A2.n1 A2.t3 149.419
R198 A2 A2.n2 76.32
R199 A2.n2 A2.n1 40.166
R200 A2.n2 A2.n0 34.811
R201 a_277_297.n1 a_277_297.n0 362.468
R202 a_277_297.t0 a_277_297.n1 185.249
R203 a_277_297.n1 a_277_297.t1 118.508
R204 a_277_297.n0 a_277_297.t3 26.595
R205 a_277_297.n0 a_277_297.t2 26.595
R206 a_27_297.t2 a_27_297.n1 230.19
R207 a_27_297.n1 a_27_297.t3 181.244
R208 a_27_297.n1 a_27_297.n0 91.913
R209 a_27_297.n0 a_27_297.t1 26.595
R210 a_27_297.n0 a_27_297.t0 26.595
R211 a_739_297.t2 a_739_297.n1 178.691
R212 a_739_297.n1 a_739_297.t1 178.549
R213 a_739_297.n1 a_739_297.n0 143.026
R214 a_739_297.n0 a_739_297.t3 26.595
R215 a_739_297.n0 a_739_297.t0 26.595
R216 A3.n0 A3.t1 296.696
R217 A3.n0 A3.t2 221.719
R218 A3.n2 A3.t3 165.485
R219 A3.n1 A3.t0 149.419
R220 A3 A3.n2 92
R221 A3.n2 A3.n1 58.911
R222 A3.n1 A3.n0 14.281
R223 A1.n0 A1.t0 221.719
R224 A1.n1 A1.t2 221.719
R225 A1.n0 A1.t1 149.419
R226 A1.n1 A1.t3 149.419
R227 A1.n2 A1.n1 76.892
R228 A1.n1 A1.n0 74.977
R229 A1 A1.n2 20.16
R230 A1.n2 A1 9.28
R231 B1.n0 B1.t0 221.719
R232 B1.n1 B1.t1 221.719
R233 B1.n0 B1.t3 149.419
R234 B1.n1 B1.t2 149.419
R235 B1 B1.n2 88.48
R236 B1.n2 B1.n0 68.729
R237 B1.n2 B1.n1 6.248
C0 X VGND 0.51fF
C1 VPB VPWR 0.17fF
C2 VPWR X 0.67fF
C3 VPWR VGND 0.17fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__o32ai_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__o32ai_1 A2 Y A1 A3 B2 B1 VGND VPWR VNB VPB
X0 VGND.t1 A3.t0 a_27_47.t2 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 a_27_47.t3 A2.t0 VGND.t2 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 Y.t0 B2.t0 a_109_297.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 a_333_297.t1 A3.t1 Y.t2 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 VGND.t0 A1.t0 a_27_47.t1 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 a_27_47.t0 B2.t1 Y.t1 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 VPWR.t0 A1.t1 a_461_297.t1 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 a_109_297.t1 B1.t0 VPWR.t1 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 a_461_297.t0 A2.t1 a_333_297.t0 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 Y.t3 B1.t1 a_27_47.t4 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
R0 A3.n0 A3.t1 235.819
R1 A3.n0 A3.t0 215.418
R2 A3 A3.n0 78.427
R3 a_27_47.n1 a_27_47.t4 224.136
R4 a_27_47.n1 a_27_47.n0 190.536
R5 a_27_47.n2 a_27_47.n1 43.173
R6 a_27_47.t0 a_27_47.n2 29.538
R7 a_27_47.n2 a_27_47.t2 27.692
R8 a_27_47.n0 a_27_47.t1 24.923
R9 a_27_47.n0 a_27_47.t3 24.923
R10 VGND.n1 VGND.n0 92.5
R11 VGND.n4 VGND.n3 92.5
R12 VGND.n2 VGND.t0 91.774
R13 VGND.n3 VGND.t1 36.923
R14 VGND.n0 VGND.t2 24.923
R15 VGND.n5 VGND.n4 5.644
R16 VGND.n2 VGND.n1 5.045
R17 VGND VGND.n5 0.362
R18 VGND.n5 VGND.n2 0.279
R19 VNB VNB.t4 6053.91
R20 VNB.t2 VNB.t3 3989.01
R21 VNB.t4 VNB.t0 2296.7
R22 VNB.t0 VNB.t2 2224.18
R23 VNB.t3 VNB.t1 2030.77
R24 A2.n0 A2.t1 236.179
R25 A2.n0 A2.t0 163.879
R26 A2.n1 A2.n0 76
R27 A2.n1 A2 12.366
R28 A2 A2.n1 2.386
R29 B2.n0 B2.t0 233.868
R30 B2.n0 B2.t1 162.548
R31 B2 B2.n0 78.374
R32 a_109_297.t0 a_109_297.t1 41.37
R33 Y.n2 Y.n0 168.078
R34 Y.n1 Y.t2 60.085
R35 Y.n1 Y.t0 60.085
R36 Y.n0 Y.t1 35.076
R37 Y.n0 Y.t3 24.923
R38 Y.n2 Y 8.564
R39 Y Y.n1 2.635
R40 Y Y.n2 0.094
R41 VPB.t0 VPB.t2 449.844
R42 VPB.t2 VPB.t1 378.816
R43 VPB.t1 VPB.t4 248.598
R44 VPB.t3 VPB.t0 213.084
R45 VPB VPB.t3 189.408
R46 a_333_297.t0 a_333_297.t1 96.53
R47 A1.n0 A1.t1 236.179
R48 A1.n0 A1.t0 163.879
R49 A1 A1.n0 82.593
R50 a_461_297.t0 a_461_297.t1 53.19
R51 VPWR.n0 VPWR.t1 154.62
R52 VPWR.n0 VPWR.t0 144.755
R53 VPWR VPWR.n0 0.039
R54 B1.n0 B1.t0 230.361
R55 B1.n0 B1.t1 158.061
R56 B1 B1.n0 78.607
C0 VPWR Y 0.29fF
C1 A2 VPWR 0.11fF
C2 A3 A2 0.11fF
C3 B2 A3 0.15fF
C4 B2 Y 0.21fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__o32ai_2.ext - technology: sky130A

.subckt sky130_fd_sc_hd__o32ai_2 A1 B1 A2 A3 Y B2 VGND VPWR VNB VPB
X0 VGND.t3 A1.t0 a_27_47.t5 VNB.t5 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 a_27_47.t2 A3.t0 VGND.t0 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 a_475_297.t1 A2.t0 a_729_297.t3 VPB.t6 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 a_729_297.t1 A1.t1 VPWR.t3 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 VPWR.t2 A1.t2 a_729_297.t0 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 a_27_47.t8 A2.t1 VGND.t5 VNB.t8 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 a_27_297.t2 B1.t0 VPWR.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 a_729_297.t2 A2.t2 a_475_297.t0 VPB.t5 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 VPWR.t1 B1.t1 a_27_297.t1 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 VGND.t4 A2.t3 a_27_47.t7 VNB.t7 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 a_27_297.t3 B2.t0 Y.t1 VPB.t9 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 a_27_47.t9 B2.t1 Y.t3 VNB.t9 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 a_27_47.t0 B1.t2 Y.t5 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 a_475_297.t3 A3.t1 Y.t7 VPB.t8 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14 Y.t6 A3.t2 a_475_297.t2 VPB.t7 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 Y.t4 B1.t3 a_27_47.t1 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X16 a_27_47.t4 A1.t3 VGND.t2 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X17 VGND.t1 A3.t3 a_27_47.t3 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X18 Y.t0 B2.t2 a_27_297.t0 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X19 Y.t2 B2.t3 a_27_47.t6 VNB.t6 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
R0 A1.n0 A1.t2 223.763
R1 A1.n1 A1.t1 212.079
R2 A1.n1 A1.t0 151.463
R3 A1.n0 A1.t3 139.779
R4 A1.n3 A1.n2 76
R5 A1.n2 A1.n0 29.212
R6 A1.n2 A1.n1 20.448
R7 A1 A1.n3 17.408
R8 A1.n3 A1 6.144
R9 a_27_47.n1 a_27_47.t4 144.156
R10 a_27_47.n7 a_27_47.t6 134.603
R11 a_27_47.n8 a_27_47.n5 93.369
R12 a_27_47.n7 a_27_47.n6 92.5
R13 a_27_47.n9 a_27_47.n8 92.5
R14 a_27_47.n5 a_27_47.n4 52.212
R15 a_27_47.n8 a_27_47.n7 46.747
R16 a_27_47.n3 a_27_47.n2 46.25
R17 a_27_47.n1 a_27_47.n0 46.25
R18 a_27_47.n0 a_27_47.t5 43.384
R19 a_27_47.n5 a_27_47.n3 42.996
R20 a_27_47.n2 a_27_47.t8 39.692
R21 a_27_47.n6 a_27_47.t1 24.923
R22 a_27_47.n6 a_27_47.t9 24.923
R23 a_27_47.n4 a_27_47.t7 24.923
R24 a_27_47.n4 a_27_47.t2 24.923
R25 a_27_47.n9 a_27_47.t3 24.923
R26 a_27_47.t0 a_27_47.n9 24.923
R27 a_27_47.n3 a_27_47.n1 6.695
R28 VGND.n1 VGND.n0 114.711
R29 VGND.n3 VGND.n2 111.959
R30 VGND.n7 VGND.n6 107.239
R31 VGND.n6 VGND.t1 103.384
R32 VGND.n6 VGND.t0 42.461
R33 VGND.n2 VGND.t2 24.923
R34 VGND.n2 VGND.t3 24.923
R35 VGND.n0 VGND.t5 24.923
R36 VGND.n0 VGND.t4 24.923
R37 VGND.n3 VGND.n1 18.421
R38 VGND.n5 VGND.n4 4.65
R39 VGND.n9 VGND.n8 4.65
R40 VGND.n8 VGND.n7 3.011
R41 VGND VGND.n10 0.605
R42 VGND.n5 VGND.n3 0.158
R43 VGND.n10 VGND.n9 0.134
R44 VGND.n9 VGND.n5 0.119
R45 VNB VNB.t6 6078.09
R46 VNB.t8 VNB.t5 4545.05
R47 VNB.t3 VNB.t2 4545.05
R48 VNB.t5 VNB.t4 2030.77
R49 VNB.t7 VNB.t8 2030.77
R50 VNB.t2 VNB.t7 2030.77
R51 VNB.t0 VNB.t3 2030.77
R52 VNB.t1 VNB.t0 2030.77
R53 VNB.t9 VNB.t1 2030.77
R54 VNB.t6 VNB.t9 2030.77
R55 A3.n1 A3.t3 351.566
R56 A3.n0 A3.t1 220.842
R57 A3.n1 A3.t2 212.079
R58 A3.n0 A3.t0 139.779
R59 A3 A3.n2 99.04
R60 A3.n2 A3.n0 27.751
R61 A3.n2 A3.n1 24.83
R62 A2.n0 A2.t0 220.842
R63 A2.n1 A2.t2 212.079
R64 A2.n1 A2.t3 148.542
R65 A2.n0 A2.t1 139.779
R66 A2.n3 A2.n2 76
R67 A2.n3 A2 28.16
R68 A2.n2 A2.n0 27.751
R69 A2.n2 A2.n1 24.83
R70 A2 A2.n3 18.944
R71 a_729_297.n1 a_729_297.n0 339.271
R72 a_729_297.n0 a_729_297.t3 26.595
R73 a_729_297.n0 a_729_297.t2 26.595
R74 a_729_297.t0 a_729_297.n1 26.595
R75 a_729_297.n1 a_729_297.t1 26.595
R76 a_475_297.n1 a_475_297.t2 233.734
R77 a_475_297.t1 a_475_297.n1 233.733
R78 a_475_297.n1 a_475_297.n0 108.146
R79 a_475_297.n0 a_475_297.t0 26.595
R80 a_475_297.n0 a_475_297.t3 26.595
R81 VPB.t0 VPB.t7 591.9
R82 VPB.t6 VPB.t3 568.224
R83 VPB.t3 VPB.t2 248.598
R84 VPB.t5 VPB.t6 248.598
R85 VPB.t8 VPB.t5 248.598
R86 VPB.t7 VPB.t8 248.598
R87 VPB.t1 VPB.t0 248.598
R88 VPB.t9 VPB.t1 248.598
R89 VPB.t4 VPB.t9 248.598
R90 VPB VPB.t4 192.367
R91 VPWR.n15 VPWR.n14 314.711
R92 VPWR.n0 VPWR.t3 201.693
R93 VPWR.n1 VPWR.t2 165.825
R94 VPWR.n14 VPWR.t0 26.595
R95 VPWR.n14 VPWR.t1 26.595
R96 VPWR.n16 VPWR.n15 6.776
R97 VPWR.n17 VPWR.n16 4.65
R98 VPWR.n3 VPWR.n2 4.65
R99 VPWR.n5 VPWR.n4 4.65
R100 VPWR.n7 VPWR.n6 4.65
R101 VPWR.n9 VPWR.n8 4.65
R102 VPWR.n11 VPWR.n10 4.65
R103 VPWR.n13 VPWR.n12 4.65
R104 VPWR.n1 VPWR.n0 4.379
R105 VPWR.n3 VPWR.n1 0.267
R106 VPWR VPWR.n18 0.247
R107 VPWR.n18 VPWR.n17 0.134
R108 VPWR.n5 VPWR.n3 0.119
R109 VPWR.n7 VPWR.n5 0.119
R110 VPWR.n9 VPWR.n7 0.119
R111 VPWR.n11 VPWR.n9 0.119
R112 VPWR.n13 VPWR.n11 0.119
R113 VPWR.n17 VPWR.n13 0.119
R114 B1.n0 B1.t0 212.079
R115 B1.n1 B1.t1 212.079
R116 B1.n0 B1.t2 139.779
R117 B1.n1 B1.t3 139.779
R118 B1.n3 B1.n2 76
R119 B1.n2 B1.n0 30.672
R120 B1.n2 B1.n1 30.672
R121 B1.n3 B1 23.04
R122 B1 B1.n3 0.512
R123 a_27_297.t2 a_27_297.n1 230.121
R124 a_27_297.n1 a_27_297.t0 196.043
R125 a_27_297.n1 a_27_297.n0 142.024
R126 a_27_297.n0 a_27_297.t1 26.595
R127 a_27_297.n0 a_27_297.t3 26.595
R128 B2.n0 B2.t0 212.079
R129 B2.n1 B2.t2 212.079
R130 B2.n0 B2.t1 139.779
R131 B2.n1 B2.t3 139.779
R132 B2 B2.n2 79.584
R133 B2.n2 B2.n0 30.672
R134 B2.n2 B2.n1 30.672
R135 Y.n5 Y.n3 230.13
R136 Y.n5 Y.n4 198.13
R137 Y.n2 Y.n1 135.508
R138 Y.n2 Y.n0 92.5
R139 Y Y.n2 37.586
R140 Y.n4 Y.t7 26.595
R141 Y.n4 Y.t6 26.595
R142 Y.n3 Y.t1 26.595
R143 Y.n3 Y.t0 26.595
R144 Y.n0 Y.t5 24.923
R145 Y.n0 Y.t4 24.923
R146 Y.n1 Y.t3 24.923
R147 Y.n1 Y.t2 24.923
R148 Y Y.n5 5.857
C0 A3 Y 0.20fF
C1 VPB VPWR 0.12fF
C2 B2 Y 0.13fF
C3 B1 Y 0.34fF
C4 VPWR VGND 0.12fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__o32ai_4.ext - technology: sky130A

.subckt sky130_fd_sc_hd__o32ai_4 A1 A2 A3 B1 Y B2 VGND VPWR VNB VPB
X0 a_1224_297.t7 A1.t0 VPWR.t6 VPB.t12 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 VPWR.t5 A1.t1 a_1224_297.t6 VPB.t11 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 a_27_297.t3 B1.t0 VPWR.t1 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 a_27_47.t15 A1.t2 VGND.t7 VNB.t15 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 a_27_297.t6 B2.t0 Y.t11 VPB.t18 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 VPWR.t0 B1.t1 a_27_297.t2 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 a_806_297.t4 A3.t0 Y.t12 VPB.t13 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 VGND.t0 A2.t0 a_27_47.t0 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 VGND.t1 A2.t1 a_27_47.t9 VNB.t9 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 a_27_47.t16 A3.t1 VGND.t8 VNB.t16 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 Y.t10 B2.t1 a_27_297.t7 VPB.t19 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 a_806_297.t3 A3.t2 Y.t13 VPB.t14 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 Y.t14 A3.t3 a_806_297.t2 VPB.t15 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13 a_27_47.t4 B1.t2 Y.t3 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14 a_27_297.t4 B2.t2 Y.t9 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 a_27_47.t5 B2.t3 Y.t7 VNB.t5 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X16 a_27_47.t6 B2.t4 Y.t6 VNB.t6 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X17 a_27_47.t3 B1.t3 Y.t2 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X18 Y.t15 A3.t4 a_806_297.t1 VPB.t16 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X19 a_27_47.t10 A2.t2 VGND.t2 VNB.t10 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X20 a_27_47.t11 A2.t3 VGND.t3 VNB.t11 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X21 a_27_47.t14 A1.t3 VGND.t6 VNB.t14 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X22 a_27_297.t1 B1.t4 VPWR.t2 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X23 Y.t1 B1.t5 a_27_47.t2 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X24 a_806_297.t5 A2.t4 a_1224_297.t1 VPB.t6 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X25 Y.t5 B2.t5 a_27_47.t7 VNB.t7 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X26 Y.t0 B1.t6 a_27_47.t1 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X27 VPWR.t7 B1.t7 a_27_297.t0 VPB.t17 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X28 VGND.t9 A3.t5 a_27_47.t17 VNB.t17 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X29 VGND.t10 A3.t6 a_27_47.t18 VNB.t18 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X30 a_1224_297.t2 A2.t5 a_806_297.t6 VPB.t7 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X31 a_1224_297.t5 A1.t4 VPWR.t4 VPB.t10 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X32 a_806_297.t7 A2.t6 a_1224_297.t3 VPB.t8 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X33 VPWR.t3 A1.t5 a_1224_297.t4 VPB.t9 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X34 Y.t8 B2.t6 a_27_297.t5 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X35 a_27_47.t19 A3.t7 VGND.t11 VNB.t19 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X36 VGND.t5 A1.t6 a_27_47.t13 VNB.t13 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X37 a_1224_297.t0 A2.t7 a_806_297.t0 VPB.t5 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X38 Y.t4 B2.t7 a_27_47.t8 VNB.t8 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X39 VGND.t4 A1.t7 a_27_47.t12 VNB.t12 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
R0 A1.n0 A1.t1 218.506
R1 A1.n7 A1.t4 218.506
R2 A1.n3 A1.t5 218.506
R3 A1.n1 A1.t0 218.506
R4 A1.n0 A1.t3 146.206
R5 A1.n7 A1.t7 146.206
R6 A1.n3 A1.t2 146.206
R7 A1.n1 A1.t6 146.206
R8 A1.n10 A1.n0 95.113
R9 A1.n9 A1.n8 76
R10 A1.n6 A1.n5 76
R11 A1.n8 A1.n0 50.693
R12 A1.n8 A1.n7 34.903
R13 A1.n7 A1.n6 34.903
R14 A1.n6 A1.n3 34.903
R15 A1.n3 A1.n2 34.903
R16 A1.n2 A1.n1 34.903
R17 A1.n5 A1.n4 26.88
R18 A1.n9 A1 24.64
R19 A1.n10 A1 22.08
R20 A1 A1.n10 7.36
R21 A1 A1.n9 4.8
R22 A1.n5 A1 2.24
R23 A1.n4 A1 0.32
R24 VPWR.n28 VPWR.n27 307.239
R25 VPWR.n32 VPWR.n31 307.239
R26 VPWR.n5 VPWR.t6 196.528
R27 VPWR.n1 VPWR.n0 174.594
R28 VPWR.n2 VPWR.t5 145.704
R29 VPWR.n0 VPWR.t4 26.595
R30 VPWR.n0 VPWR.t3 26.595
R31 VPWR.n27 VPWR.t1 26.595
R32 VPWR.n27 VPWR.t0 26.595
R33 VPWR.n31 VPWR.t2 26.595
R34 VPWR.n31 VPWR.t7 26.595
R35 VPWR.n2 VPWR.n1 11.191
R36 VPWR.n4 VPWR.n3 4.65
R37 VPWR.n6 VPWR.n5 4.65
R38 VPWR.n8 VPWR.n7 4.65
R39 VPWR.n10 VPWR.n9 4.65
R40 VPWR.n12 VPWR.n11 4.65
R41 VPWR.n14 VPWR.n13 4.65
R42 VPWR.n16 VPWR.n15 4.65
R43 VPWR.n18 VPWR.n17 4.65
R44 VPWR.n20 VPWR.n19 4.65
R45 VPWR.n22 VPWR.n21 4.65
R46 VPWR.n24 VPWR.n23 4.65
R47 VPWR.n26 VPWR.n25 4.65
R48 VPWR.n30 VPWR.n29 4.65
R49 VPWR.n29 VPWR.n28 4.517
R50 VPWR.n33 VPWR.n32 3.508
R51 VPWR VPWR.n33 0.585
R52 VPWR.n4 VPWR.n2 0.23
R53 VPWR.n33 VPWR.n30 0.151
R54 VPWR.n6 VPWR.n4 0.119
R55 VPWR.n8 VPWR.n6 0.119
R56 VPWR.n10 VPWR.n8 0.119
R57 VPWR.n12 VPWR.n10 0.119
R58 VPWR.n14 VPWR.n12 0.119
R59 VPWR.n16 VPWR.n14 0.119
R60 VPWR.n18 VPWR.n16 0.119
R61 VPWR.n20 VPWR.n18 0.119
R62 VPWR.n22 VPWR.n20 0.119
R63 VPWR.n24 VPWR.n22 0.119
R64 VPWR.n26 VPWR.n24 0.119
R65 VPWR.n30 VPWR.n26 0.119
R66 a_1224_297.n2 a_1224_297.n0 190.978
R67 a_1224_297.n2 a_1224_297.n1 152.578
R68 a_1224_297.n5 a_1224_297.n4 146.035
R69 a_1224_297.n4 a_1224_297.n3 107.635
R70 a_1224_297.n4 a_1224_297.n2 77.552
R71 a_1224_297.t6 a_1224_297.n5 45.31
R72 a_1224_297.n0 a_1224_297.t3 26.595
R73 a_1224_297.n0 a_1224_297.t0 26.595
R74 a_1224_297.n1 a_1224_297.t1 26.595
R75 a_1224_297.n1 a_1224_297.t2 26.595
R76 a_1224_297.n3 a_1224_297.t4 26.595
R77 a_1224_297.n3 a_1224_297.t7 26.595
R78 a_1224_297.n5 a_1224_297.t5 26.595
R79 VPB.t6 VPB.t12 556.386
R80 VPB.t1 VPB.t16 556.386
R81 VPB.t10 VPB.t11 304.828
R82 VPB.t18 VPB.t17 257.476
R83 VPB.t9 VPB.t10 248.598
R84 VPB.t12 VPB.t9 248.598
R85 VPB.t7 VPB.t6 248.598
R86 VPB.t8 VPB.t7 248.598
R87 VPB.t5 VPB.t8 248.598
R88 VPB.t13 VPB.t5 248.598
R89 VPB.t15 VPB.t13 248.598
R90 VPB.t14 VPB.t15 248.598
R91 VPB.t16 VPB.t14 248.598
R92 VPB.t0 VPB.t1 248.598
R93 VPB.t2 VPB.t0 248.598
R94 VPB.t17 VPB.t2 248.598
R95 VPB.t19 VPB.t18 248.598
R96 VPB.t3 VPB.t19 248.598
R97 VPB.t4 VPB.t3 248.598
R98 VPB VPB.t4 189.408
R99 B1.n0 B1.t0 218.506
R100 B1.n2 B1.t1 218.506
R101 B1.n5 B1.t4 218.506
R102 B1.n3 B1.t7 218.506
R103 B1.n0 B1.t3 146.206
R104 B1.n2 B1.t6 146.206
R105 B1.n5 B1.t2 146.206
R106 B1.n3 B1.t5 146.206
R107 B1.n4 B1 81.12
R108 B1.n8 B1.n1 76
R109 B1.n7 B1.n6 76
R110 B1.n6 B1.n2 35.734
R111 B1.n5 B1.n4 35.734
R112 B1.n1 B1.n0 34.903
R113 B1.n2 B1.n1 34.903
R114 B1.n6 B1.n5 34.072
R115 B1.n4 B1.n3 34.072
R116 B1.n7 B1 21.76
R117 B1.n8 B1 19.52
R118 B1 B1.n8 9.92
R119 B1 B1.n7 7.68
R120 a_27_297.n4 a_27_297.n3 292.5
R121 a_27_297.t3 a_27_297.n5 233.918
R122 a_27_297.n2 a_27_297.t5 180.11
R123 a_27_297.n2 a_27_297.n1 150.897
R124 a_27_297.n5 a_27_297.n0 150.897
R125 a_27_297.n5 a_27_297.n4 75.67
R126 a_27_297.n4 a_27_297.n2 58.514
R127 a_27_297.n3 a_27_297.t6 29.55
R128 a_27_297.n0 a_27_297.t2 26.595
R129 a_27_297.n0 a_27_297.t1 26.595
R130 a_27_297.n3 a_27_297.t0 26.595
R131 a_27_297.n1 a_27_297.t7 26.595
R132 a_27_297.n1 a_27_297.t4 26.595
R133 VGND.n5 VGND.n2 114.795
R134 VGND.n4 VGND.n3 114.711
R135 VGND.n11 VGND.n10 114.711
R136 VGND.n17 VGND.n16 114.711
R137 VGND.n1 VGND.n0 114.711
R138 VGND.n25 VGND.n24 107.239
R139 VGND.n24 VGND.t8 39.692
R140 VGND.n24 VGND.t10 39.692
R141 VGND.n2 VGND.t6 34.153
R142 VGND.n2 VGND.t4 33.23
R143 VGND.n3 VGND.t7 24.923
R144 VGND.n3 VGND.t5 24.923
R145 VGND.n10 VGND.t3 24.923
R146 VGND.n10 VGND.t1 24.923
R147 VGND.n16 VGND.t2 24.923
R148 VGND.n16 VGND.t0 24.923
R149 VGND.n0 VGND.t11 24.923
R150 VGND.n0 VGND.t9 24.923
R151 VGND.n29 VGND.n1 15.057
R152 VGND.n5 VGND.n4 8.2
R153 VGND.n7 VGND.n6 4.65
R154 VGND.n9 VGND.n8 4.65
R155 VGND.n13 VGND.n12 4.65
R156 VGND.n15 VGND.n14 4.65
R157 VGND.n19 VGND.n18 4.65
R158 VGND.n21 VGND.n20 4.65
R159 VGND.n23 VGND.n22 4.65
R160 VGND.n26 VGND.n25 4.65
R161 VGND.n28 VGND.n27 4.65
R162 VGND.n18 VGND.n17 3.388
R163 VGND.n12 VGND.n11 2.635
R164 VGND VGND.n29 0.962
R165 VGND.n7 VGND.n5 0.211
R166 VGND.n29 VGND.n28 0.134
R167 VGND.n9 VGND.n7 0.119
R168 VGND.n13 VGND.n9 0.119
R169 VGND.n15 VGND.n13 0.119
R170 VGND.n19 VGND.n15 0.119
R171 VGND.n21 VGND.n19 0.119
R172 VGND.n23 VGND.n21 0.119
R173 VGND.n26 VGND.n23 0.119
R174 VGND.n28 VGND.n26 0.119
R175 a_27_47.n20 a_27_47.t14 138.824
R176 a_27_47.n5 a_27_47.t8 136.727
R177 a_27_47.n7 a_27_47.n2 92.5
R178 a_27_47.n6 a_27_47.n3 92.5
R179 a_27_47.n5 a_27_47.n4 92.5
R180 a_27_47.n9 a_27_47.n7 55.425
R181 a_27_47.n18 a_27_47.t13 54.461
R182 a_27_47.n12 a_27_47.n11 53.696
R183 a_27_47.n20 a_27_47.n19 53.696
R184 a_27_47.n11 a_27_47.n10 52.6
R185 a_27_47.n16 a_27_47.n15 52.6
R186 a_27_47.n21 a_27_47.n20 52.599
R187 a_27_47.n7 a_27_47.n6 52.114
R188 a_27_47.n6 a_27_47.n5 51.2
R189 a_27_47.n11 a_27_47.n9 50.878
R190 a_27_47.n12 a_27_47.n1 46.25
R191 a_27_47.n14 a_27_47.n13 46.25
R192 a_27_47.n17 a_27_47.n0 46.25
R193 a_27_47.n19 a_27_47.n18 46.25
R194 a_27_47.n16 a_27_47.n14 43.154
R195 a_27_47.n9 a_27_47.n8 42.06
R196 a_27_47.n17 a_27_47.n16 41.649
R197 a_27_47.n13 a_27_47.t0 28.615
R198 a_27_47.n3 a_27_47.t2 27.692
R199 a_27_47.n0 a_27_47.t11 24.923
R200 a_27_47.n1 a_27_47.t16 24.923
R201 a_27_47.n8 a_27_47.t17 24.923
R202 a_27_47.n8 a_27_47.t3 24.923
R203 a_27_47.n4 a_27_47.t7 24.923
R204 a_27_47.n4 a_27_47.t5 24.923
R205 a_27_47.n3 a_27_47.t6 24.923
R206 a_27_47.n2 a_27_47.t1 24.923
R207 a_27_47.n2 a_27_47.t4 24.923
R208 a_27_47.n10 a_27_47.t18 24.923
R209 a_27_47.n10 a_27_47.t19 24.923
R210 a_27_47.n15 a_27_47.t9 24.923
R211 a_27_47.n15 a_27_47.t10 24.923
R212 a_27_47.n21 a_27_47.t12 24.923
R213 a_27_47.t15 a_27_47.n21 24.923
R214 a_27_47.n19 a_27_47.n17 7.089
R215 a_27_47.n14 a_27_47.n12 6.695
R216 VNB VNB.t8 6053.91
R217 VNB.t11 VNB.t13 4545.05
R218 VNB.t16 VNB.t0 3771.43
R219 VNB.t18 VNB.t16 2804.4
R220 VNB.t12 VNB.t14 2490.11
R221 VNB.t6 VNB.t2 2103.3
R222 VNB.t15 VNB.t12 2030.77
R223 VNB.t13 VNB.t15 2030.77
R224 VNB.t9 VNB.t11 2030.77
R225 VNB.t10 VNB.t9 2030.77
R226 VNB.t0 VNB.t10 2030.77
R227 VNB.t19 VNB.t18 2030.77
R228 VNB.t17 VNB.t19 2030.77
R229 VNB.t3 VNB.t17 2030.77
R230 VNB.t1 VNB.t3 2030.77
R231 VNB.t4 VNB.t1 2030.77
R232 VNB.t2 VNB.t4 2030.77
R233 VNB.t7 VNB.t6 2030.77
R234 VNB.t5 VNB.t7 2030.77
R235 VNB.t8 VNB.t5 2030.77
R236 B2.n1 B2.t0 218.506
R237 B2.n3 B2.t1 218.506
R238 B2.n0 B2.t2 218.506
R239 B2.n8 B2.t6 218.506
R240 B2.n1 B2.t4 146.206
R241 B2.n3 B2.t5 146.206
R242 B2.n0 B2.t3 146.206
R243 B2.n8 B2.t7 146.206
R244 B2.n9 B2.n8 108.41
R245 B2.n5 B2.n4 76
R246 B2.n7 B2.n6 76
R247 B2.n2 B2.n1 34.903
R248 B2.n3 B2.n2 34.903
R249 B2.n4 B2.n3 34.903
R250 B2.n4 B2.n0 34.903
R251 B2.n7 B2.n0 34.903
R252 B2.n8 B2.n7 34.903
R253 B2.n6 B2 24.96
R254 B2.n9 B2 21.44
R255 B2 B2.n9 8
R256 B2.n6 B2 4.48
R257 B2 B2.n5 1.92
R258 Y.n3 Y.n1 190.978
R259 Y.n12 Y.n0 190.978
R260 Y.n11 Y.n3 178.823
R261 Y.n3 Y.n2 152.578
R262 Y.n14 Y.n13 147.068
R263 Y.n9 Y.n8 135.508
R264 Y.n6 Y.n4 135.508
R265 Y.n9 Y.n7 92.5
R266 Y.n6 Y.n5 92.5
R267 Y.n11 Y.n10 48
R268 Y.n13 Y.t11 26.595
R269 Y.n13 Y.t10 26.595
R270 Y.n1 Y.t12 26.595
R271 Y.n1 Y.t14 26.595
R272 Y.n2 Y.t13 26.595
R273 Y.n2 Y.t15 26.595
R274 Y.n0 Y.t9 26.595
R275 Y.n0 Y.t8 26.595
R276 Y.n4 Y.t2 24.923
R277 Y.n4 Y.t0 24.923
R278 Y.n5 Y.t3 24.923
R279 Y.n5 Y.t1 24.923
R280 Y.n7 Y.t6 24.923
R281 Y.n7 Y.t5 24.923
R282 Y.n8 Y.t7 24.923
R283 Y.n8 Y.t4 24.923
R284 Y.n10 Y.n6 22.016
R285 Y.n10 Y.n9 21.76
R286 Y.n12 Y.n11 11.67
R287 Y.n14 Y.n12 5.238
R288 Y Y.n14 2.332
R289 A3.n2 A3.t0 278.34
R290 A3.n3 A3.t3 218.506
R291 A3.n5 A3.t2 218.506
R292 A3.n0 A3.t4 218.506
R293 A3.n12 A3.t5 161.164
R294 A3.n11 A3.t7 146.206
R295 A3.n6 A3.t6 146.206
R296 A3.n2 A3.t1 146.206
R297 A3.n8 A3.n7 76
R298 A3.n10 A3.n9 76
R299 A3.n13 A3.n12 76
R300 A3.n5 A3.n4 68.144
R301 A3.n12 A3.n11 54.848
R302 A3.n6 A3.n0 53.186
R303 A3.n8 A3.n1 26.88
R304 A3.n9 A3 25.28
R305 A3.n13 A3 22.72
R306 A3.n7 A3.n6 14.958
R307 A3.n11 A3.n10 14.958
R308 A3.n3 A3.n2 9.972
R309 A3 A3.n13 6.72
R310 A3.n9 A3 4.16
R311 A3.n4 A3.n3 1.662
R312 A3.n7 A3.n5 1.662
R313 A3.n10 A3.n0 1.662
R314 A3 A3.n8 1.6
R315 A3.n1 A3 0.96
R316 a_806_297.n3 a_806_297.t1 224.115
R317 a_806_297.n1 a_806_297.t5 224.115
R318 a_806_297.n5 a_806_297.n4 150.898
R319 a_806_297.n1 a_806_297.n0 150.897
R320 a_806_297.n3 a_806_297.n2 150.897
R321 a_806_297.n4 a_806_297.n1 51.2
R322 a_806_297.n4 a_806_297.n3 51.2
R323 a_806_297.n2 a_806_297.t2 26.595
R324 a_806_297.n2 a_806_297.t3 26.595
R325 a_806_297.n0 a_806_297.t6 26.595
R326 a_806_297.n0 a_806_297.t7 26.595
R327 a_806_297.n5 a_806_297.t0 26.595
R328 a_806_297.t4 a_806_297.n5 26.595
R329 A2.n1 A2.t4 218.506
R330 A2.n0 A2.t5 218.506
R331 A2.n5 A2.t6 218.506
R332 A2.n6 A2.t7 218.506
R333 A2.n1 A2.t3 146.206
R334 A2.n0 A2.t1 146.206
R335 A2.n5 A2.t2 146.206
R336 A2.n6 A2.t0 146.206
R337 A2 A2.n2 78.88
R338 A2.n4 A2.n3 76
R339 A2.n8 A2.n7 76
R340 A2.n2 A2.n1 34.903
R341 A2.n2 A2.n0 34.903
R342 A2.n4 A2.n0 34.903
R343 A2.n5 A2.n4 34.903
R344 A2.n7 A2.n5 34.903
R345 A2.n7 A2.n6 34.903
R346 A2.n3 A2 24
R347 A2.n8 A2 21.44
R348 A2 A2.n8 8
R349 A2.n3 A2 5.44
C0 VPWR VGND 0.21fF
C1 A3 Y 0.33fF
C2 B2 Y 0.42fF
C3 VPB VPWR 0.20fF
C4 B1 Y 0.52fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__o41a_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__o41a_1 A1 A2 A3 A4 B1 X VGND VPWR VNB VPB
X0 VGND.t0 A4.t0 a_321_47.t0 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 a_321_47.t4 A3.t0 VGND.t4 VNB.t5 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 a_103_21.t2 B1.t0 VPWR.t2 VPB.t5 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 VPWR.t1 a_103_21.t3 X.t1 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 VGND.t3 a_103_21.t4 X.t0 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 VGND.t2 A2.t0 a_321_47.t3 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 a_321_47.t2 A1.t0 VGND.t1 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 a_511_297.t0 A3.t1 a_393_297.t1 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 a_619_297.t1 A2.t1 a_511_297.t1 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 a_321_47.t1 B1.t1 a_103_21.t1 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 a_393_297.t0 A4.t1 a_103_21.t0 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 VPWR.t0 A1.t1 a_619_297.t0 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
R0 A4.n0 A4.t1 233.007
R1 A4.n0 A4.t0 162.917
R2 A4 A4.n0 87.054
R3 a_321_47.n2 a_321_47.n1 167.417
R4 a_321_47.n1 a_321_47.t2 140.466
R5 a_321_47.n1 a_321_47.n0 52.431
R6 a_321_47.n0 a_321_47.t3 36.923
R7 a_321_47.n0 a_321_47.t4 35.076
R8 a_321_47.t0 a_321_47.n2 24.923
R9 a_321_47.n2 a_321_47.t1 24.923
R10 VGND.n8 VGND.t3 197.787
R11 VGND.n3 VGND.n0 110.707
R12 VGND.n2 VGND.n1 107.239
R13 VGND.n0 VGND.t1 36
R14 VGND.n0 VGND.t2 36
R15 VGND.n1 VGND.t4 35.076
R16 VGND.n1 VGND.t0 35.076
R17 VGND.n9 VGND.n8 12.429
R18 VGND.n5 VGND.n4 4.65
R19 VGND.n7 VGND.n6 4.65
R20 VGND.n3 VGND.n2 3.524
R21 VGND.n5 VGND.n3 0.176
R22 VGND.n9 VGND.n7 0.132
R23 VGND VGND.n9 0.129
R24 VGND.n7 VGND.n5 0.119
R25 VNB VNB.t4 6658.31
R26 VNB.t4 VNB.t1 4545.05
R27 VNB.t3 VNB.t2 2610.99
R28 VNB.t5 VNB.t3 2610.99
R29 VNB.t0 VNB.t5 2562.64
R30 VNB.t1 VNB.t0 2030.77
R31 A3.n0 A3.t1 236.179
R32 A3.n0 A3.t0 163.879
R33 A3 A3.n0 87.054
R34 B1.n0 B1.t0 262.574
R35 B1.n0 B1.t1 157.306
R36 B1 B1.n0 81.18
R37 VPWR.n1 VPWR.n0 167.457
R38 VPWR.n1 VPWR.t0 150.143
R39 VPWR.n0 VPWR.t2 26.595
R40 VPWR.n0 VPWR.t1 26.595
R41 VPWR VPWR.n1 0.245
R42 a_103_21.n0 a_103_21.t3 234.17
R43 a_103_21.n0 a_103_21.t4 162.697
R44 a_103_21.n2 a_103_21.n1 138.117
R45 a_103_21.n1 a_103_21.t1 108.082
R46 a_103_21.n1 a_103_21.n0 78.742
R47 a_103_21.t0 a_103_21.n2 60.085
R48 a_103_21.n2 a_103_21.t2 42.355
R49 VPB.t5 VPB.t2 396.573
R50 VPB VPB.t0 387.694
R51 VPB.t2 VPB.t3 349.221
R52 VPB.t4 VPB.t1 319.626
R53 VPB.t3 VPB.t4 319.626
R54 VPB.t0 VPB.t5 248.598
R55 X.n2 X.n1 292.5
R56 X.n1 X.n0 146.431
R57 X X.n5 94.194
R58 X.n6 X.n5 92.5
R59 X.n1 X.t1 55.16
R60 X.n5 X.t0 47.076
R61 X.n6 X 11.105
R62 X.n4 X 10.429
R63 X.n0 X 6.374
R64 X.n4 X 5.688
R65 X X.n4 4.517
R66 X.n3 X.n2 4.266
R67 X.n2 X 3.779
R68 X.n0 X 1.892
R69 X X.n6 1.694
R70 X X.n3 0.474
R71 X.n3 X 0.243
R72 A2.n0 A2.t1 236.179
R73 A2.n0 A2.t0 163.879
R74 A2 A2.n0 85.859
R75 A1.n0 A1.t1 236.179
R76 A1.n0 A1.t0 163.879
R77 A1 A1.n0 84.96
R78 a_393_297.t0 a_393_297.t1 86.68
R79 a_511_297.t0 a_511_297.t1 76.83
R80 a_619_297.t0 a_619_297.t1 76.83
C0 X VPWR 0.15fF
C1 A2 A3 0.27fF
C2 A2 VPWR 0.12fF
C3 A4 A3 0.22fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__o41a_2.ext - technology: sky130A

.subckt sky130_fd_sc_hd__o41a_2 A1 A2 A3 A4 B1 X VGND VPWR VNB VPB
X0 VGND.t1 A2.t0 a_393_47.t2 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 a_496_297.t0 A4.t0 a_79_21.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 a_393_47.t3 A3.t0 VGND.t2 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 VPWR.t3 A1.t0 a_697_297.t1 VPB.t6 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 VPWR.t2 a_79_21.t3 X.t3 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 VGND.t3 a_79_21.t4 X.t1 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 a_79_21.t1 B1.t0 VPWR.t0 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 VGND.t0 A4.t1 a_393_47.t0 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 a_697_297.t0 A2.t1 a_597_297.t1 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 a_393_47.t4 A1.t1 VGND.t5 VNB.t6 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 X.t2 a_79_21.t5 VPWR.t1 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 a_393_47.t1 B1.t1 a_79_21.t2 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 a_597_297.t0 A3.t1 a_496_297.t1 VPB.t5 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13 X.t0 a_79_21.t6 VGND.t4 VNB.t5 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
R0 A2.n0 A2.t1 239.503
R1 A2.n0 A2.t0 167.203
R2 A2.n1 A2.n0 76
R3 A2.n1 A2 11.054
R4 A2 A2.n1 2.133
R5 a_393_47.n1 a_393_47.t4 150.595
R6 a_393_47.n2 a_393_47.n1 95.932
R7 a_393_47.n1 a_393_47.n0 52.818
R8 a_393_47.n0 a_393_47.t2 39.692
R9 a_393_47.n2 a_393_47.t1 34.153
R10 a_393_47.t0 a_393_47.n2 33.23
R11 a_393_47.n0 a_393_47.t3 24.923
R12 VGND.n3 VGND.n2 115.927
R13 VGND.n1 VGND.n0 110.854
R14 VGND.n8 VGND.t3 109.725
R15 VGND.n12 VGND.t4 108.334
R16 VGND.n0 VGND.t2 40.615
R17 VGND.n2 VGND.t5 36
R18 VGND.n2 VGND.t1 28.615
R19 VGND.n0 VGND.t0 24.923
R20 VGND.n13 VGND.n12 4.65
R21 VGND.n5 VGND.n4 4.65
R22 VGND.n7 VGND.n6 4.65
R23 VGND.n9 VGND.n8 4.65
R24 VGND.n11 VGND.n10 4.65
R25 VGND.n3 VGND.n1 3.773
R26 VGND.n5 VGND.n3 0.196
R27 VGND.n7 VGND.n5 0.119
R28 VGND.n9 VGND.n7 0.119
R29 VGND.n11 VGND.n9 0.119
R30 VGND.n13 VGND.n11 0.119
R31 VGND VGND.n13 0.02
R32 VNB VNB.t5 6053.91
R33 VNB.t4 VNB.t1 4835.16
R34 VNB.t1 VNB.t0 2490.11
R35 VNB.t0 VNB.t3 2441.76
R36 VNB.t2 VNB.t6 2417.58
R37 VNB.t3 VNB.t2 2417.58
R38 VNB.t5 VNB.t4 2030.77
R39 A4.n0 A4.t0 239.038
R40 A4.n0 A4.t1 166.738
R41 A4.n1 A4.n0 76
R42 A4.n1 A4 11.054
R43 A4 A4.n1 2.133
R44 a_79_21.n1 a_79_21.t3 205.652
R45 a_79_21.n0 a_79_21.t5 205.652
R46 a_79_21.n1 a_79_21.t4 133.353
R47 a_79_21.n0 a_79_21.t6 133.353
R48 a_79_21.n2 a_79_21.n1 132.889
R49 a_79_21.n3 a_79_21.n2 125.464
R50 a_79_21.n2 a_79_21.t2 108.801
R51 a_79_21.t0 a_79_21.n3 92.59
R52 a_79_21.n1 a_79_21.n0 54.713
R53 a_79_21.n3 a_79_21.t1 26.595
R54 a_496_297.t0 a_496_297.t1 69.935
R55 VPB.t4 VPB.t1 449.844
R56 VPB.t1 VPB.t0 446.884
R57 VPB.t0 VPB.t5 298.909
R58 VPB.t2 VPB.t6 295.95
R59 VPB.t5 VPB.t2 295.95
R60 VPB.t3 VPB.t4 248.598
R61 VPB VPB.t3 189.408
R62 A3.n0 A3.t1 239.503
R63 A3.n0 A3.t0 167.203
R64 A3.n1 A3.n0 76
R65 A3.n1 A3 11.054
R66 A3 A3.n1 2.133
R67 A1.n0 A1.t0 239.503
R68 A1.n0 A1.t1 167.203
R69 A1 A1.n0 91.104
R70 a_697_297.t0 a_697_297.t1 68.95
R71 VPWR.n2 VPWR.t3 171.872
R72 VPWR.n5 VPWR.t1 151.631
R73 VPWR.n0 VPWR.t0 60.085
R74 VPWR.n0 VPWR.t2 56.858
R75 VPWR.n1 VPWR.n0 13.803
R76 VPWR.n4 VPWR.n3 4.65
R77 VPWR.n6 VPWR.n5 4.65
R78 VPWR.n2 VPWR.n1 3.199
R79 VPWR.n4 VPWR.n2 0.16
R80 VPWR.n6 VPWR.n4 0.119
R81 VPWR VPWR.n6 0.02
R82 X.n5 X.n4 292.5
R83 X.n6 X.n5 147.104
R84 X X.n0 94.245
R85 X.n1 X.n0 92.5
R86 X.n5 X.t3 26.595
R87 X.n5 X.t2 26.595
R88 X.n0 X.t1 24.923
R89 X.n0 X.t0 24.923
R90 X.n1 X 11.442
R91 X.n6 X 10.71
R92 X X.n2 10.472
R93 X.n4 X.n3 6.4
R94 X.n2 X 5.352
R95 X.n4 X 4.848
R96 X.n2 X 4.46
R97 X X.n6 2.439
R98 X.n3 X 2.327
R99 X.n3 X 1.939
R100 X X.n1 1.745
R101 B1.n0 B1.t0 264.563
R102 B1.n0 B1.t1 149.419
R103 B1 B1.n0 86.777
R104 a_597_297.t0 a_597_297.t1 68.95
C0 VPWR VGND 0.12fF
C1 A4 A3 0.26fF
C2 X VGND 0.27fF
C3 VPB VPWR 0.10fF
C4 VPWR X 0.35fF
C5 A3 A2 0.26fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__o41a_4.ext - technology: sky130A

.subckt sky130_fd_sc_hd__o41a_4 A1 A2 A3 A4 B1 X VGND VPWR VNB VPB
X0 a_467_47.t9 A4.t0 VGND.t7 VNB.t9 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 a_467_47.t4 A3.t0 VGND.t4 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 VGND.t2 A1.t0 a_467_47.t2 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 a_467_47.t6 B1.t0 a_79_21.t5 VNB.t6 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 a_467_47.t1 A2.t0 VGND.t1 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 a_79_21.t3 B1.t1 VPWR.t7 VPB.t13 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 VPWR.t1 A1.t1 a_1083_297.t3 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 VPWR.t5 a_79_21.t6 X.t7 VPB.t7 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 a_1083_297.t0 A2.t1 a_889_297.t1 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 VGND.t5 A3.t1 a_467_47.t5 VNB.t5 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 a_79_21.t4 B1.t2 a_467_47.t7 VNB.t7 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 X.t6 a_79_21.t7 VPWR.t4 VPB.t6 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 a_889_297.t0 A2.t2 a_1083_297.t1 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13 VPWR.t3 a_79_21.t8 X.t5 VPB.t5 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14 VGND.t8 a_79_21.t9 X.t3 VNB.t10 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X15 VGND.t9 a_79_21.t10 X.t2 VNB.t11 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X16 a_639_297.t3 A3.t2 a_889_297.t3 VPB.t11 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17 VGND.t0 A2.t3 a_467_47.t0 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X18 a_889_297.t2 A3.t3 a_639_297.t2 VPB.t10 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X19 X.t1 a_79_21.t11 VGND.t10 VNB.t12 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X20 a_639_297.t1 A4.t1 a_79_21.t1 VPB.t9 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X21 VPWR.t6 B1.t3 a_79_21.t2 VPB.t12 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X22 VGND.t6 A4.t2 a_467_47.t8 VNB.t8 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X23 a_1083_297.t2 A1.t2 VPWR.t0 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X24 a_79_21.t0 A4.t3 a_639_297.t0 VPB.t8 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X25 a_467_47.t3 A1.t3 VGND.t3 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X26 X.t4 a_79_21.t12 VPWR.t2 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X27 X.t0 a_79_21.t13 VGND.t11 VNB.t13 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
R0 A4.n0 A4.t1 221.719
R1 A4.n1 A4.t3 221.719
R2 A4.n0 A4.t0 149.419
R3 A4.n1 A4.t2 149.419
R4 A4.n3 A4.n2 76
R5 A4.n2 A4.n0 37.488
R6 A4.n2 A4.n1 37.488
R7 A4 A4.n3 21.12
R8 A4.n3 A4 8.32
R9 VGND.n36 VGND.t11 194.283
R10 VGND.n31 VGND.n30 114.711
R11 VGND.n17 VGND.n16 114.609
R12 VGND.n1 VGND.n0 114.285
R13 VGND.n13 VGND.n12 110.514
R14 VGND.n26 VGND.t9 109.244
R15 VGND.n3 VGND.n2 92.5
R16 VGND.n7 VGND.n6 92.5
R17 VGND.n2 VGND.t1 24.923
R18 VGND.n6 VGND.t0 24.923
R19 VGND.n0 VGND.t3 24.923
R20 VGND.n0 VGND.t2 24.923
R21 VGND.n12 VGND.t4 24.923
R22 VGND.n12 VGND.t5 24.923
R23 VGND.n16 VGND.t7 24.923
R24 VGND.n16 VGND.t6 24.923
R25 VGND.n30 VGND.t10 24.923
R26 VGND.n30 VGND.t8 24.923
R27 VGND.n14 VGND.n13 5.647
R28 VGND.n37 VGND.n36 4.65
R29 VGND.n5 VGND.n4 4.65
R30 VGND.n9 VGND.n8 4.65
R31 VGND.n11 VGND.n10 4.65
R32 VGND.n15 VGND.n14 4.65
R33 VGND.n19 VGND.n18 4.65
R34 VGND.n21 VGND.n20 4.65
R35 VGND.n23 VGND.n22 4.65
R36 VGND.n25 VGND.n24 4.65
R37 VGND.n27 VGND.n26 4.65
R38 VGND.n29 VGND.n28 4.65
R39 VGND.n33 VGND.n32 4.65
R40 VGND.n35 VGND.n34 4.65
R41 VGND.n8 VGND.n7 3.871
R42 VGND.n32 VGND.n31 3.764
R43 VGND.n18 VGND.n17 2.635
R44 VGND.n4 VGND.n3 0.609
R45 VGND.n5 VGND.n1 0.509
R46 VGND.n9 VGND.n5 0.119
R47 VGND.n11 VGND.n9 0.119
R48 VGND.n15 VGND.n11 0.119
R49 VGND.n19 VGND.n15 0.119
R50 VGND.n21 VGND.n19 0.119
R51 VGND.n23 VGND.n21 0.119
R52 VGND.n25 VGND.n23 0.119
R53 VGND.n27 VGND.n25 0.119
R54 VGND.n29 VGND.n27 0.119
R55 VGND.n33 VGND.n29 0.119
R56 VGND.n35 VGND.n33 0.119
R57 VGND.n37 VGND.n35 0.119
R58 VGND VGND.n37 0.02
R59 a_467_47.n6 a_467_47.t7 231.794
R60 a_467_47.n1 a_467_47.t3 182.431
R61 a_467_47.n3 a_467_47.n1 99.764
R62 a_467_47.n6 a_467_47.n5 63.9
R63 a_467_47.n5 a_467_47.n3 63.247
R64 a_467_47.n1 a_467_47.n0 51.506
R65 a_467_47.n3 a_467_47.n2 51.506
R66 a_467_47.n5 a_467_47.n4 51.506
R67 a_467_47.n0 a_467_47.t1 48
R68 a_467_47.n7 a_467_47.n6 42.273
R69 a_467_47.n0 a_467_47.t2 38.769
R70 a_467_47.n2 a_467_47.t0 28.615
R71 a_467_47.n7 a_467_47.t6 28.615
R72 a_467_47.n4 a_467_47.t5 24.923
R73 a_467_47.n4 a_467_47.t9 24.923
R74 a_467_47.n2 a_467_47.t4 24.923
R75 a_467_47.t8 a_467_47.n7 24.923
R76 VNB VNB.t13 6053.91
R77 VNB.t11 VNB.t7 4545.05
R78 VNB.t0 VNB.t1 3674.73
R79 VNB.t1 VNB.t2 2997.8
R80 VNB.t4 VNB.t0 2127.47
R81 VNB.t6 VNB.t8 2127.47
R82 VNB.t2 VNB.t3 2030.77
R83 VNB.t5 VNB.t4 2030.77
R84 VNB.t9 VNB.t5 2030.77
R85 VNB.t8 VNB.t9 2030.77
R86 VNB.t7 VNB.t6 2030.77
R87 VNB.t12 VNB.t11 2030.77
R88 VNB.t10 VNB.t12 2030.77
R89 VNB.t13 VNB.t10 2030.77
R90 A3.n0 A3.t2 221.719
R91 A3.n1 A3.t3 221.719
R92 A3.n0 A3.t0 149.419
R93 A3.n1 A3.t1 149.419
R94 A3.n3 A3.n2 76
R95 A3.n2 A3.n0 37.488
R96 A3.n2 A3.n1 37.488
R97 A3 A3.n3 16
R98 A3.n3 A3 13.44
R99 A1.n1 A1.t2 221.719
R100 A1.n2 A1.t1 221.719
R101 A1.n1 A1.t3 149.419
R102 A1.n2 A1.t0 149.419
R103 A1.n1 A1.n0 126.877
R104 A1.n4 A1.n3 76
R105 A1.n3 A1.n2 40.166
R106 A1.n3 A1.n1 34.811
R107 A1.n4 A1 17.6
R108 A1.n0 A1 15.04
R109 A1.n0 A1 13.12
R110 A1 A1.n4 11.84
R111 B1.n0 B1.t1 300.267
R112 B1.n0 B1.t3 221.719
R113 B1.n2 B1.t0 165.485
R114 B1.n1 B1.t2 149.419
R115 B1 B1.n2 80.48
R116 B1.n2 B1.n1 58.911
R117 B1.n1 B1.n0 14.281
R118 a_79_21.n11 a_79_21.n9 232.125
R119 a_79_21.n5 a_79_21.t6 221.719
R120 a_79_21.n6 a_79_21.t7 221.719
R121 a_79_21.n2 a_79_21.t8 221.719
R122 a_79_21.n0 a_79_21.t12 221.719
R123 a_79_21.n5 a_79_21.t10 149.419
R124 a_79_21.n6 a_79_21.t11 149.419
R125 a_79_21.n2 a_79_21.t9 149.419
R126 a_79_21.n0 a_79_21.t13 149.419
R127 a_79_21.n13 a_79_21.n12 122.64
R128 a_79_21.n11 a_79_21.n10 108.9
R129 a_79_21.n4 a_79_21.n1 100.436
R130 a_79_21.n4 a_79_21.n3 76
R131 a_79_21.n8 a_79_21.n7 76
R132 a_79_21.n12 a_79_21.n8 38.981
R133 a_79_21.n7 a_79_21.n6 38.381
R134 a_79_21.n3 a_79_21.n2 37.488
R135 a_79_21.n1 a_79_21.n0 37.488
R136 a_79_21.n7 a_79_21.n5 36.596
R137 a_79_21.n10 a_79_21.t3 30.535
R138 a_79_21.n10 a_79_21.t2 26.595
R139 a_79_21.n9 a_79_21.t1 26.595
R140 a_79_21.n9 a_79_21.t0 26.595
R141 a_79_21.t5 a_79_21.n13 24.923
R142 a_79_21.n13 a_79_21.t4 24.923
R143 a_79_21.n8 a_79_21.n4 24.727
R144 a_79_21.n12 a_79_21.n11 12.617
R145 A2.n0 A2.t1 229.752
R146 A2.n2 A2.t2 221.719
R147 A2.n6 A2.t3 164.593
R148 A2.n1 A2.t0 149.419
R149 A2.n6 A2.n5 77.655
R150 A2.n5 A2.n4 76
R151 A2.n7 A2.n6 76
R152 A2.n2 A2.n1 39.274
R153 A2.n1 A2.n0 27.67
R154 A2.n7 A2 26.56
R155 A2.n4 A2.n3 25.28
R156 A2.n5 A2.n2 3.57
R157 A2.n3 A2 2.88
R158 A2 A2.n7 2.88
R159 A2.n4 A2 1.28
R160 VPWR.n1 VPWR.t6 196.528
R161 VPWR.n17 VPWR.t2 195.621
R162 VPWR.n12 VPWR.n11 174.594
R163 VPWR.n2 VPWR.n0 170.327
R164 VPWR.n6 VPWR.n5 132.865
R165 VPWR.n11 VPWR.t4 26.595
R166 VPWR.n11 VPWR.t3 26.595
R167 VPWR.n5 VPWR.t7 26.595
R168 VPWR.n5 VPWR.t5 26.595
R169 VPWR.n0 VPWR.t0 26.595
R170 VPWR.n0 VPWR.t1 26.595
R171 VPWR.n7 VPWR.n6 9.788
R172 VPWR.n2 VPWR.n1 6.022
R173 VPWR.n4 VPWR.n3 4.65
R174 VPWR.n8 VPWR.n7 4.65
R175 VPWR.n10 VPWR.n9 4.65
R176 VPWR.n14 VPWR.n13 4.65
R177 VPWR.n16 VPWR.n15 4.65
R178 VPWR.n18 VPWR.n17 4.65
R179 VPWR.n13 VPWR.n12 3.764
R180 VPWR.n4 VPWR.n2 0.134
R181 VPWR.n8 VPWR.n4 0.119
R182 VPWR.n10 VPWR.n8 0.119
R183 VPWR.n14 VPWR.n10 0.119
R184 VPWR.n16 VPWR.n14 0.119
R185 VPWR.n18 VPWR.n16 0.119
R186 VPWR VPWR.n18 0.02
R187 VPB.t11 VPB.t0 580.062
R188 VPB.t12 VPB.t8 556.386
R189 VPB.t13 VPB.t12 260.436
R190 VPB.t3 VPB.t2 248.598
R191 VPB.t1 VPB.t3 248.598
R192 VPB.t0 VPB.t1 248.598
R193 VPB.t10 VPB.t11 248.598
R194 VPB.t9 VPB.t10 248.598
R195 VPB.t8 VPB.t9 248.598
R196 VPB.t7 VPB.t13 248.598
R197 VPB.t6 VPB.t7 248.598
R198 VPB.t5 VPB.t6 248.598
R199 VPB.t4 VPB.t5 248.598
R200 VPB VPB.t4 189.408
R201 a_1083_297.n1 a_1083_297.t1 238.015
R202 a_1083_297.t2 a_1083_297.n1 236.789
R203 a_1083_297.n1 a_1083_297.n0 110.507
R204 a_1083_297.n0 a_1083_297.t3 26.595
R205 a_1083_297.n0 a_1083_297.t0 26.595
R206 X.n5 X.n3 140.856
R207 X.n5 X.n4 108.216
R208 X.n2 X.n0 87.175
R209 X.n2 X.n1 52.818
R210 X.n3 X.t7 26.595
R211 X.n3 X.t6 26.595
R212 X.n4 X.t5 26.595
R213 X.n4 X.t4 26.595
R214 X.n0 X.t2 24.923
R215 X.n0 X.t1 24.923
R216 X.n1 X.t3 24.923
R217 X.n1 X.t0 24.923
R218 X X.n5 16.787
R219 X.n6 X 14.523
R220 X.n6 X.n2 11.452
R221 X X.n6 2.215
R222 a_889_297.n1 a_889_297.n0 398.711
R223 a_889_297.n0 a_889_297.t3 26.595
R224 a_889_297.n0 a_889_297.t2 26.595
R225 a_889_297.t1 a_889_297.n1 26.595
R226 a_889_297.n1 a_889_297.t0 26.595
R227 a_639_297.n0 a_639_297.t0 239.197
R228 a_639_297.n0 a_639_297.t3 233.296
R229 a_639_297.n1 a_639_297.n0 91.914
R230 a_639_297.n1 a_639_297.t2 26.595
R231 a_639_297.t1 a_639_297.n1 26.595
C0 VPWR VGND 0.17fF
C1 X VGND 0.48fF
C2 VPB VPWR 0.16fF
C3 VPWR X 0.71fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__o41ai_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__o41ai_1 A1 A2 A3 A4 Y B1 VGND VPWR VNB VPB
X0 a_348_297.t1 A3.t0 a_193_297.t1 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_109_47.t0 A1.t0 VGND.t0 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 a_193_297.t0 A4.t0 Y.t0 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 VPWR.t0 A1.t1 a_432_297.t0 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 VGND.t2 A4.t1 a_109_47.t2 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 VGND.t1 A2.t0 a_109_47.t1 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 a_109_47.t4 A3.t1 VGND.t3 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 a_432_297.t1 A2.t1 a_348_297.t0 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 Y.t1 B1.t0 VPWR.t1 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 a_109_47.t3 B1.t1 Y.t2 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
R0 A3.n0 A3.t0 241.534
R1 A3.n0 A3.t1 169.234
R2 A3.n1 A3.n0 76
R3 A3.n1 A3 11.4
R4 A3 A3.n1 2.2
R5 a_193_297.t0 a_193_297.t1 123.125
R6 a_348_297.t0 a_348_297.t1 53.19
R7 VPB.t1 VPB.t4 458.722
R8 VPB.t3 VPB.t2 295.95
R9 VPB.t4 VPB.t3 248.598
R10 VPB.t0 VPB.t1 248.598
R11 VPB VPB.t0 189.408
R12 A1.n0 A1.t1 239.503
R13 A1.n0 A1.t0 167.203
R14 A1 A1.n0 88.544
R15 VGND.n2 VGND.n1 117.78
R16 VGND.n2 VGND.n0 117.538
R17 VGND.n1 VGND.t1 39.692
R18 VGND.n1 VGND.t0 24.923
R19 VGND.n0 VGND.t3 24.923
R20 VGND.n0 VGND.t2 24.923
R21 VGND VGND.n2 0.451
R22 a_109_47.t0 a_109_47.n2 133.933
R23 a_109_47.n2 a_109_47.n0 99.065
R24 a_109_47.n0 a_109_47.t3 83.215
R25 a_109_47.n2 a_109_47.n1 53.206
R26 a_109_47.n0 a_109_47.t2 31.173
R27 a_109_47.n1 a_109_47.t1 24.923
R28 a_109_47.n1 a_109_47.t4 24.923
R29 VNB VNB.t3 6053.91
R30 VNB.t3 VNB.t2 3747.25
R31 VNB.t1 VNB.t0 2417.58
R32 VNB.t4 VNB.t1 2030.77
R33 VNB.t2 VNB.t4 2030.77
R34 A4.n0 A4.t0 269.026
R35 A4.n0 A4.t1 165.485
R36 A4.n1 A4.n0 76
R37 A4.n1 A4 11.96
R38 A4 A4.n1 2.308
R39 Y Y.n0 139.93
R40 Y.n1 Y.t2 83.131
R41 Y.n0 Y.t0 26.595
R42 Y.n0 Y.t1 26.595
R43 Y Y.n1 22.901
R44 Y Y.n2 15.058
R45 Y.n2 Y 10.541
R46 Y.n2 Y 6.4
R47 Y.n1 Y 5.55
R48 a_432_297.t0 a_432_297.t1 68.95
R49 VPWR.n0 VPWR.t1 155.644
R50 VPWR.n0 VPWR.t0 150.825
R51 VPWR VPWR.n0 0.038
R52 A2.n0 A2.t1 239.503
R53 A2.n0 A2.t0 167.203
R54 A2 A2.n0 87.019
R55 B1.n0 B1.t0 234.39
R56 B1.n0 B1.t1 162.09
R57 B1 B1.n0 84
C0 VPWR Y 0.23fF
C1 A2 VPWR 0.12fF
C2 A3 A2 0.27fF
C3 B1 Y 0.10fF
C4 A4 A3 0.25fF
C5 A4 Y 0.13fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__o41ai_2.ext - technology: sky130A

.subckt sky130_fd_sc_hd__o41ai_2 A1 A2 A3 A4 Y B1 VGND VPWR VNB VPB
X0 a_27_47.t1 A2.t0 VGND.t0 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 VGND.t6 A4.t0 a_27_47.t8 VNB.t8 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 VGND.t2 A3.t0 a_27_47.t2 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 VGND.t1 A2.t1 a_27_47.t0 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 VGND.t4 A1.t0 a_27_47.t6 VNB.t6 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 a_27_47.t3 A3.t1 VGND.t3 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 VPWR.t1 B1.t0 Y.t1 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 a_27_47.t4 B1.t1 Y.t3 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 a_299_297.t1 A3.t2 a_549_297.t3 VPB.t7 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 a_549_297.t2 A3.t3 a_299_297.t0 VPB.t6 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 a_299_297.t3 A4.t1 Y.t5 VPB.t9 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 Y.t4 A4.t2 a_299_297.t2 VPB.t8 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 a_743_297.t3 A1.t1 VPWR.t3 VPB.t5 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13 VPWR.t2 A1.t2 a_743_297.t2 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14 a_743_297.t1 A2.t2 a_549_297.t1 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 a_27_47.t9 A4.t3 VGND.t7 VNB.t9 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X16 Y.t0 B1.t2 VPWR.t0 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17 a_27_47.t7 A1.t3 VGND.t5 VNB.t7 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X18 a_549_297.t0 A2.t3 a_743_297.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X19 Y.t2 B1.t3 a_27_47.t5 VNB.t5 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
R0 A2.n0 A2.t2 221.719
R1 A2.n3 A2.t3 221.719
R2 A2.n0 A2.t0 138.173
R3 A2.n3 A2.t1 138.173
R4 A2.n4 A2.n3 95.754
R5 A2.n2 A2.n1 76
R6 A2.n1 A2.n0 26.865
R7 A2.n4 A2.n2 24
R8 A2 A2.n4 4.8
R9 A2.n2 A2 0.64
R10 VGND.n16 VGND.t7 195.032
R11 VGND.n6 VGND.t2 190.339
R12 VGND.n3 VGND.n0 124.921
R13 VGND.n2 VGND.n1 114.711
R14 VGND.n11 VGND.n10 114.711
R15 VGND.n0 VGND.t5 24.923
R16 VGND.n0 VGND.t4 24.923
R17 VGND.n1 VGND.t0 24.923
R18 VGND.n1 VGND.t1 24.923
R19 VGND.n10 VGND.t3 24.923
R20 VGND.n10 VGND.t6 24.923
R21 VGND.n3 VGND.n2 10.723
R22 VGND.n12 VGND.n11 5.27
R23 VGND.n5 VGND.n4 4.65
R24 VGND.n7 VGND.n6 4.65
R25 VGND.n9 VGND.n8 4.65
R26 VGND.n13 VGND.n12 4.65
R27 VGND.n15 VGND.n14 4.65
R28 VGND.n17 VGND.n16 3.953
R29 VGND VGND.n17 0.359
R30 VGND.n5 VGND.n3 0.327
R31 VGND.n17 VGND.n15 0.139
R32 VGND.n7 VGND.n5 0.119
R33 VGND.n9 VGND.n7 0.119
R34 VGND.n13 VGND.n9 0.119
R35 VGND.n15 VGND.n13 0.119
R36 a_27_47.n0 a_27_47.t5 140.979
R37 a_27_47.n6 a_27_47.t7 127.91
R38 a_27_47.n5 a_27_47.t0 89.51
R39 a_27_47.n0 a_27_47.t4 81.281
R40 a_27_47.n2 a_27_47.n0 59.108
R41 a_27_47.n2 a_27_47.n1 53.206
R42 a_27_47.n4 a_27_47.n3 53.206
R43 a_27_47.n7 a_27_47.n6 53.205
R44 a_27_47.n5 a_27_47.n4 48.941
R45 a_27_47.n4 a_27_47.n2 38.4
R46 a_27_47.n6 a_27_47.n5 38.4
R47 a_27_47.n1 a_27_47.t8 24.923
R48 a_27_47.n1 a_27_47.t9 24.923
R49 a_27_47.n3 a_27_47.t2 24.923
R50 a_27_47.n3 a_27_47.t3 24.923
R51 a_27_47.n7 a_27_47.t6 24.923
R52 a_27_47.t1 a_27_47.n7 24.923
R53 VNB VNB.t5 6053.91
R54 VNB.t2 VNB.t0 4738.46
R55 VNB.t4 VNB.t9 4545.05
R56 VNB.t6 VNB.t7 2030.77
R57 VNB.t1 VNB.t6 2030.77
R58 VNB.t0 VNB.t1 2030.77
R59 VNB.t3 VNB.t2 2030.77
R60 VNB.t8 VNB.t3 2030.77
R61 VNB.t9 VNB.t8 2030.77
R62 VNB.t5 VNB.t4 2030.77
R63 A4.n2 A4.t2 235.167
R64 A4.n0 A4.t1 218.506
R65 A4.n3 A4.t3 163.462
R66 A4.n0 A4.t0 149.419
R67 A4 A4.n1 84.64
R68 A4.n4 A4.n3 76
R69 A4 A4.n4 22.08
R70 A4.n1 A4.n0 18.075
R71 A4.n4 A4 7.36
R72 A4.n3 A4.n2 0.595
R73 A3.n0 A3.t2 216.899
R74 A3.n1 A3.t3 216.899
R75 A3.n0 A3.t0 144.599
R76 A3.n1 A3.t1 144.599
R77 A3.n3 A3.n0 90.46
R78 A3 A3.n2 86.88
R79 A3.n2 A3.n0 53.02
R80 A3.n3 A3 16
R81 A3.n2 A3.n1 14.46
R82 A3 A3.n3 13.44
R83 A1.n1 A1.t1 221.719
R84 A1.n2 A1.t2 221.719
R85 A1.n1 A1.t3 149.419
R86 A1.n2 A1.t0 149.419
R87 A1.n1 A1.n0 118.844
R88 A1.n4 A1.n3 76
R89 A1.n3 A1.n2 38.381
R90 A1.n3 A1.n1 36.596
R91 A1 A1.n4 21.44
R92 A1.n0 A1 20.48
R93 A1.n0 A1 8.96
R94 A1.n4 A1 8
R95 B1.n0 B1.t0 216.899
R96 B1.n1 B1.t2 216.899
R97 B1.n0 B1.t1 141.386
R98 B1.n1 B1.t3 141.386
R99 B1 B1.n1 115.605
R100 B1.n1 B1.n0 65.303
R101 Y.n2 Y.n0 213.474
R102 Y.n2 Y.n1 112.936
R103 Y Y.n3 94.245
R104 Y.n1 Y.t1 26.595
R105 Y.n1 Y.t0 26.595
R106 Y.n0 Y.t5 26.595
R107 Y.n0 Y.t4 26.595
R108 Y.n3 Y.t3 24.923
R109 Y.n3 Y.t2 24.923
R110 Y Y.n4 11.982
R111 Y.n4 Y 6.536
R112 Y Y.n2 5.991
R113 Y.n4 Y 4.654
R114 VPWR.n1 VPWR.t1 196.528
R115 VPWR.n2 VPWR.n0 168.612
R116 VPWR.n5 VPWR.t0 151.631
R117 VPWR.n0 VPWR.t3 26.595
R118 VPWR.n0 VPWR.t2 26.595
R119 VPWR.n4 VPWR.n3 4.65
R120 VPWR.n6 VPWR.n5 4.65
R121 VPWR.n2 VPWR.n1 4.013
R122 VPWR.n4 VPWR.n2 0.137
R123 VPWR.n6 VPWR.n4 0.119
R124 VPWR VPWR.n6 0.02
R125 VPB.t7 VPB.t0 580.062
R126 VPB.t3 VPB.t8 556.386
R127 VPB.t4 VPB.t5 248.598
R128 VPB.t1 VPB.t4 248.598
R129 VPB.t0 VPB.t1 248.598
R130 VPB.t6 VPB.t7 248.598
R131 VPB.t9 VPB.t6 248.598
R132 VPB.t8 VPB.t9 248.598
R133 VPB.t2 VPB.t3 248.598
R134 VPB VPB.t2 189.408
R135 a_549_297.n1 a_549_297.n0 382.615
R136 a_549_297.n0 a_549_297.t3 26.595
R137 a_549_297.n0 a_549_297.t2 26.595
R138 a_549_297.n1 a_549_297.t1 26.595
R139 a_549_297.t0 a_549_297.n1 26.595
R140 a_299_297.t1 a_299_297.n1 262.34
R141 a_299_297.n1 a_299_297.t2 259.292
R142 a_299_297.n1 a_299_297.n0 87.183
R143 a_299_297.n0 a_299_297.t0 26.595
R144 a_299_297.n0 a_299_297.t3 26.595
R145 a_743_297.n0 a_743_297.t0 238.015
R146 a_743_297.n0 a_743_297.t3 194.203
R147 a_743_297.n1 a_743_297.n0 110.508
R148 a_743_297.n1 a_743_297.t2 26.595
R149 a_743_297.t1 a_743_297.n1 26.595
C0 VPB VPWR 0.12fF
C1 VPWR Y 0.40fF
C2 VPWR VGND 0.13fF
C3 A4 Y 0.14fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__o41ai_4.ext - technology: sky130A

.subckt sky130_fd_sc_hd__o41ai_4 A1 A2 A3 A4 Y B1 VGND VPWR VNB VPB
X0 VGND.t13 A2.t0 a_27_47.t17 VNB.t17 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 a_467_297.t3 A4.t0 Y.t10 VPB.t13 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 VGND.t12 A2.t1 a_27_47.t16 VNB.t16 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 VPWR.t7 A1.t0 a_1243_297.t7 VPB.t18 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 VGND.t15 A1.t1 a_27_47.t19 VNB.t19 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 a_27_47.t1 A4.t1 VGND.t1 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 Y.t9 A4.t2 a_467_297.t2 VPB.t12 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 a_27_47.t2 A4.t3 VGND.t2 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 VPWR.t3 B1.t0 Y.t11 VPB.t19 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 a_27_47.t15 A2.t2 VGND.t11 VNB.t15 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 a_27_47.t14 A2.t3 VGND.t10 VNB.t14 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 VGND.t3 A4.t4 a_27_47.t3 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 a_27_47.t0 A1.t2 VGND.t0 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 VGND.t5 A3.t0 a_27_47.t5 VNB.t5 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14 Y.t0 B1.t1 VPWR.t0 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 a_1243_297.t6 A1.t3 VPWR.t6 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16 a_27_47.t8 A1.t4 VGND.t8 VNB.t8 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X17 VGND.t4 A4.t5 a_27_47.t4 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X18 VGND.t6 A3.t1 a_27_47.t6 VNB.t6 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X19 VPWR.t1 B1.t2 Y.t1 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X20 VPWR.t5 A1.t5 a_1243_297.t5 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X21 a_27_47.t10 B1.t3 Y.t2 VNB.t10 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X22 a_27_47.t11 B1.t4 Y.t3 VNB.t11 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X23 a_467_297.t1 A4.t6 Y.t8 VPB.t11 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X24 a_1243_297.t0 A2.t4 a_885_297.t3 VPB.t9 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X25 Y.t7 A4.t7 a_467_297.t0 VPB.t10 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X26 a_27_47.t7 A3.t2 VGND.t7 VNB.t7 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X27 VGND.t9 A1.t6 a_27_47.t9 VNB.t9 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X28 a_885_297.t2 A2.t5 a_1243_297.t3 VPB.t8 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X29 a_27_47.t18 A3.t3 VGND.t14 VNB.t18 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X30 Y.t4 B1.t5 a_27_47.t12 VNB.t12 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X31 a_1243_297.t2 A2.t6 a_885_297.t1 VPB.t7 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X32 a_467_297.t4 A3.t4 a_885_297.t7 VPB.t14 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X33 a_885_297.t0 A2.t7 a_1243_297.t1 VPB.t6 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X34 a_885_297.t6 A3.t5 a_467_297.t5 VPB.t15 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X35 a_467_297.t6 A3.t6 a_885_297.t5 VPB.t16 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X36 Y.t5 B1.t6 VPWR.t2 VPB.t5 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X37 a_1243_297.t4 A1.t7 VPWR.t4 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X38 a_885_297.t4 A3.t7 a_467_297.t7 VPB.t17 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X39 Y.t6 B1.t7 a_27_47.t13 VNB.t13 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
R0 A2.n6 A2.t6 221.719
R1 A2.n1 A2.t4 221.719
R2 A2.n2 A2.t5 221.719
R3 A2.n7 A2.t7 221.719
R4 A2.n6 A2.t2 149.419
R5 A2.n1 A2.t3 149.419
R6 A2.n2 A2.t1 149.419
R7 A2.n7 A2.t0 149.419
R8 A2 A2.n3 90.4
R9 A2.n8 A2.n7 79.57
R10 A2.n4 A2.n0 76
R11 A2.n6 A2.n5 76
R12 A2.n7 A2.n6 74.977
R13 A2.n6 A2.n0 71.407
R14 A2.n3 A2.n2 68.729
R15 A2 A2.n8 23.04
R16 A2.n5 A2 21.76
R17 A2 A2.n4 17.92
R18 A2.n4 A2 11.52
R19 A2.n5 A2 7.68
R20 A2.n8 A2 6.4
R21 A2.n3 A2.n1 6.248
R22 A2.n2 A2.n0 3.57
R23 a_27_47.n2 a_27_47.t11 175.576
R24 a_27_47.n1 a_27_47.t13 136.63
R25 a_27_47.n16 a_27_47.t8 127.91
R26 a_27_47.n1 a_27_47.n0 92.5
R27 a_27_47.n10 a_27_47.t7 92.303
R28 a_27_47.n11 a_27_47.t17 92.303
R29 a_27_47.n3 a_27_47.t3 81.64
R30 a_27_47.n5 a_27_47.n4 53.206
R31 a_27_47.n7 a_27_47.n6 53.206
R32 a_27_47.n9 a_27_47.n8 53.206
R33 a_27_47.n13 a_27_47.n12 53.206
R34 a_27_47.n15 a_27_47.n14 53.206
R35 a_27_47.n17 a_27_47.n16 53.205
R36 a_27_47.n2 a_27_47.n1 51.2
R37 a_27_47.n5 a_27_47.n3 50.413
R38 a_27_47.n7 a_27_47.n5 38.4
R39 a_27_47.n9 a_27_47.n7 38.4
R40 a_27_47.n10 a_27_47.n9 38.4
R41 a_27_47.n13 a_27_47.n11 38.4
R42 a_27_47.n15 a_27_47.n13 38.4
R43 a_27_47.n16 a_27_47.n15 38.4
R44 a_27_47.n3 a_27_47.n2 33.687
R45 a_27_47.n0 a_27_47.t12 24.923
R46 a_27_47.n0 a_27_47.t10 24.923
R47 a_27_47.n4 a_27_47.t4 24.923
R48 a_27_47.n4 a_27_47.t1 24.923
R49 a_27_47.n6 a_27_47.t6 24.923
R50 a_27_47.n6 a_27_47.t2 24.923
R51 a_27_47.n8 a_27_47.t5 24.923
R52 a_27_47.n8 a_27_47.t18 24.923
R53 a_27_47.n12 a_27_47.t16 24.923
R54 a_27_47.n12 a_27_47.t15 24.923
R55 a_27_47.n14 a_27_47.t19 24.923
R56 a_27_47.n14 a_27_47.t14 24.923
R57 a_27_47.n17 a_27_47.t9 24.923
R58 a_27_47.t0 a_27_47.n17 24.923
R59 a_27_47.n11 a_27_47.n10 14.305
R60 VGND.n3 VGND.n0 124.575
R61 VGND.n2 VGND.n1 114.711
R62 VGND.n7 VGND.n6 114.711
R63 VGND.n13 VGND.n12 114.711
R64 VGND.n21 VGND.n20 114.711
R65 VGND.n27 VGND.n26 114.711
R66 VGND.n31 VGND.n30 114.711
R67 VGND.n37 VGND.n36 114.711
R68 VGND.n0 VGND.t8 24.923
R69 VGND.n0 VGND.t9 24.923
R70 VGND.n1 VGND.t0 24.923
R71 VGND.n1 VGND.t15 24.923
R72 VGND.n6 VGND.t10 24.923
R73 VGND.n6 VGND.t12 24.923
R74 VGND.n12 VGND.t11 24.923
R75 VGND.n12 VGND.t13 24.923
R76 VGND.n20 VGND.t7 24.923
R77 VGND.n20 VGND.t5 24.923
R78 VGND.n26 VGND.t14 24.923
R79 VGND.n26 VGND.t6 24.923
R80 VGND.n30 VGND.t2 24.923
R81 VGND.n30 VGND.t4 24.923
R82 VGND.n36 VGND.t1 24.923
R83 VGND.n36 VGND.t3 24.923
R84 VGND.n28 VGND.n27 14.305
R85 VGND.n32 VGND.n31 14.305
R86 VGND.n3 VGND.n2 9.234
R87 VGND.n22 VGND.n21 8.282
R88 VGND.n38 VGND.n37 8.282
R89 VGND.n14 VGND.n13 6.776
R90 VGND.n5 VGND.n4 4.65
R91 VGND.n9 VGND.n8 4.65
R92 VGND.n11 VGND.n10 4.65
R93 VGND.n15 VGND.n14 4.65
R94 VGND.n17 VGND.n16 4.65
R95 VGND.n19 VGND.n18 4.65
R96 VGND.n23 VGND.n22 4.65
R97 VGND.n25 VGND.n24 4.65
R98 VGND.n29 VGND.n28 4.65
R99 VGND.n33 VGND.n32 4.65
R100 VGND.n35 VGND.n34 4.65
R101 VGND.n39 VGND.n38 4.65
R102 VGND.n8 VGND.n7 0.752
R103 VGND VGND.n40 0.603
R104 VGND.n5 VGND.n3 0.31
R105 VGND.n40 VGND.n39 0.134
R106 VGND.n9 VGND.n5 0.119
R107 VGND.n11 VGND.n9 0.119
R108 VGND.n15 VGND.n11 0.119
R109 VGND.n17 VGND.n15 0.119
R110 VGND.n19 VGND.n17 0.119
R111 VGND.n23 VGND.n19 0.119
R112 VGND.n25 VGND.n23 0.119
R113 VGND.n29 VGND.n25 0.119
R114 VGND.n33 VGND.n29 0.119
R115 VGND.n35 VGND.n33 0.119
R116 VGND.n39 VGND.n35 0.119
R117 VNB VNB.t13 6053.91
R118 VNB.t7 VNB.t17 4545.05
R119 VNB.t11 VNB.t3 4545.05
R120 VNB.t9 VNB.t8 2030.77
R121 VNB.t0 VNB.t9 2030.77
R122 VNB.t19 VNB.t0 2030.77
R123 VNB.t14 VNB.t19 2030.77
R124 VNB.t16 VNB.t14 2030.77
R125 VNB.t15 VNB.t16 2030.77
R126 VNB.t17 VNB.t15 2030.77
R127 VNB.t5 VNB.t7 2030.77
R128 VNB.t18 VNB.t5 2030.77
R129 VNB.t6 VNB.t18 2030.77
R130 VNB.t2 VNB.t6 2030.77
R131 VNB.t4 VNB.t2 2030.77
R132 VNB.t1 VNB.t4 2030.77
R133 VNB.t3 VNB.t1 2030.77
R134 VNB.t12 VNB.t11 2030.77
R135 VNB.t10 VNB.t12 2030.77
R136 VNB.t13 VNB.t10 2030.77
R137 A4.n9 A4.t7 232.213
R138 A4.n1 A4.t0 221.719
R139 A4.n0 A4.t2 221.719
R140 A4.n6 A4.t6 221.719
R141 A4.n9 A4.t4 159.913
R142 A4.n1 A4.t3 149.419
R143 A4.n0 A4.t5 149.419
R144 A4.n6 A4.t1 149.419
R145 A4.n3 A4.n2 76
R146 A4.n5 A4.n4 76
R147 A4.n8 A4.n7 76
R148 A4.n10 A4.n9 76
R149 A4.n2 A4.n1 37.488
R150 A4.n2 A4.n0 37.488
R151 A4.n5 A4.n0 37.488
R152 A4.n6 A4.n5 37.488
R153 A4.n7 A4.n6 36.596
R154 A4.n4 A4 23.68
R155 A4.n10 A4.n8 23.68
R156 A4 A4.n3 21.12
R157 A4.n3 A4 8.32
R158 A4.n4 A4 5.76
R159 A4.n8 A4 2.88
R160 A4 A4.n10 2.88
R161 Y.n6 Y.n4 192.917
R162 Y.n6 Y.n5 154.517
R163 Y.n10 Y.n9 132.322
R164 Y.n1 Y.n0 109.574
R165 Y.n3 Y.n2 109.574
R166 Y.n10 Y.n8 92.5
R167 Y.n7 Y.n6 41.788
R168 Y.n4 Y.t10 26.595
R169 Y.n4 Y.t9 26.595
R170 Y.n5 Y.t8 26.595
R171 Y.n5 Y.t7 26.595
R172 Y.n0 Y.t1 26.595
R173 Y.n0 Y.t5 26.595
R174 Y.n2 Y.t11 26.595
R175 Y.n2 Y.t0 26.595
R176 Y.n8 Y.t3 24.923
R177 Y.n8 Y.t4 24.923
R178 Y.n9 Y.t2 24.923
R179 Y.n9 Y.t6 24.923
R180 Y.n3 Y 21.458
R181 Y Y.n1 16.941
R182 Y.n11 Y.n10 16.592
R183 Y Y.n11 14.786
R184 Y.n7 Y.n3 13.929
R185 Y.n3 Y 11.67
R186 Y Y.n7 3.751
R187 Y.n1 Y 3.296
R188 Y.n3 Y 3.296
R189 Y.n11 Y 0.22
R190 a_467_297.n3 a_467_297.t0 238.527
R191 a_467_297.n1 a_467_297.t4 219.512
R192 a_467_297.n1 a_467_297.n0 154.517
R193 a_467_297.n3 a_467_297.n2 152.759
R194 a_467_297.n5 a_467_297.n4 87.182
R195 a_467_297.n4 a_467_297.n3 87.062
R196 a_467_297.n4 a_467_297.n1 74.149
R197 a_467_297.n2 a_467_297.t2 26.595
R198 a_467_297.n2 a_467_297.t1 26.595
R199 a_467_297.n0 a_467_297.t5 26.595
R200 a_467_297.n0 a_467_297.t6 26.595
R201 a_467_297.n5 a_467_297.t7 26.595
R202 a_467_297.t3 a_467_297.n5 26.595
R203 VPB.t14 VPB.t6 556.386
R204 VPB.t19 VPB.t10 556.386
R205 VPB.t18 VPB.t2 248.598
R206 VPB.t0 VPB.t18 248.598
R207 VPB.t1 VPB.t0 248.598
R208 VPB.t9 VPB.t1 248.598
R209 VPB.t8 VPB.t9 248.598
R210 VPB.t7 VPB.t8 248.598
R211 VPB.t6 VPB.t7 248.598
R212 VPB.t15 VPB.t14 248.598
R213 VPB.t16 VPB.t15 248.598
R214 VPB.t17 VPB.t16 248.598
R215 VPB.t13 VPB.t17 248.598
R216 VPB.t12 VPB.t13 248.598
R217 VPB.t11 VPB.t12 248.598
R218 VPB.t10 VPB.t11 248.598
R219 VPB.t3 VPB.t19 248.598
R220 VPB.t4 VPB.t3 248.598
R221 VPB.t5 VPB.t4 248.598
R222 VPB VPB.t5 189.408
R223 A1.n0 A1.t7 221.719
R224 A1.n4 A1.t0 221.719
R225 A1.n5 A1.t3 221.719
R226 A1.n8 A1.t5 221.719
R227 A1.n0 A1.t4 149.419
R228 A1.n4 A1.t6 149.419
R229 A1.n5 A1.t2 149.419
R230 A1.n8 A1.t1 149.419
R231 A1 A1.n9 85.6
R232 A1.n1 A1.n0 84.033
R233 A1.n3 A1.n2 76
R234 A1.n7 A1.n6 76
R235 A1.n3 A1.n0 70.514
R236 A1.n6 A1.n4 63.374
R237 A1.n1 A1 20.16
R238 A1.n2 A1 18.88
R239 A1.n9 A1.n8 16.066
R240 A1 A1.n7 15.68
R241 A1.n7 A1 13.76
R242 A1.n6 A1.n5 11.603
R243 A1.n2 A1 10.56
R244 A1 A1.n1 9.28
R245 A1.n4 A1.n3 4.462
R246 a_1243_297.n1 a_1243_297.t1 219.512
R247 a_1243_297.n3 a_1243_297.t4 174.569
R248 a_1243_297.n1 a_1243_297.n0 154.517
R249 a_1243_297.n5 a_1243_297.n4 109.574
R250 a_1243_297.n3 a_1243_297.n2 109.574
R251 a_1243_297.n4 a_1243_297.n1 38.4
R252 a_1243_297.n4 a_1243_297.n3 38.4
R253 a_1243_297.n2 a_1243_297.t7 26.595
R254 a_1243_297.n2 a_1243_297.t6 26.595
R255 a_1243_297.n0 a_1243_297.t3 26.595
R256 a_1243_297.n0 a_1243_297.t2 26.595
R257 a_1243_297.n5 a_1243_297.t5 26.595
R258 a_1243_297.t0 a_1243_297.n5 26.595
R259 VPWR.n30 VPWR.t3 196.528
R260 VPWR.n3 VPWR.n0 184.458
R261 VPWR.n35 VPWR.n34 174.594
R262 VPWR.n2 VPWR.n1 174.594
R263 VPWR.n40 VPWR.t2 151.631
R264 VPWR.n34 VPWR.t0 26.595
R265 VPWR.n34 VPWR.t1 26.595
R266 VPWR.n1 VPWR.t6 26.595
R267 VPWR.n1 VPWR.t5 26.595
R268 VPWR.n0 VPWR.t4 26.595
R269 VPWR.n0 VPWR.t7 26.595
R270 VPWR.n3 VPWR.n2 9.234
R271 VPWR.n5 VPWR.n4 4.65
R272 VPWR.n7 VPWR.n6 4.65
R273 VPWR.n9 VPWR.n8 4.65
R274 VPWR.n11 VPWR.n10 4.65
R275 VPWR.n13 VPWR.n12 4.65
R276 VPWR.n15 VPWR.n14 4.65
R277 VPWR.n17 VPWR.n16 4.65
R278 VPWR.n19 VPWR.n18 4.65
R279 VPWR.n21 VPWR.n20 4.65
R280 VPWR.n23 VPWR.n22 4.65
R281 VPWR.n25 VPWR.n24 4.65
R282 VPWR.n27 VPWR.n26 4.65
R283 VPWR.n29 VPWR.n28 4.65
R284 VPWR.n31 VPWR.n30 4.65
R285 VPWR.n33 VPWR.n32 4.65
R286 VPWR.n37 VPWR.n36 4.65
R287 VPWR.n39 VPWR.n38 4.65
R288 VPWR.n41 VPWR.n40 4.65
R289 VPWR.n36 VPWR.n35 3.764
R290 VPWR.n5 VPWR.n3 0.31
R291 VPWR.n7 VPWR.n5 0.119
R292 VPWR.n9 VPWR.n7 0.119
R293 VPWR.n11 VPWR.n9 0.119
R294 VPWR.n13 VPWR.n11 0.119
R295 VPWR.n15 VPWR.n13 0.119
R296 VPWR.n17 VPWR.n15 0.119
R297 VPWR.n19 VPWR.n17 0.119
R298 VPWR.n21 VPWR.n19 0.119
R299 VPWR.n23 VPWR.n21 0.119
R300 VPWR.n25 VPWR.n23 0.119
R301 VPWR.n27 VPWR.n25 0.119
R302 VPWR.n29 VPWR.n27 0.119
R303 VPWR.n31 VPWR.n29 0.119
R304 VPWR.n33 VPWR.n31 0.119
R305 VPWR.n37 VPWR.n33 0.119
R306 VPWR.n39 VPWR.n37 0.119
R307 VPWR.n41 VPWR.n39 0.119
R308 VPWR VPWR.n41 0.02
R309 B1.n9 B1.t6 234.39
R310 B1.n2 B1.t0 221.719
R311 B1.n4 B1.t1 221.719
R312 B1.n0 B1.t2 221.719
R313 B1.n9 B1.t7 162.09
R314 B1.n2 B1.t4 149.419
R315 B1.n4 B1.t5 149.419
R316 B1.n0 B1.t3 149.419
R317 B1.n6 B1.n5 76
R318 B1.n8 B1.n7 76
R319 B1.n10 B1.n9 76
R320 B1.n3 B1.n2 37.488
R321 B1.n4 B1.n3 37.488
R322 B1.n5 B1.n4 37.488
R323 B1.n5 B1.n0 37.488
R324 B1.n8 B1.n0 37.488
R325 B1.n6 B1.n1 26.88
R326 B1.n7 B1 24.96
R327 B1.n9 B1.n8 24.1
R328 B1.n10 B1 21.44
R329 B1 B1.n10 8
R330 B1.n7 B1 4.48
R331 B1 B1.n6 1.92
R332 B1.n1 B1 0.64
R333 A3.n1 A3.t4 221.719
R334 A3.n0 A3.t5 221.719
R335 A3.n6 A3.t6 221.719
R336 A3.n7 A3.t7 221.719
R337 A3.n1 A3.t2 149.419
R338 A3.n0 A3.t0 149.419
R339 A3.n6 A3.t3 149.419
R340 A3.n7 A3.t1 149.419
R341 A3.n1 A3 120.596
R342 A3.n3 A3.n2 76
R343 A3.n5 A3.n4 76
R344 A3.n9 A3.n8 76
R345 A3.n5 A3.n0 38.381
R346 A3.n2 A3.n1 37.488
R347 A3.n2 A3.n0 37.488
R348 A3.n8 A3.n6 37.488
R349 A3.n8 A3.n7 37.488
R350 A3.n6 A3.n5 36.596
R351 A3.n3 A3 18.56
R352 A3.n4 A3 16.32
R353 A3 A3.n9 16
R354 A3.n9 A3 13.44
R355 A3.n4 A3 13.12
R356 A3 A3.n3 10.88
R357 a_885_297.n5 a_885_297.n4 216.005
R358 a_885_297.n3 a_885_297.n2 211.932
R359 a_885_297.n3 a_885_297.n1 152.759
R360 a_885_297.n4 a_885_297.n0 152.759
R361 a_885_297.n4 a_885_297.n3 102.4
R362 a_885_297.n2 a_885_297.t5 26.595
R363 a_885_297.n2 a_885_297.t4 26.595
R364 a_885_297.n1 a_885_297.t7 26.595
R365 a_885_297.n1 a_885_297.t6 26.595
R366 a_885_297.n0 a_885_297.t1 26.595
R367 a_885_297.n0 a_885_297.t0 26.595
R368 a_885_297.t3 a_885_297.n5 26.595
R369 a_885_297.n5 a_885_297.t2 26.595
C0 A4 Y 0.31fF
C1 VPB VPWR 0.20fF
C2 VPWR Y 0.71fF
C3 VPWR VGND 0.21fF
C4 B1 Y 0.47fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__o211a_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__o211a_1 C1 B1 A2 A1 X VGND VPWR VNB VPB
X0 VGND.t0 A1.t0 a_215_47.t0 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 a_510_47.t1 B1.t0 a_215_47.t1 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 a_79_21.t0 C1.t0 VPWR.t1 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 VPWR.t3 B1.t1 a_79_21.t3 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 a_79_21.t2 A2.t0 a_297_297.t1 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 a_297_297.t0 A1.t1 VPWR.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 a_79_21.t1 C1.t1 a_510_47.t0 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 VPWR.t2 a_79_21.t4 X.t0 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 VGND.t1 a_79_21.t5 X.t1 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 a_215_47.t2 A2.t1 VGND.t2 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
R0 A1.n0 A1.t1 241.534
R1 A1.n0 A1.t0 169.234
R2 A1 A1.n0 81.44
R3 a_215_47.t0 a_215_47.n0 188.05
R4 a_215_47.n0 a_215_47.t1 56.307
R5 a_215_47.n0 a_215_47.t2 24.923
R6 VGND.n1 VGND.n0 117.811
R7 VGND.n1 VGND.t1 112.685
R8 VGND.n0 VGND.t0 30.461
R9 VGND.n0 VGND.t2 29.538
R10 VGND VGND.n1 0.208
R11 VNB VNB.t3 6053.91
R12 VNB.t3 VNB.t0 4545.05
R13 VNB.t4 VNB.t2 2852.75
R14 VNB.t2 VNB.t1 2417.58
R15 VNB.t0 VNB.t4 2296.7
R16 B1.n0 B1.t1 239.503
R17 B1.n0 B1.t0 167.203
R18 B1 B1.n0 81.44
R19 a_510_47.t0 a_510_47.t1 64.615
R20 C1.n0 C1.t0 212.079
R21 C1 C1.n0 141.547
R22 C1.n0 C1.t1 139.779
R23 VPWR.n0 VPWR.t0 196.528
R24 VPWR.n2 VPWR.n1 168.689
R25 VPWR.n3 VPWR.t2 159.459
R26 VPWR.n1 VPWR.t1 34.475
R27 VPWR.n1 VPWR.t3 34.475
R28 VPWR.n5 VPWR.n4 4.65
R29 VPWR.n2 VPWR.n0 3.98
R30 VPWR.n4 VPWR.n3 0.752
R31 VPWR.n5 VPWR.n2 0.143
R32 VPWR.n6 VPWR.n5 0.119
R33 VPWR VPWR.n6 0.02
R34 a_79_21.n0 a_79_21.t4 239.546
R35 a_79_21.n2 a_79_21.n0 195.339
R36 a_79_21.n0 a_79_21.t5 167.246
R37 a_79_21.t0 a_79_21.n3 148.51
R38 a_79_21.n3 a_79_21.t1 131.783
R39 a_79_21.n2 a_79_21.n1 107.635
R40 a_79_21.n1 a_79_21.t3 60.085
R41 a_79_21.n3 a_79_21.n2 53.835
R42 a_79_21.n1 a_79_21.t2 26.595
R43 VPB.t3 VPB.t0 556.386
R44 VPB.t2 VPB.t4 349.221
R45 VPB.t4 VPB.t1 295.95
R46 VPB.t0 VPB.t2 281.152
R47 VPB VPB.t3 189.408
R48 A2.n0 A2.t0 233.007
R49 A2.n0 A2.t1 160.707
R50 A2 A2.n0 78.133
R51 a_297_297.t0 a_297_297.t1 64.025
R52 X.n1 X.n0 147.08
R53 X.n2 X.t1 83.131
R54 X.n3 X.n2 62.247
R55 X.n0 X.t0 26.595
R56 X X.n1 10.397
R57 X.n2 X 5.55
R58 X X.n3 4.705
R59 X.n1 X 2.366
C0 X VGND 0.17fF
C1 X VPWR 0.22fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__o211a_2.ext - technology: sky130A

.subckt sky130_fd_sc_hd__o211a_2 C1 B1 A2 A1 X VPWR VGND VNB VPB
X0 a_27_47.t0 B1.t0 VPWR.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 VGND.t2 a_27_47.t4 X.t1 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 VPWR.t4 C1.t0 a_27_47.t2 VPB.t5 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 VPWR.t3 A1.t0 a_373_297.t0 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 a_182_47.t2 A2.t0 VGND.t0 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 X.t3 a_27_47.t5 VPWR.t2 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 a_182_47.t0 B1.t1 a_110_47.t0 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 X.t0 a_27_47.t6 VGND.t1 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 a_373_297.t1 A2.t1 a_27_47.t1 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 a_110_47.t1 C1.t1 a_27_47.t3 VNB.t5 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 VPWR.t1 a_27_47.t7 X.t2 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 VGND.t3 A1.t1 a_182_47.t1 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
R0 B1.n0 B1.t0 235.47
R1 B1.n0 B1.t1 163.17
R2 B1 B1.n0 80.072
R3 VPWR.n2 VPWR.t1 574.869
R4 VPWR.n10 VPWR.n9 163.438
R5 VPWR.n1 VPWR.n0 159.454
R6 VPWR.n0 VPWR.t2 39.4
R7 VPWR.n0 VPWR.t3 37.43
R8 VPWR.n9 VPWR.t0 27.58
R9 VPWR.n9 VPWR.t4 27.58
R10 VPWR.n4 VPWR.n3 4.65
R11 VPWR.n6 VPWR.n5 4.65
R12 VPWR.n8 VPWR.n7 4.65
R13 VPWR.n11 VPWR.n10 3.949
R14 VPWR.n2 VPWR.n1 3.901
R15 VPWR.n4 VPWR.n2 0.261
R16 VPWR.n11 VPWR.n8 0.137
R17 VPWR VPWR.n11 0.122
R18 VPWR.n6 VPWR.n4 0.119
R19 VPWR.n8 VPWR.n6 0.119
R20 a_27_47.n5 a_27_47.t2 258.79
R21 a_27_47.n1 a_27_47.t7 216.652
R22 a_27_47.n2 a_27_47.t5 213.686
R23 a_27_47.n7 a_27_47.n6 146.25
R24 a_27_47.n2 a_27_47.t6 142.745
R25 a_27_47.n1 a_27_47.t4 139.779
R26 a_27_47.n5 a_27_47.t3 137.396
R27 a_27_47.n4 a_27_47.n3 98.594
R28 a_27_47.n7 a_27_47.n0 66.98
R29 a_27_47.t0 a_27_47.n7 41.37
R30 a_27_47.n0 a_27_47.t1 36.445
R31 a_27_47.n3 a_27_47.n2 26.672
R32 a_27_47.n6 a_27_47.n5 22.54
R33 a_27_47.n3 a_27_47.n1 22.341
R34 a_27_47.n6 a_27_47.n4 4.557
R35 VPB.t0 VPB.t1 523.831
R36 VPB.t4 VPB.t3 319.626
R37 VPB.t3 VPB.t2 254.517
R38 VPB.t5 VPB.t0 254.517
R39 VPB.t1 VPB.t4 213.084
R40 VPB VPB.t5 192.367
R41 X X.n0 419.77
R42 X X.n1 75.805
R43 X.n0 X.t2 27.58
R44 X.n0 X.t3 27.58
R45 X.n1 X.t1 25.846
R46 X.n1 X.t0 25.846
R47 VGND.n2 VGND.t2 149.144
R48 VGND.n5 VGND.t0 134.306
R49 VGND.n1 VGND.n0 112.108
R50 VGND.n0 VGND.t1 29.538
R51 VGND.n0 VGND.t3 29.538
R52 VGND.n4 VGND.n3 4.65
R53 VGND.n2 VGND.n1 4.027
R54 VGND.n6 VGND.n5 3.826
R55 VGND VGND.n6 0.355
R56 VGND.n4 VGND.n2 0.225
R57 VGND.n6 VGND.n4 0.143
R58 VNB VNB.t5 6078.09
R59 VNB.t0 VNB.t1 4520.88
R60 VNB.t4 VNB.t2 2272.53
R61 VNB.t2 VNB.t3 2079.12
R62 VNB.t1 VNB.t4 2079.12
R63 VNB.t5 VNB.t0 1740.66
R64 C1.n0 C1.t0 220.365
R65 C1.n0 C1.t1 157.65
R66 C1 C1.n0 80.848
R67 A1.n0 A1.t0 237.733
R68 A1.n0 A1.t1 165.433
R69 A1 A1.n0 85.696
R70 a_373_297.t0 a_373_297.t1 41.37
R71 A2.n0 A2.t1 220.606
R72 A2.n0 A2.t0 160.171
R73 A2 A2.n0 82.012
R74 a_182_47.n1 a_182_47.n0 248.326
R75 a_182_47.n1 a_182_47.t0 77.354
R76 a_182_47.n0 a_182_47.t1 25.846
R77 a_182_47.n0 a_182_47.t2 25.846
R78 a_110_47.t0 a_110_47.t1 38.769
C0 VPWR X 0.21fF
C1 X VGND 0.21fF
C2 A2 A1 0.12fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__o211a_4.ext - technology: sky130A

.subckt sky130_fd_sc_hd__o211a_4 A1 X C1 A2 B1 VGND VPWR VNB VPB
X0 VGND.t7 A1.t0 a_474_47.t5 VNB.t11 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 VPWR.t9 a_79_21.t8 X.t7 VPB.t11 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 VPWR.t4 A1.t1 a_1122_297.t1 VPB.t7 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 X.t6 a_79_21.t9 VPWR.t8 VPB.t10 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 a_79_21.t4 B1.t0 VPWR.t2 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 VGND.t0 a_79_21.t10 X.t3 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 VGND.t1 a_79_21.t11 X.t2 VNB.t5 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 VPWR.t0 C1.t0 a_79_21.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 a_950_297.t1 A1.t2 VPWR.t5 VPB.t6 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 a_557_47.t1 B1.t1 a_474_47.t0 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 a_474_47.t1 B1.t2 a_748_47.t1 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 VGND.t4 A2.t0 a_474_47.t2 VNB.t8 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 VPWR.t7 a_79_21.t12 X.t5 VPB.t9 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13 X.t1 a_79_21.t13 VGND.t2 VNB.t6 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14 a_79_21.t1 C1.t1 a_557_47.t0 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X15 a_474_47.t4 A1.t3 VGND.t6 VNB.t10 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X16 a_79_21.t2 C1.t2 VPWR.t1 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17 a_748_47.t0 C1.t3 a_79_21.t3 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X18 a_474_47.t3 A2.t1 VGND.t5 VNB.t9 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X19 VPWR.t3 B1.t3 a_79_21.t5 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X20 a_79_21.t6 A2.t2 a_950_297.t0 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X21 a_1122_297.t0 A2.t3 a_79_21.t7 VPB.t5 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X22 X.t4 a_79_21.t14 VPWR.t6 VPB.t8 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X23 X.t0 a_79_21.t15 VGND.t3 VNB.t7 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
R0 A1.n0 A1.t2 236.179
R1 A1.n1 A1.t1 231.961
R2 A1 A1.n0 166.544
R3 A1.n0 A1.t0 163.879
R4 A1.n1 A1.t3 159.661
R5 A1 A1.n1 85.12
R6 a_474_47.t0 a_474_47.n3 284.586
R7 a_474_47.n1 a_474_47.t4 129.919
R8 a_474_47.n3 a_474_47.n1 56.247
R9 a_474_47.n1 a_474_47.n0 52.431
R10 a_474_47.n3 a_474_47.n2 43.173
R11 a_474_47.n2 a_474_47.t1 30.461
R12 a_474_47.n2 a_474_47.t5 28.615
R13 a_474_47.n0 a_474_47.t2 25.846
R14 a_474_47.n0 a_474_47.t3 25.846
R15 VGND.n23 VGND.t3 190.315
R16 VGND.n14 VGND.t1 179.046
R17 VGND.n3 VGND.n0 120.465
R18 VGND.n2 VGND.n1 107.128
R19 VGND.n19 VGND.n18 106.463
R20 VGND.n1 VGND.t5 38.769
R21 VGND.n1 VGND.t7 33.23
R22 VGND.n0 VGND.t6 25.846
R23 VGND.n0 VGND.t4 25.846
R24 VGND.n18 VGND.t2 24.923
R25 VGND.n18 VGND.t0 24.923
R26 VGND.n24 VGND.n23 4.65
R27 VGND.n5 VGND.n4 4.65
R28 VGND.n7 VGND.n6 4.65
R29 VGND.n9 VGND.n8 4.65
R30 VGND.n11 VGND.n10 4.65
R31 VGND.n13 VGND.n12 4.65
R32 VGND.n15 VGND.n14 4.65
R33 VGND.n17 VGND.n16 4.65
R34 VGND.n20 VGND.n19 4.65
R35 VGND.n22 VGND.n21 4.65
R36 VGND.n3 VGND.n2 3.874
R37 VGND.n5 VGND.n3 0.215
R38 VGND.n7 VGND.n5 0.119
R39 VGND.n9 VGND.n7 0.119
R40 VGND.n11 VGND.n9 0.119
R41 VGND.n13 VGND.n11 0.119
R42 VGND.n15 VGND.n13 0.119
R43 VGND.n17 VGND.n15 0.119
R44 VGND.n20 VGND.n17 0.119
R45 VGND.n22 VGND.n20 0.119
R46 VGND.n24 VGND.n22 0.119
R47 VGND VGND.n24 0.022
R48 VNB VNB.t7 6078.09
R49 VNB.t5 VNB.t2 4738.46
R50 VNB.t0 VNB.t1 2876.92
R51 VNB.t11 VNB.t9 2610.99
R52 VNB.t3 VNB.t11 2272.53
R53 VNB.t8 VNB.t10 2079.12
R54 VNB.t9 VNB.t8 2079.12
R55 VNB.t1 VNB.t3 2079.12
R56 VNB.t6 VNB.t5 2030.77
R57 VNB.t4 VNB.t6 2030.77
R58 VNB.t7 VNB.t4 2030.77
R59 VNB.t2 VNB.t0 1740.66
R60 a_79_21.n2 a_79_21.n1 306.255
R61 a_79_21.n20 a_79_21.n19 292.5
R62 a_79_21.n2 a_79_21.n0 230.507
R63 a_79_21.n16 a_79_21.t8 225.224
R64 a_79_21.n14 a_79_21.t14 212.079
R65 a_79_21.n9 a_79_21.t12 212.079
R66 a_79_21.n5 a_79_21.t9 212.079
R67 a_79_21.n18 a_79_21.n3 187.411
R68 a_79_21.n4 a_79_21.t15 173.372
R69 a_79_21.n6 a_79_21.t10 139.779
R70 a_79_21.n10 a_79_21.t13 139.779
R71 a_79_21.n13 a_79_21.t11 139.779
R72 a_79_21.n8 a_79_21.n4 97.76
R73 a_79_21.n19 a_79_21.n18 79.761
R74 a_79_21.n15 a_79_21.n14 76
R75 a_79_21.n12 a_79_21.n11 76
R76 a_79_21.n8 a_79_21.n7 76
R77 a_79_21.n17 a_79_21.n16 76
R78 a_79_21.n19 a_79_21.n2 58.05
R79 a_79_21.t0 a_79_21.n20 52.205
R80 a_79_21.n20 a_79_21.t4 47.28
R81 a_79_21.n3 a_79_21.t3 43.384
R82 a_79_21.n1 a_79_21.t2 41.37
R83 a_79_21.n3 a_79_21.t1 38.769
R84 a_79_21.n1 a_79_21.t5 35.46
R85 a_79_21.n0 a_79_21.t7 27.58
R86 a_79_21.n0 a_79_21.t6 27.58
R87 a_79_21.n7 a_79_21.n6 21.909
R88 a_79_21.n17 a_79_21.n15 21.76
R89 a_79_21.n15 a_79_21.n12 21.76
R90 a_79_21.n12 a_79_21.n8 21.76
R91 a_79_21.n18 a_79_21.n17 14.4
R92 a_79_21.n11 a_79_21.n10 10.224
R93 a_79_21.n6 a_79_21.n5 4.381
R94 a_79_21.n10 a_79_21.n9 2.921
R95 a_79_21.n14 a_79_21.n13 1.46
R96 X.n2 X.n1 205.081
R97 X.n2 X.n0 164.227
R98 X.n5 X.n4 163.771
R99 X.n5 X.n3 107.182
R100 X X.n2 70.623
R101 X.n1 X.t7 27.58
R102 X.n1 X.t4 27.58
R103 X.n0 X.t5 27.58
R104 X.n0 X.t6 27.58
R105 X X.n5 25.1
R106 X.n3 X.t3 24.923
R107 X.n3 X.t0 24.923
R108 X.n4 X.t2 24.923
R109 X.n4 X.t1 24.923
R110 VPWR.n1 VPWR.n0 309.888
R111 VPWR.n11 VPWR.n10 308.015
R112 VPWR.n6 VPWR.n5 306.463
R113 VPWR.n2 VPWR.t4 196.11
R114 VPWR.n20 VPWR.t8 192.21
R115 VPWR.n16 VPWR.n15 164.63
R116 VPWR.n0 VPWR.t5 35.46
R117 VPWR.n0 VPWR.t3 27.58
R118 VPWR.n5 VPWR.t1 27.58
R119 VPWR.n5 VPWR.t0 27.58
R120 VPWR.n10 VPWR.t2 27.58
R121 VPWR.n10 VPWR.t9 27.58
R122 VPWR.n15 VPWR.t6 27.58
R123 VPWR.n15 VPWR.t7 27.58
R124 VPWR.n4 VPWR.n3 4.65
R125 VPWR.n7 VPWR.n6 4.65
R126 VPWR.n9 VPWR.n8 4.65
R127 VPWR.n12 VPWR.n11 4.65
R128 VPWR.n14 VPWR.n13 4.65
R129 VPWR.n17 VPWR.n16 4.65
R130 VPWR.n19 VPWR.n18 4.65
R131 VPWR.n2 VPWR.n1 3.898
R132 VPWR.n21 VPWR.n20 3.865
R133 VPWR.n4 VPWR.n2 0.142
R134 VPWR.n21 VPWR.n19 0.139
R135 VPWR VPWR.n21 0.121
R136 VPWR.n7 VPWR.n4 0.119
R137 VPWR.n9 VPWR.n7 0.119
R138 VPWR.n12 VPWR.n9 0.119
R139 VPWR.n14 VPWR.n12 0.119
R140 VPWR.n17 VPWR.n14 0.119
R141 VPWR.n19 VPWR.n17 0.119
R142 VPB VPB.t10 423.208
R143 VPB.t2 VPB.t0 387.694
R144 VPB.t1 VPB.t3 319.626
R145 VPB.t3 VPB.t6 278.193
R146 VPB.t5 VPB.t7 254.517
R147 VPB.t4 VPB.t5 254.517
R148 VPB.t6 VPB.t4 254.517
R149 VPB.t0 VPB.t1 254.517
R150 VPB.t11 VPB.t2 254.517
R151 VPB.t8 VPB.t11 254.517
R152 VPB.t9 VPB.t8 254.517
R153 VPB.t10 VPB.t9 254.517
R154 a_1122_297.t0 a_1122_297.t1 55.16
R155 B1.n0 B1.t0 239.038
R156 B1.n1 B1.t3 236.179
R157 B1.n0 B1.t1 166.738
R158 B1.n1 B1.t2 163.879
R159 B1 B1.n0 146.675
R160 B1 B1.n1 87.054
R161 C1.n1 C1.t0 212.079
R162 C1.n0 C1.t2 212.079
R163 C1.n1 C1.t1 163.879
R164 C1.n0 C1.t3 139.779
R165 C1.n2 C1.n0 32.908
R166 C1 C1.n2 32.897
R167 C1.n2 C1.n1 18.678
R168 a_950_297.t0 a_950_297.t1 55.16
R169 a_557_47.t0 a_557_47.t1 38.769
R170 a_748_47.t0 a_748_47.t1 51.692
R171 A2.n0 A2.t3 212.079
R172 A2.n1 A2.t2 212.079
R173 A2.n0 A2.t0 139.779
R174 A2.n1 A2.t1 139.779
R175 A2 A2.n2 31.938
R176 A2.n2 A2.n1 30.615
R177 A2.n2 A2.n0 20.809
C0 A1 A2 0.38fF
C1 B1 A1 0.14fF
C2 VPWR X 0.49fF
C3 VPWR VGND 0.14fF
C4 B1 C1 0.35fF
C5 X VGND 0.33fF
C6 VPB VPWR 0.13fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__o211ai_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__o211ai_1 A1 A2 Y C1 B1 VGND VPWR VNB VPB
X0 a_110_297.t0 A1.t0 VPWR.t1 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 VGND.t0 A1.t1 a_27_47.t0 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 Y.t1 A2.t0 a_110_297.t1 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 VPWR.t0 B1.t0 Y.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 a_27_47.t1 A2.t1 VGND.t1 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 a_326_47.t0 B1.t1 a_27_47.t2 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 Y.t3 C1.t0 VPWR.t2 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 Y.t2 C1.t1 a_326_47.t1 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
R0 A1.n0 A1.t0 233.287
R1 A1.n0 A1.t1 160.987
R2 A1 A1.n0 82.4
R3 VPWR.n1 VPWR.n0 310.197
R4 VPWR.n1 VPWR.t1 150.721
R5 VPWR.n0 VPWR.t2 45.31
R6 VPWR.n0 VPWR.t0 31.52
R7 VPWR VPWR.n1 0.054
R8 a_110_297.t0 a_110_297.t1 41.37
R9 VPB.t0 VPB.t2 319.626
R10 VPB.t3 VPB.t0 319.626
R11 VPB.t1 VPB.t3 213.084
R12 VPB VPB.t1 195.327
R13 a_27_47.t0 a_27_47.n0 179.681
R14 a_27_47.n0 a_27_47.t1 36.923
R15 a_27_47.n0 a_27_47.t2 35.076
R16 VGND VGND.n0 109.991
R17 VGND.n0 VGND.t0 38.769
R18 VGND.n0 VGND.t1 33.23
R19 VNB VNB.t0 6102.26
R20 VNB.t2 VNB.t3 2610.99
R21 VNB.t0 VNB.t2 2610.99
R22 VNB.t3 VNB.t1 1740.66
R23 A2.n0 A2.t0 236.179
R24 A2.n0 A2.t1 163.879
R25 A2 A2.n0 92.986
R26 Y.n1 Y.n0 147.111
R27 Y.n2 Y.n1 71.003
R28 Y.n1 Y.t3 63.04
R29 Y.n2 Y.t2 57.23
R30 Y.n0 Y.t1 39.4
R31 Y.n0 Y.t0 37.43
R32 Y Y.n2 2.253
R33 B1.n0 B1.t0 230.92
R34 B1.n0 B1.t1 163.879
R35 B1.n1 B1.n0 76
R36  B1.n1 8.992
R37 B1.n1 B1 1.422
R38 a_326_47.t0 a_326_47.t1 38.769
R39 C1.n0 C1.t0 230.574
R40 C1.n0 C1.t1 158.274
R41 C1 C1.n0 87.054
C0 A1 A2 0.11fF
C1 Y VGND 0.13fF
C2 C1 Y 0.19fF
C3 B1 C1 0.12fF
C4 VPWR Y 0.32fF
C5 A2 Y 0.11fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__o211ai_2.ext - technology: sky130A

.subckt sky130_fd_sc_hd__o211ai_2 A1 A2 B1 Y C1 VGND VPWR VNB VPB
X0 a_286_47.t3 A1.t0 VGND.t1 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 VPWR.t1 B1.t0 Y.t1 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 a_286_47.t4 A2.t0 VGND.t2 VNB.t6 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 Y.t6 A2.t1 a_487_297.t1 VPB.t6 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 VGND.t0 A1.t1 a_286_47.t2 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 Y.t2 C1.t0 a_27_47.t1 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 VGND.t3 A2.t2 a_286_47.t5 VNB.t7 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 a_487_297.t0 A2.t3 Y.t7 VPB.t7 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 a_27_47.t3 B1.t1 a_286_47.t0 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 VPWR.t4 C1.t1 Y.t3 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 VPWR.t3 A1.t2 a_487_297.t3 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 a_27_47.t0 C1.t2 Y.t4 VNB.t5 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 Y.t5 C1.t3 VPWR.t5 VPB.t5 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13 a_487_297.t2 A1.t3 VPWR.t2 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14 a_286_47.t1 B1.t2 a_27_47.t2 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X15 Y.t0 B1.t3 VPWR.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
R0 A1.n0 A1.t3 212.079
R1 A1.n1 A1.t2 212.079
R2 A1.n0 A1.t1 139.779
R3 A1.n1 A1.t0 139.779
R4 A1 A1.n2 54.793
R5 A1.n2 A1.n1 26.592
R6 A1.n2 A1.n0 25.077
R7 VGND.n2 VGND.t0 194.475
R8 VGND.n5 VGND.t2 190.673
R9 VGND.n1 VGND.n0 106.463
R10 VGND.n0 VGND.t1 25.846
R11 VGND.n0 VGND.t3 25.846
R12 VGND.n4 VGND.n3 4.65
R13 VGND.n6 VGND.n5 3.984
R14 VGND.n2 VGND.n1 3.853
R15 VGND VGND.n6 0.601
R16 VGND.n4 VGND.n2 0.262
R17 VGND.n6 VGND.n4 0.138
R18 a_286_47.n2 a_286_47.n1 179.052
R19 a_286_47.n3 a_286_47.n2 144.919
R20 a_286_47.n2 a_286_47.n0 92.5
R21 a_286_47.n1 a_286_47.t0 25.846
R22 a_286_47.n1 a_286_47.t1 25.846
R23 a_286_47.n0 a_286_47.t5 25.846
R24 a_286_47.n0 a_286_47.t4 25.846
R25 a_286_47.n3 a_286_47.t2 25.846
R26 a_286_47.t3 a_286_47.n3 25.846
R27 VNB VNB.t4 6198.96
R28 VNB.t0 VNB.t6 4786.81
R29 VNB.t3 VNB.t2 2079.12
R30 VNB.t7 VNB.t3 2079.12
R31 VNB.t6 VNB.t7 2079.12
R32 VNB.t1 VNB.t0 2079.12
R33 VNB.t5 VNB.t1 2079.12
R34 VNB.t4 VNB.t5 2079.12
R35 B1.n0 B1.t0 212.079
R36 B1.n1 B1.t3 212.079
R37 B1.n0 B1.t1 139.779
R38 B1.n1 B1.t2 139.779
R39 B1.n2 B1.n0 33.085
R40 B1 B1.n2 32.741
R41 B1.n2 B1.n1 19
R42 Y.n2 Y.n0 239.725
R43 Y.n2 Y.n1 168.353
R44 Y.n4 Y.n3 160.64
R45 Y Y.n5 92.693
R46 Y.n4 Y.n2 45.176
R47 Y Y.n4 33.357
R48 Y.n0 Y.t7 27.58
R49 Y.n0 Y.t6 27.58
R50 Y.n1 Y.t1 27.58
R51 Y.n1 Y.t0 27.58
R52 Y.n3 Y.t3 27.58
R53 Y.n3 Y.t5 27.58
R54 Y.n5 Y.t4 25.846
R55 Y.n5 Y.t2 25.846
R56 VPWR.n10 VPWR.t5 575.112
R57 VPWR.n1 VPWR.t1 191.794
R58 VPWR.n2 VPWR.n0 168.517
R59 VPWR.n6 VPWR.n5 164.214
R60 VPWR.n5 VPWR.t0 27.58
R61 VPWR.n5 VPWR.t4 27.58
R62 VPWR.n0 VPWR.t2 27.58
R63 VPWR.n0 VPWR.t3 27.58
R64 VPWR.n4 VPWR.n3 4.65
R65 VPWR.n7 VPWR.n6 4.65
R66 VPWR.n9 VPWR.n8 4.65
R67 VPWR.n11 VPWR.n10 4.65
R68 VPWR.n2 VPWR.n1 4.038
R69 VPWR.n4 VPWR.n2 0.138
R70 VPWR.n7 VPWR.n4 0.119
R71 VPWR.n9 VPWR.n7 0.119
R72 VPWR.n11 VPWR.n9 0.119
R73 VPWR VPWR.n11 0.022
R74 VPB.t1 VPB.t6 585.981
R75 VPB.t3 VPB.t2 254.517
R76 VPB.t7 VPB.t3 254.517
R77 VPB.t6 VPB.t7 254.517
R78 VPB.t0 VPB.t1 254.517
R79 VPB.t4 VPB.t0 254.517
R80 VPB.t5 VPB.t4 254.517
R81 VPB VPB.t5 207.165
R82 A2.n0 A2.t3 212.079
R83 A2.n1 A2.t1 212.079
R84 A2.n0 A2.t2 139.779
R85 A2.n1 A2.t0 139.779
R86 A2 A2.n2 49.632
R87 A2.n2 A2.n0 26.043
R88 A2.n2 A2.n1 25.41
R89 a_487_297.t1 a_487_297.n1 601.007
R90 a_487_297.n1 a_487_297.t2 275.231
R91 a_487_297.n1 a_487_297.n0 138.665
R92 a_487_297.n0 a_487_297.t3 27.58
R93 a_487_297.n0 a_487_297.t0 27.58
R94 C1.n0 C1.t1 212.079
R95 C1.n1 C1.t3 212.079
R96 C1.n0 C1.t2 139.779
R97 C1.n1 C1.t0 139.779
R98 C1 C1.n1 125.824
R99 C1.n1 C1.n0 62.806
R100 a_27_47.t1 a_27_47.n1 234.036
R101 a_27_47.n1 a_27_47.t3 229.129
R102 a_27_47.n1 a_27_47.n0 49.967
R103 a_27_47.n0 a_27_47.t2 25.846
R104 a_27_47.n0 a_27_47.t0 25.846
C0 A2 Y 0.13fF
C1 VPWR Y 0.48fF
C2 VPWR VGND 0.10fF
C3 C1 Y 0.14fF
C4 B1 Y 0.26fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__o211ai_4.ext - technology: sky130A

.subckt sky130_fd_sc_hd__o211ai_4 A1 B1 A2 C1 Y VGND VPWR VNB VPB
X0 VPWR.t11 A1.t0 a_110_297.t3 VPB.t11 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 Y.t15 A2.t0 a_110_297.t4 VPB.t12 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 a_806_47.t3 B1.t0 a_27_47.t5 VNB.t11 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 a_110_297.t5 A2.t1 Y.t14 VPB.t13 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 a_110_297.t2 A1.t1 VPWR.t10 VPB.t10 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 VGND.t7 A1.t2 a_27_47.t11 VNB.t15 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 VPWR.t2 B1.t1 Y.t2 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 a_110_297.t1 A1.t3 VPWR.t9 VPB.t9 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 a_27_47.t3 A2.t2 VGND.t3 VNB.t7 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 VPWR.t8 A1.t4 a_110_297.t0 VPB.t8 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 VPWR.t4 C1.t0 Y.t4 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 a_27_47.t7 B1.t2 a_1314_47.t0 VNB.t10 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 Y.t5 C1.t1 VPWR.t5 VPB.t5 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13 a_27_47.t10 A1.t5 VGND.t6 VNB.t14 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14 VPWR.t6 C1.t2 Y.t6 VPB.t6 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 Y.t3 B1.t3 VPWR.t3 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16 VGND.t5 A1.t6 a_27_47.t9 VNB.t13 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X17 Y.t13 A2.t3 a_110_297.t6 VPB.t14 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X18 a_27_47.t8 A1.t7 VGND.t4 VNB.t12 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X19 Y.t7 C1.t3 a_978_47.t1 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X20 Y.t8 C1.t4 a_806_47.t0 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X21 a_27_47.t2 A2.t4 VGND.t2 VNB.t6 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X22 a_27_47.t6 B1.t4 a_806_47.t2 VNB.t9 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X23 a_110_297.t7 A2.t5 Y.t12 VPB.t15 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X24 a_806_47.t1 C1.t5 Y.t9 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X25 VPWR.t0 B1.t5 Y.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X26 VGND.t1 A2.t6 a_27_47.t1 VNB.t5 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X27 a_978_47.t0 B1.t6 a_27_47.t4 VNB.t8 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X28 a_1314_47.t1 C1.t6 Y.t10 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X29 Y.t11 C1.t7 VPWR.t7 VPB.t7 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X30 Y.t1 B1.t7 VPWR.t1 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X31 VGND.t0 A2.t7 a_27_47.t0 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
R0 A1.n3 A1.n0 245.646
R1 A1.n0 A1.t4 236.179
R2 A1.n4 A1.t0 212.079
R3 A1.n1 A1.t3 212.079
R4 A1.n5 A1.t1 212.079
R5 A1.n0 A1.t7 163.879
R6 A1.n4 A1.t5 139.779
R7 A1.n1 A1.t2 139.779
R8 A1.n5 A1.t6 139.779
R9 A1.n3 A1.n2 76
R10 A1 A1.n6 37.552
R11 A1.n6 A1.n5 34.275
R12 A1.n6 A1.n4 17.256
R13 A1.n2 A1.n1 13.145
R14 A1 A1.n3 3.672
R15 a_110_297.n3 a_110_297.n2 356.951
R16 a_110_297.n5 a_110_297.n4 350.436
R17 a_110_297.n3 a_110_297.n1 292.5
R18 a_110_297.n4 a_110_297.n0 292.5
R19 a_110_297.n4 a_110_297.n3 66.45
R20 a_110_297.n0 a_110_297.t4 27.58
R21 a_110_297.n0 a_110_297.t7 27.58
R22 a_110_297.n1 a_110_297.t6 27.58
R23 a_110_297.n1 a_110_297.t1 27.58
R24 a_110_297.n2 a_110_297.t3 27.58
R25 a_110_297.n2 a_110_297.t2 27.58
R26 a_110_297.t0 a_110_297.n5 27.58
R27 a_110_297.n5 a_110_297.t5 27.58
R28 VPWR.n2 VPWR.t0 414.956
R29 VPWR.n15 VPWR.n14 309.566
R30 VPWR.n29 VPWR.n28 306.463
R31 VPWR.n11 VPWR.n10 306.463
R32 VPWR.n6 VPWR.n5 306.463
R33 VPWR.n1 VPWR.n0 306.255
R34 VPWR.n33 VPWR.t10 258.994
R35 VPWR.n14 VPWR.t1 31.52
R36 VPWR.n14 VPWR.t8 31.52
R37 VPWR.n28 VPWR.t9 27.58
R38 VPWR.n28 VPWR.t11 27.58
R39 VPWR.n10 VPWR.t3 27.58
R40 VPWR.n10 VPWR.t2 27.58
R41 VPWR.n5 VPWR.t5 26.595
R42 VPWR.n5 VPWR.t6 26.595
R43 VPWR.n0 VPWR.t7 26.595
R44 VPWR.n0 VPWR.t4 26.595
R45 VPWR.n12 VPWR.n11 4.894
R46 VPWR.n4 VPWR.n3 4.65
R47 VPWR.n7 VPWR.n6 4.65
R48 VPWR.n9 VPWR.n8 4.65
R49 VPWR.n13 VPWR.n12 4.65
R50 VPWR.n17 VPWR.n16 4.65
R51 VPWR.n19 VPWR.n18 4.65
R52 VPWR.n21 VPWR.n20 4.65
R53 VPWR.n23 VPWR.n22 4.65
R54 VPWR.n25 VPWR.n24 4.65
R55 VPWR.n27 VPWR.n26 4.65
R56 VPWR.n30 VPWR.n29 4.65
R57 VPWR.n32 VPWR.n31 4.65
R58 VPWR.n34 VPWR.n33 4.65
R59 VPWR.n2 VPWR.n1 3.748
R60 VPWR.n16 VPWR.n15 1.882
R61 VPWR.n4 VPWR.n2 0.161
R62 VPWR.n7 VPWR.n4 0.119
R63 VPWR.n9 VPWR.n7 0.119
R64 VPWR.n13 VPWR.n9 0.119
R65 VPWR.n17 VPWR.n13 0.119
R66 VPWR.n19 VPWR.n17 0.119
R67 VPWR.n21 VPWR.n19 0.119
R68 VPWR.n23 VPWR.n21 0.119
R69 VPWR.n25 VPWR.n23 0.119
R70 VPWR.n27 VPWR.n25 0.119
R71 VPWR.n30 VPWR.n27 0.119
R72 VPWR.n32 VPWR.n30 0.119
R73 VPWR.n34 VPWR.n32 0.119
R74 VPWR VPWR.n34 0.02
R75 VPB.t8 VPB.t1 278.193
R76 VPB.t2 VPB.t3 254.517
R77 VPB.t1 VPB.t2 254.517
R78 VPB.t13 VPB.t8 254.517
R79 VPB.t12 VPB.t13 254.517
R80 VPB.t15 VPB.t12 254.517
R81 VPB.t14 VPB.t15 254.517
R82 VPB.t9 VPB.t14 254.517
R83 VPB.t11 VPB.t9 254.517
R84 VPB.t10 VPB.t11 254.517
R85 VPB.t7 VPB.t0 248.598
R86 VPB.t4 VPB.t7 248.598
R87 VPB.t5 VPB.t4 248.598
R88 VPB.t6 VPB.t5 248.598
R89 VPB.t3 VPB.t6 248.598
R90 VPB VPB.t10 192.367
R91 A2.n0 A2.t1 196.012
R92 A2.n2 A2.t0 196.012
R93 A2.n5 A2.t5 196.012
R94 A2.n8 A2.t3 196.012
R95 A2.n0 A2.t6 139.779
R96 A2.n2 A2.t4 139.779
R97 A2.n5 A2.t7 139.779
R98 A2.n8 A2.t2 139.779
R99 A2.n4 A2.n1 92.118
R100 A2 A2.n9 81.688
R101 A2.n4 A2.n3 76
R102 A2.n7 A2.n6 76
R103 A2.n1 A2.n0 20.928
R104 A2.n7 A2.n4 16.118
R105 A2.n9 A2.n8 13.318
R106 A2 A2.n7 10.429
R107 A2.n3 A2.n2 9.513
R108 A2.n6 A2.n5 1.902
R109 Y.n6 Y.n5 336.532
R110 Y.n6 Y.n4 292.5
R111 Y.n10 Y.n0 292.5
R112 Y.n9 Y.n1 292.5
R113 Y.n8 Y.n2 292.5
R114 Y.n7 Y.n3 292.5
R115 Y.n13 Y.n12 152.233
R116 Y Y.n13 134.376
R117 Y.n13 Y.n11 92.5
R118 Y.n7 Y.n6 81.95
R119 Y.n8 Y.n7 43.776
R120 Y.n10 Y.n9 43.008
R121 Y.n9 Y.n8 43.008
R122 Y Y.n10 28.702
R123 Y.n3 Y.t2 27.58
R124 Y.n3 Y.t1 27.58
R125 Y.n5 Y.t12 27.58
R126 Y.n5 Y.t13 27.58
R127 Y.n4 Y.t14 27.58
R128 Y.n4 Y.t15 27.58
R129 Y.n2 Y.t6 26.595
R130 Y.n2 Y.t3 26.595
R131 Y.n1 Y.t4 26.595
R132 Y.n1 Y.t5 26.595
R133 Y.n0 Y.t0 26.595
R134 Y.n0 Y.t11 26.595
R135 Y.n12 Y.t9 24.923
R136 Y.n12 Y.t7 24.923
R137 Y.n11 Y.t10 24.923
R138 Y.n11 Y.t8 24.923
R139 B1 B1.n0 252.972
R140 B1.n0 B1.t5 241.534
R141 B1.n2 B1.t1 212.079
R142 B1.n4 B1.t3 212.079
R143 B1.n1 B1.t7 212.079
R144 B1.n0 B1.t2 169.234
R145 B1.n2 B1.t4 139.779
R146 B1.n4 B1.t6 139.779
R147 B1.n1 B1.t0 139.779
R148 B1.n6 B1.n5 76
R149 B1.n6 B1.n3 36.962
R150 B1.n3 B1.n1 33.176
R151 B1.n3 B1.n2 17.921
R152 B1.n5 B1.n4 13.145
R153 B1 B1.n6 0.463
R154 a_27_47.n7 a_27_47.t7 197.924
R155 a_27_47.n6 a_27_47.t9 157.66
R156 a_27_47.n2 a_27_47.n1 149.251
R157 a_27_47.n6 a_27_47.n5 92.5
R158 a_27_47.n2 a_27_47.n0 92.5
R159 a_27_47.n4 a_27_47.n3 92.5
R160 a_27_47.n9 a_27_47.n8 92.5
R161 a_27_47.n8 a_27_47.n7 82.703
R162 a_27_47.n4 a_27_47.n2 63.195
R163 a_27_47.n8 a_27_47.n4 45.866
R164 a_27_47.n0 a_27_47.t5 29.538
R165 a_27_47.n0 a_27_47.t8 27.692
R166 a_27_47.n3 a_27_47.t1 25.846
R167 a_27_47.n3 a_27_47.t2 25.846
R168 a_27_47.n5 a_27_47.t11 25.846
R169 a_27_47.n5 a_27_47.t10 25.846
R170 a_27_47.n1 a_27_47.t4 25.846
R171 a_27_47.n1 a_27_47.t6 25.846
R172 a_27_47.t0 a_27_47.n9 25.846
R173 a_27_47.n9 a_27_47.t3 25.846
R174 a_27_47.n7 a_27_47.n6 0.457
R175 a_806_47.n1 a_806_47.n0 305.533
R176 a_806_47.t2 a_806_47.n1 25.846
R177 a_806_47.n1 a_806_47.t3 25.846
R178 a_806_47.n0 a_806_47.t0 24.923
R179 a_806_47.n0 a_806_47.t1 24.923
R180 VNB VNB.t13 6078.09
R181 VNB.t3 VNB.t10 2272.53
R182 VNB.t12 VNB.t11 2224.18
R183 VNB.t5 VNB.t12 2127.47
R184 VNB.t9 VNB.t8 2079.12
R185 VNB.t11 VNB.t9 2079.12
R186 VNB.t6 VNB.t5 2079.12
R187 VNB.t4 VNB.t6 2079.12
R188 VNB.t7 VNB.t4 2079.12
R189 VNB.t15 VNB.t7 2079.12
R190 VNB.t14 VNB.t15 2079.12
R191 VNB.t13 VNB.t14 2079.12
R192 VNB.t1 VNB.t3 2030.77
R193 VNB.t2 VNB.t1 2030.77
R194 VNB.t0 VNB.t2 2030.77
R195 VNB.t8 VNB.t0 2030.77
R196 VGND.n7 VGND.n6 113.205
R197 VGND.n3 VGND.n2 110.2
R198 VGND.n1 VGND.n0 106.463
R199 VGND.n13 VGND.n12 106.463
R200 VGND.n2 VGND.t4 27.692
R201 VGND.n2 VGND.t1 25.846
R202 VGND.n0 VGND.t2 25.846
R203 VGND.n0 VGND.t0 25.846
R204 VGND.n6 VGND.t3 25.846
R205 VGND.n6 VGND.t7 25.846
R206 VGND.n12 VGND.t6 25.846
R207 VGND.n12 VGND.t5 25.846
R208 VGND.n5 VGND.n4 4.65
R209 VGND.n9 VGND.n8 4.65
R210 VGND.n11 VGND.n10 4.65
R211 VGND.n8 VGND.n7 4.517
R212 VGND.n14 VGND.n13 3.949
R213 VGND.n3 VGND.n1 3.931
R214 VGND.n5 VGND.n3 0.292
R215 VGND.n14 VGND.n11 0.137
R216 VGND VGND.n14 0.122
R217 VGND.n9 VGND.n5 0.119
R218 VGND.n11 VGND.n9 0.119
R219 C1.n0 C1.t7 212.079
R220 C1.n5 C1.t0 212.079
R221 C1.n2 C1.t1 212.079
R222 C1.n3 C1.t2 212.079
R223 C1.n0 C1.t6 139.779
R224 C1.n5 C1.t4 139.779
R225 C1.n2 C1.t5 139.779
R226 C1.n3 C1.t3 139.779
R227 C1.n7 C1.n4 92.118
R228 C1 C1.n1 82.874
R229 C1.n7 C1.n6 76
R230 C1.n4 C1.n3 52.581
R231 C1.n1 C1.n0 32.133
R232 C1.n6 C1.n5 20.448
R233 C1 C1.n7 9.244
R234 C1.n4 C1.n2 8.763
R235 a_1314_47.t0 a_1314_47.t1 59.076
R236 a_978_47.t0 a_978_47.t1 49.846
C0 B1 Y 0.65fF
C1 A1 A2 0.56fF
C2 Y VGND 0.25fF
C3 B1 C1 0.43fF
C4 A1 Y 0.31fF
C5 A1 B1 0.14fF
C6 VPWR Y 0.52fF
C7 VPB VPWR 0.16fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__o221a_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__o221a_1 A2 X B1 C1 A1 B2 VGND VPWR VNB VPB
X0 a_240_47.t3 A2.t0 VGND.t2 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 X.t1 a_51_297.t4 VGND.t0 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 VGND.t1 A1.t0 a_240_47.t1 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 a_51_297.t0 B2.t0 a_245_297.t1 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 a_149_47.t2 C1.t0 a_51_297.t2 VNB.t5 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 a_240_47.t0 B1.t0 a_149_47.t0 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 VPWR.t1 A1.t1 a_512_297.t0 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 X.t0 a_51_297.t5 VPWR.t2 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 a_149_47.t1 B2.t1 a_240_47.t2 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 a_245_297.t0 B1.t1 VPWR.t3 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 VPWR.t0 C1.t1 a_51_297.t3 VPB.t5 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 a_512_297.t1 A2.t1 a_51_297.t1 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
R0 A2.n0 A2.t1 233.573
R1 A2.n0 A2.t0 161.273
R2 A2 A2.n0 82.501
R3 VGND.n1 VGND.t2 204.383
R4 VGND.n1 VGND.n0 84.145
R5 VGND.n0 VGND.t0 24.923
R6 VGND.n0 VGND.t1 24.923
R7 VGND VGND.n1 0.706
R8 a_240_47.n1 a_240_47.n0 229.82
R9 a_240_47.n0 a_240_47.t1 24.923
R10 a_240_47.n0 a_240_47.t3 24.923
R11 a_240_47.n1 a_240_47.t2 24.923
R12 a_240_47.t0 a_240_47.n1 24.923
R13 VNB VNB.t5 7053.3
R14 VNB.t3 VNB.t4 4545.05
R15 VNB.t5 VNB.t0 2200
R16 VNB.t2 VNB.t1 2030.77
R17 VNB.t4 VNB.t2 2030.77
R18 VNB.t0 VNB.t3 2030.77
R19 a_51_297.n1 a_51_297.t5 234.481
R20 a_51_297.n2 a_51_297.n1 190.346
R21 a_51_297.n1 a_51_297.t4 162.181
R22 a_51_297.n5 a_51_297.n4 146.25
R23 a_51_297.n3 a_51_297.t3 145.986
R24 a_51_297.n3 a_51_297.t2 137.864
R25 a_51_297.n5 a_51_297.n0 109.335
R26 a_51_297.n4 a_51_297.n3 90.108
R27 a_51_297.n0 a_51_297.t1 26.595
R28 a_51_297.t0 a_51_297.n5 26.595
R29 a_51_297.n4 a_51_297.n2 12.04
R30 X.n0 X.t0 180.04
R31 X X.t1 132.564
R32 X.n0 X 4.608
R33 X X.n0 1.732
R34 A1.n0 A1.t1 241.534
R35 A1.n0 A1.t0 169.234
R36 A1 A1.n0 77.564
R37 B2.n0 B2.t0 234.801
R38 B2.n0 B2.t1 162.501
R39 B2.n1 B2.n0 76
R40 B2 B2.n1 11.4
R41 B2.n1 B2 2.2
R42 a_245_297.t0 a_245_297.t1 41.37
R43 VPB.t1 VPB.t4 577.102
R44 VPB VPB.t5 310.747
R45 VPB.t2 VPB.t3 284.112
R46 VPB.t5 VPB.t0 284.112
R47 VPB.t4 VPB.t2 213.084
R48 VPB.t0 VPB.t1 213.084
R49 C1.n0 C1.t1 212.079
R50 C1 C1.n0 141.979
R51 C1.n0 C1.t0 139.779
R52 a_149_47.n0 a_149_47.t1 327.084
R53 a_149_47.n0 a_149_47.t2 30.461
R54 a_149_47.t0 a_149_47.n0 25.846
R55 B1.n0 B1.t1 241.534
R56 B1.n0 B1.t0 169.234
R57 B1 B1.n0 78.133
R58 a_512_297.t0 a_512_297.t1 41.37
R59 VPWR.n2 VPWR.n1 177.129
R60 VPWR.n2 VPWR.n0 169.715
R61 VPWR.n0 VPWR.t2 38.415
R62 VPWR.n1 VPWR.t3 34.475
R63 VPWR.n1 VPWR.t0 30.535
R64 VPWR.n0 VPWR.t1 26.595
R65 VPWR VPWR.n2 0.176
C0 X VGND 0.22fF
C1 VPWR X 0.22fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__o221a_2.ext - technology: sky130A

.subckt sky130_fd_sc_hd__o221a_2 B2 A2 X B1 C1 A1 VGND VPWR VNB VPB
X0 VPWR.t3 a_38_47.t4 X.t3 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 VPWR.t1 A1.t0 a_497_297.t1 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 X.t2 a_38_47.t5 VPWR.t2 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 a_141_47.t0 B2.t0 a_225_47.t0 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 a_497_297.t0 A2.t0 a_38_47.t2 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 VGND.t0 A1.t1 a_225_47.t1 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 VPWR.t0 C1.t0 a_38_47.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 a_237_297.t1 B1.t0 VPWR.t4 VPB.t6 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 a_38_47.t3 B2.t1 a_237_297.t0 VPB.t5 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 a_225_47.t2 A2.t1 VGND.t3 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 X.t1 a_38_47.t6 VGND.t2 VNB.t5 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 a_141_47.t1 C1.t1 a_38_47.t1 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 VGND.t1 a_38_47.t7 X.t0 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 a_225_47.t3 B1.t1 a_141_47.t2 VNB.t6 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
R0 a_38_47.n7 a_38_47.t1 226.774
R1 a_38_47.n0 a_38_47.t4 212.079
R2 a_38_47.n1 a_38_47.t5 212.079
R3 a_38_47.n4 a_38_47.n2 191.924
R4 a_38_47.t0 a_38_47.n7 169.343
R5 a_38_47.n4 a_38_47.n3 146.25
R6 a_38_47.n6 a_38_47.n5 146.25
R7 a_38_47.n0 a_38_47.t7 139.779
R8 a_38_47.n1 a_38_47.t6 139.779
R9 a_38_47.n7 a_38_47.n6 64.218
R10 a_38_47.n2 a_38_47.n0 37.975
R11 a_38_47.n3 a_38_47.t2 26.595
R12 a_38_47.n5 a_38_47.t3 26.595
R13 a_38_47.n2 a_38_47.n1 23.369
R14 a_38_47.n6 a_38_47.n4 10.955
R15 X X.n0 172.76
R16 X X.n1 101.698
R17 X.n0 X.t3 26.595
R18 X.n0 X.t2 26.595
R19 X.n1 X.t0 24.923
R20 X.n1 X.t1 24.923
R21 VPWR.n2 VPWR.t3 550.954
R22 VPWR.n12 VPWR.n11 170.114
R23 VPWR.n1 VPWR.n0 165.765
R24 VPWR.n0 VPWR.t2 38.415
R25 VPWR.n11 VPWR.t0 33.49
R26 VPWR.n11 VPWR.t4 31.52
R27 VPWR.n0 VPWR.t1 26.595
R28 VPWR.n13 VPWR.n12 8.664
R29 VPWR.n4 VPWR.n3 4.65
R30 VPWR.n6 VPWR.n5 4.65
R31 VPWR.n8 VPWR.n7 4.65
R32 VPWR.n10 VPWR.n9 4.65
R33 VPWR.n2 VPWR.n1 3.876
R34 VPWR.n4 VPWR.n2 0.242
R35 VPWR.n13 VPWR.n10 0.132
R36 VPWR VPWR.n13 0.13
R37 VPWR.n6 VPWR.n4 0.119
R38 VPWR.n8 VPWR.n6 0.119
R39 VPWR.n10 VPWR.n8 0.119
R40 VPB.t5 VPB.t1 547.507
R41 VPB VPB.t0 290.031
R42 VPB.t2 VPB.t3 284.112
R43 VPB.t0 VPB.t6 284.112
R44 VPB.t3 VPB.t4 248.598
R45 VPB.t6 VPB.t5 221.962
R46 VPB.t1 VPB.t2 213.084
R47 A1.n0 A1.t0 241.534
R48 A1.n0 A1.t1 169.234
R49 A1 A1.n0 80.266
R50 a_497_297.t0 a_497_297.t1 41.37
R51 B2.n0 B2.t1 233.868
R52 B2.n0 B2.t0 161.568
R53 B2.n1 B2.n0 76
R54 B2.n1 B2 12.579
R55 B2 B2.n1 2.427
R56 a_225_47.n1 a_225_47.n0 229.82
R57 a_225_47.n0 a_225_47.t1 24.923
R58 a_225_47.n0 a_225_47.t2 24.923
R59 a_225_47.t0 a_225_47.n1 24.923
R60 a_225_47.n1 a_225_47.t3 24.923
R61 a_141_47.t0 a_141_47.n0 331.323
R62 a_141_47.n0 a_141_47.t2 24.923
R63 a_141_47.n0 a_141_47.t1 24.923
R64 VNB VNB.t1 6972.59
R65 VNB.t0 VNB.t3 4545.05
R66 VNB.t5 VNB.t4 2030.77
R67 VNB.t2 VNB.t5 2030.77
R68 VNB.t3 VNB.t2 2030.77
R69 VNB.t6 VNB.t0 2030.77
R70 VNB.t1 VNB.t6 2030.77
R71 A2.n0 A2.t0 233.573
R72 A2.n0 A2.t1 161.273
R73 A2.n1 A2.n0 76
R74 A2.n1 A2 11.96
R75 A2 A2.n1 2.308
R76 VGND.n1 VGND.t1 199.091
R77 VGND.n0 VGND.t3 193.925
R78 VGND.n3 VGND.n2 74.837
R79 VGND.n2 VGND.t2 24.923
R80 VGND.n2 VGND.t0 24.923
R81 VGND.n8 VGND.n0 13.928
R82 VGND.n5 VGND.n4 4.65
R83 VGND.n7 VGND.n6 4.65
R84 VGND.n4 VGND.n3 3.764
R85 VGND.n5 VGND.n1 0.861
R86 VGND VGND.n8 0.492
R87 VGND.n8 VGND.n7 0.134
R88 VGND.n7 VGND.n5 0.119
R89 C1.n0 C1.t0 212.079
R90 C1.n0 C1.t1 133.353
R91 C1 C1.n0 132.074
R92 B1.n0 B1.t0 241.534
R93 B1.n0 B1.t1 169.234
R94 B1 B1.n0 78.04
R95 a_237_297.t0 a_237_297.t1 44.325
C0 VPWR X 0.26fF
C1 B2 A2 0.12fF
C2 X VGND 0.27fF
C3 A2 A1 0.10fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__o221a_4.ext - technology: sky130A

.subckt sky130_fd_sc_hd__o221a_4 C1 A1 A2 B1 B2 X VGND VPWR VNB VPB
X0 a_27_47.t1 B1.t0 a_277_47.t2 VNB.t6 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 a_109_47.t2 A2.t0 a_717_297.t1 VPB.t8 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 a_717_297.t2 A1.t0 VPWR.t8 VPB.t11 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 VGND.t7 A2.t1 a_277_47.t6 VNB.t10 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 a_277_297.t3 B2.t0 a_109_47.t3 VPB.t9 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 a_109_47.t4 B2.t1 a_277_297.t2 VPB.t10 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 VPWR.t3 a_109_47.t8 X.t7 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 X.t3 a_109_47.t9 VGND.t3 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 a_277_297.t1 B1.t1 VPWR.t6 VPB.t6 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 X.t6 a_109_47.t10 VPWR.t2 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 a_277_47.t5 A1.t1 VGND.t5 VNB.t9 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 a_277_47.t7 A2.t2 VGND.t6 VNB.t11 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 X.t2 a_109_47.t11 VGND.t2 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 VPWR.t4 C1.t0 a_109_47.t0 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14 a_27_47.t4 C1.t1 a_109_47.t5 VNB.t12 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X15 a_27_47.t2 B2.t2 a_277_47.t3 VNB.t7 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X16 VGND.t1 a_109_47.t12 X.t1 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X17 VGND.t4 A1.t2 a_277_47.t0 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X18 VGND.t0 a_109_47.t13 X.t0 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X19 a_277_47.t1 B1.t2 a_27_47.t0 VNB.t5 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X20 a_277_47.t4 B2.t3 a_27_47.t3 VNB.t8 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X21 VPWR.t1 a_109_47.t14 X.t5 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X22 VPWR.t5 B1.t3 a_277_297.t0 VPB.t5 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X23 X.t4 a_109_47.t15 VPWR.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X24 VPWR.t7 A1.t3 a_717_297.t3 VPB.t13 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X25 a_109_47.t6 C1.t2 VPWR.t9 VPB.t12 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X26 a_717_297.t0 A2.t3 a_109_47.t1 VPB.t7 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X27 a_109_47.t7 C1.t3 a_27_47.t5 VNB.t13 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
R0 B1.n1 B1.t1 241.534
R1 B1.n0 B1.t3 241.534
R2 B1.n1 B1.t2 169.234
R3 B1.n0 B1.t0 169.234
R4 B1.n2 B1.n0 162.716
R5 B1.n2 B1.n1 76
R6 B1 B1.n2 5.688
R7 a_277_47.n2 a_277_47.n1 133.853
R8 a_277_47.n2 a_277_47.n0 92.5
R9 a_277_47.n5 a_277_47.n4 89.082
R10 a_277_47.n4 a_277_47.n2 77.33
R11 a_277_47.n4 a_277_47.n3 51.267
R12 a_277_47.n3 a_277_47.t6 24.923
R13 a_277_47.n3 a_277_47.t5 24.923
R14 a_277_47.n1 a_277_47.t3 24.923
R15 a_277_47.n1 a_277_47.t1 24.923
R16 a_277_47.n0 a_277_47.t2 24.923
R17 a_277_47.n0 a_277_47.t4 24.923
R18 a_277_47.t0 a_277_47.n5 24.923
R19 a_277_47.n5 a_277_47.t7 24.923
R20 a_27_47.t1 a_27_47.n3 224.448
R21 a_27_47.n2 a_27_47.t5 134.628
R22 a_27_47.n3 a_27_47.n0 92.5
R23 a_27_47.n2 a_27_47.n1 50.599
R24 a_27_47.n3 a_27_47.n2 48.872
R25 a_27_47.n1 a_27_47.t0 24.923
R26 a_27_47.n1 a_27_47.t4 24.923
R27 a_27_47.n0 a_27_47.t3 24.923
R28 a_27_47.n0 a_27_47.t2 24.923
R29 VNB VNB.t13 6053.91
R30 VNB.t6 VNB.t9 4545.05
R31 VNB.t1 VNB.t3 2030.77
R32 VNB.t2 VNB.t1 2030.77
R33 VNB.t0 VNB.t2 2030.77
R34 VNB.t4 VNB.t0 2030.77
R35 VNB.t11 VNB.t4 2030.77
R36 VNB.t10 VNB.t11 2030.77
R37 VNB.t9 VNB.t10 2030.77
R38 VNB.t8 VNB.t6 2030.77
R39 VNB.t7 VNB.t8 2030.77
R40 VNB.t5 VNB.t7 2030.77
R41 VNB.t12 VNB.t5 2030.77
R42 VNB.t13 VNB.t12 2030.77
R43 A2.n0 A2.t3 212.079
R44 A2.n1 A2.t0 212.079
R45 A2.n0 A2.t2 139.779
R46 A2.n1 A2.t1 139.779
R47 A2 A2.n2 95.2
R48 A2.n2 A2.n0 30.672
R49 A2.n2 A2.n1 30.672
R50 a_717_297.n1 a_717_297.n0 638.833
R51 a_717_297.n0 a_717_297.t1 26.595
R52 a_717_297.n0 a_717_297.t2 26.595
R53 a_717_297.n1 a_717_297.t3 26.595
R54 a_717_297.t0 a_717_297.n1 26.595
R55 a_109_47.n13 a_109_47.n9 292.5
R56 a_109_47.n15 a_109_47.n14 292.5
R57 a_109_47.n0 a_109_47.t8 212.079
R58 a_109_47.n2 a_109_47.t10 212.079
R59 a_109_47.n5 a_109_47.t14 212.079
R60 a_109_47.n6 a_109_47.t15 212.079
R61 a_109_47.n14 a_109_47.n13 155.857
R62 a_109_47.n12 a_109_47.n11 146.733
R63 a_109_47.n0 a_109_47.t13 139.779
R64 a_109_47.n2 a_109_47.t11 139.779
R65 a_109_47.n5 a_109_47.t12 139.779
R66 a_109_47.n6 a_109_47.t9 139.779
R67 a_109_47.n14 a_109_47.n8 114.52
R68 a_109_47.n4 a_109_47.n1 104.8
R69 a_109_47.n12 a_109_47.n10 98.629
R70 a_109_47.n13 a_109_47.n12 81.971
R71 a_109_47.n8 a_109_47.n7 76
R72 a_109_47.n4 a_109_47.n3 76
R73 a_109_47.n3 a_109_47.n2 35.054
R74 a_109_47.n1 a_109_47.n0 30.672
R75 a_109_47.n7 a_109_47.n5 30.672
R76 a_109_47.n7 a_109_47.n6 30.672
R77 a_109_47.n9 a_109_47.t3 26.595
R78 a_109_47.n9 a_109_47.t4 26.595
R79 a_109_47.n10 a_109_47.t0 26.595
R80 a_109_47.n10 a_109_47.t6 26.595
R81 a_109_47.n15 a_109_47.t1 26.595
R82 a_109_47.t2 a_109_47.n15 26.595
R83 a_109_47.n8 a_109_47.n4 24.96
R84 a_109_47.n11 a_109_47.t5 24.923
R85 a_109_47.n11 a_109_47.t7 24.923
R86 VPB.t5 VPB.t11 556.386
R87 VPB.t2 VPB.t3 248.598
R88 VPB.t1 VPB.t2 248.598
R89 VPB.t0 VPB.t1 248.598
R90 VPB.t13 VPB.t0 248.598
R91 VPB.t7 VPB.t13 248.598
R92 VPB.t8 VPB.t7 248.598
R93 VPB.t11 VPB.t8 248.598
R94 VPB.t9 VPB.t5 248.598
R95 VPB.t10 VPB.t9 248.598
R96 VPB.t6 VPB.t10 248.598
R97 VPB.t4 VPB.t6 248.598
R98 VPB.t12 VPB.t4 248.598
R99 VPB VPB.t12 189.408
R100 A1.n1 A1.t3 241.534
R101 A1.n0 A1.t0 240.482
R102 A1.n3 A1.n0 171.339
R103 A1.n1 A1.t2 169.234
R104 A1.n0 A1.t1 168.182
R105 A1.n2 A1.n1 76
R106 A1 A1.n3 3.446
R107 A1.n2 A1 2.816
R108 A1.n3 A1.n2 0.768
R109 VPWR.n28 VPWR.n27 314.004
R110 VPWR.n6 VPWR.n5 314.004
R111 VPWR.n1 VPWR.n0 314.004
R112 VPWR.n18 VPWR.n17 292.5
R113 VPWR.n14 VPWR.n13 292.5
R114 VPWR.n2 VPWR.t3 202.206
R115 VPWR.n32 VPWR.t9 153.228
R116 VPWR.n17 VPWR.t5 28.565
R117 VPWR.n13 VPWR.t8 26.595
R118 VPWR.n27 VPWR.t6 26.595
R119 VPWR.n27 VPWR.t4 26.595
R120 VPWR.n5 VPWR.t0 26.595
R121 VPWR.n5 VPWR.t7 26.595
R122 VPWR.n0 VPWR.t2 26.595
R123 VPWR.n0 VPWR.t1 26.595
R124 VPWR.n4 VPWR.n3 4.65
R125 VPWR.n8 VPWR.n7 4.65
R126 VPWR.n10 VPWR.n9 4.65
R127 VPWR.n12 VPWR.n11 4.65
R128 VPWR.n16 VPWR.n15 4.65
R129 VPWR.n20 VPWR.n19 4.65
R130 VPWR.n22 VPWR.n21 4.65
R131 VPWR.n24 VPWR.n23 4.65
R132 VPWR.n26 VPWR.n25 4.65
R133 VPWR.n29 VPWR.n28 4.65
R134 VPWR.n31 VPWR.n30 4.65
R135 VPWR.n33 VPWR.n32 4.65
R136 VPWR.n15 VPWR.n14 4.234
R137 VPWR.n2 VPWR.n1 3.784
R138 VPWR.n19 VPWR.n18 3.764
R139 VPWR.n7 VPWR.n6 1.882
R140 VPWR.n4 VPWR.n2 0.233
R141 VPWR.n8 VPWR.n4 0.119
R142 VPWR.n10 VPWR.n8 0.119
R143 VPWR.n12 VPWR.n10 0.119
R144 VPWR.n16 VPWR.n12 0.119
R145 VPWR.n20 VPWR.n16 0.119
R146 VPWR.n22 VPWR.n20 0.119
R147 VPWR.n24 VPWR.n22 0.119
R148 VPWR.n26 VPWR.n24 0.119
R149 VPWR.n29 VPWR.n26 0.119
R150 VPWR.n31 VPWR.n29 0.119
R151 VPWR.n33 VPWR.n31 0.119
R152 VPWR VPWR.n33 0.02
R153 VGND.n17 VGND.t5 195.842
R154 VGND.n0 VGND.t0 193.644
R155 VGND.n2 VGND.n1 115.464
R156 VGND.n14 VGND.n13 115.464
R157 VGND.n8 VGND.n7 74.837
R158 VGND.n1 VGND.t2 24.923
R159 VGND.n1 VGND.t1 24.923
R160 VGND.n7 VGND.t3 24.923
R161 VGND.n7 VGND.t4 24.923
R162 VGND.n13 VGND.t6 24.923
R163 VGND.n13 VGND.t7 24.923
R164 VGND.n15 VGND.n14 17.317
R165 VGND.n9 VGND.n8 11.294
R166 VGND.n3 VGND.n2 5.27
R167 VGND.n18 VGND.n17 4.894
R168 VGND.n4 VGND.n3 4.65
R169 VGND.n6 VGND.n5 4.65
R170 VGND.n10 VGND.n9 4.65
R171 VGND.n12 VGND.n11 4.65
R172 VGND.n16 VGND.n15 4.65
R173 VGND.n19 VGND.n18 4.65
R174 VGND VGND.n20 0.723
R175 VGND.n4 VGND.n0 0.645
R176 VGND.n20 VGND.n19 0.134
R177 VGND.n6 VGND.n4 0.119
R178 VGND.n10 VGND.n6 0.119
R179 VGND.n12 VGND.n10 0.119
R180 VGND.n16 VGND.n12 0.119
R181 VGND.n19 VGND.n16 0.119
R182 B2.n0 B2.t0 212.079
R183 B2.n1 B2.t1 212.079
R184 B2.n0 B2.t3 139.779
R185 B2.n1 B2.t2 139.779
R186 B2 B2.n2 77.268
R187 B2.n2 B2.n0 30.672
R188 B2.n2 B2.n1 30.672
R189 a_277_297.n1 a_277_297.n0 638.834
R190 a_277_297.n0 a_277_297.t0 26.595
R191 a_277_297.n0 a_277_297.t3 26.595
R192 a_277_297.n1 a_277_297.t2 26.595
R193 a_277_297.t1 a_277_297.n1 26.595
R194 X.n2 X.n0 213.963
R195 X.n2 X.n1 111.272
R196 X.n5 X.n3 88.89
R197 X.n5 X.n4 52.624
R198 X X.n5 36.181
R199 X.n0 X.t5 26.595
R200 X.n0 X.t4 26.595
R201 X.n1 X.t7 26.595
R202 X.n1 X.t6 26.595
R203 X.n4 X.t0 24.923
R204 X.n4 X.t2 24.923
R205 X.n3 X.t1 24.923
R206 X.n3 X.t3 24.923
R207 X X.n2 18.964
R208 C1.n0 C1.t0 212.079
R209 C1.n1 C1.t2 212.079
R210 C1.n0 C1.t1 139.779
R211 C1.n1 C1.t3 139.779
R212 C1 C1.n1 112.481
R213 C1.n1 C1.n0 61.345
C0 VPWR X 0.48fF
C1 VPWR VGND 0.16fF
C2 B1 B2 0.33fF
C3 X VGND 0.51fF
C4 A1 A2 0.33fF
C5 VPB VPWR 0.15fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__o221ai_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__o221ai_1 A2 Y B1 C1 A1 B2 VGND VPWR VNB VPB
X0 a_109_47.t0 B1.t0 a_213_123.t0 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 Y.t2 B2.t0 a_295_297.t0 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 VPWR.t2 A1.t0 a_493_297.t1 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 a_213_123.t2 B2.t1 a_109_47.t1 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 a_295_297.t1 B1.t1 VPWR.t1 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 a_493_297.t0 A2.t0 Y.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 VPWR.t0 C1.t0 Y.t1 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 VGND.t0 A2.t1 a_213_123.t1 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 a_213_123.t3 A1.t1 VGND.t1 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 a_109_47.t2 C1.t1 Y.t3 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
R0 B1.n0 B1.t1 235.47
R1 B1.n0 B1.t0 163.17
R2 B1 B1.n0 83.951
R3 a_213_123.t0 a_213_123.n1 174.528
R4 a_213_123.n1 a_213_123.t3 168.142
R5 a_213_123.n1 a_213_123.n0 92.5
R6 a_213_123.n2 a_213_123.t0 64.8
R7 a_213_123.n0 a_213_123.t1 41.538
R8 a_213_123.n0 a_213_123.t2 24.923
R9 a_109_47.n0 a_109_47.t2 282.237
R10 a_109_47.n0 a_109_47.t1 24.923
R11 a_109_47.t0 a_109_47.n0 24.923
R12 VNB VNB.t3 6078.09
R13 VNB.t3 VNB.t0 4496.7
R14 VNB.t2 VNB.t1 2465.93
R15 VNB.t1 VNB.t4 2030.77
R16 VNB.t0 VNB.t2 2030.77
R17 B2.n0 B2.t0 241.534
R18 B2.n0 B2.t1 169.234
R19 B2 B2.n0 81.624
R20 a_295_297.t0 a_295_297.t1 47.28
R21 Y.n2 Y.t3 192.39
R22 Y.n2 Y.t1 155.79
R23 Y.n1 Y.n0 96.575
R24 Y Y.n2 69.558
R25 Y.n0 Y.t0 62.055
R26 Y.n0 Y.t2 26.595
R27 Y Y.n1 4.568
R28 Y.n1 Y 3.843
R29 VPB.t1 VPB.t3 538.629
R30 VPB.t2 VPB.t0 355.14
R31 VPB.t3 VPB.t2 230.841
R32 VPB.t0 VPB.t4 213.084
R33 VPB VPB.t1 204.205
R34 A1.n0 A1.t0 230.791
R35 A1.n0 A1.t1 158.491
R36 A1 A1.n0 77.53
R37 a_493_297.t0 a_493_297.t1 41.37
R38 VPWR.n0 VPWR.t2 155.966
R39 VPWR.n6 VPWR.n5 146.25
R40 VPWR.n2 VPWR.n1 146.25
R41 VPWR.n1 VPWR.t1 29.55
R42 VPWR.n5 VPWR.t0 29.55
R43 VPWR.n4 VPWR.n3 4.65
R44 VPWR.n7 VPWR.n6 4.369
R45 VPWR.n3 VPWR.n2 0.344
R46 VPWR.n4 VPWR.n0 0.141
R47 VPWR.n7 VPWR.n4 0.135
R48 VPWR VPWR.n7 0.125
R49 A2.n0 A2.t0 241.534
R50 A2.n0 A2.t1 169.234
R51 A2 A2.n0 116.532
R52 C1.n0 C1.t0 236.932
R53 C1.n0 C1.t1 205.73
R54 C1 C1.n0 85.115
R55 VGND VGND.n0 118.154
R56 VGND.n0 VGND.t1 24.923
R57 VGND.n0 VGND.t0 24.923
C0 Y VPWR 0.44fF
C1 C1 Y 0.17fF
C2 A2 VPWR 0.16fF
C3 B1 Y 0.14fF
C4 B1 B2 0.11fF
C5 B2 Y 0.13fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__o221ai_2.ext - technology: sky130A

.subckt sky130_fd_sc_hd__o221ai_2 B1 B2 Y A2 A1 C1 VGND VPWR VNB VPB
X0 Y.t7 A2.t0 a_734_297.t3 VPB.t8 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_300_47.t5 B2.t0 a_28_47.t3 VNB.t7 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 Y.t1 C1.t0 VPWR.t4 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 a_300_47.t6 B1.t0 a_28_47.t4 VNB.t8 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 a_300_47.t3 A2.t1 VGND.t3 VNB.t5 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 a_300_47.t1 A1.t0 VGND.t1 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 a_734_297.t0 A1.t1 VPWR.t0 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 a_28_47.t0 C1.t1 Y.t2 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 Y.t3 C1.t2 a_28_47.t1 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 VPWR.t3 C1.t3 Y.t4 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 VPWR.t5 B1.t1 a_382_297.t3 VPB.t9 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 a_382_297.t1 B2.t1 Y.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 a_28_47.t5 B1.t2 a_300_47.t7 VNB.t9 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 a_28_47.t2 B2.t2 a_300_47.t4 VNB.t6 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14 VGND.t0 A1.t2 a_300_47.t0 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X15 Y.t5 B2.t3 a_382_297.t0 VPB.t6 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16 VPWR.t1 A1.t3 a_734_297.t1 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17 VGND.t2 A2.t2 a_300_47.t2 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X18 a_382_297.t2 B1.t3 VPWR.t2 VPB.t5 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X19 a_734_297.t2 A2.t3 Y.t6 VPB.t7 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
R0 A2.n0 A2.t3 212.079
R1 A2.n1 A2.t0 212.079
R2 A2.n0 A2.t2 139.779
R3 A2.n1 A2.t1 139.779
R4 A2 A2.n2 81.12
R5 A2.n2 A2.n0 30.672
R6 A2.n2 A2.n1 30.672
R7 a_734_297.n1 a_734_297.n0 496.201
R8 a_734_297.n0 a_734_297.t1 26.595
R9 a_734_297.n0 a_734_297.t2 26.595
R10 a_734_297.n1 a_734_297.t3 26.595
R11 a_734_297.t0 a_734_297.n1 26.595
R12 Y.n2 Y.n0 415.604
R13 Y.n2 Y.n1 292.5
R14 Y.n5 Y.n4 144.625
R15 Y.n5 Y.n3 98.657
R16 Y Y.n2 64.563
R17 Y Y.n5 56.051
R18 Y.n3 Y.t4 26.595
R19 Y.n3 Y.t1 26.595
R20 Y.n1 Y.t0 26.595
R21 Y.n1 Y.t5 26.595
R22 Y.n0 Y.t6 26.595
R23 Y.n0 Y.t7 26.595
R24 Y.n4 Y.t2 24.923
R25 Y.n4 Y.t3 24.923
R26 VPB.t4 VPB.t5 556.386
R27 VPB.t9 VPB.t1 295.95
R28 VPB.t7 VPB.t2 248.598
R29 VPB.t8 VPB.t7 248.598
R30 VPB.t1 VPB.t8 248.598
R31 VPB.t0 VPB.t9 248.598
R32 VPB.t6 VPB.t0 248.598
R33 VPB.t5 VPB.t6 248.598
R34 VPB.t3 VPB.t4 248.598
R35 VPB VPB.t3 195.327
R36 B2.n0 B2.t1 212.079
R37 B2.n1 B2.t3 212.079
R38 B2.n0 B2.t2 139.779
R39 B2.n1 B2.t0 139.779
R40 B2 B2.n2 77.268
R41 B2.n2 B2.n0 30.672
R42 B2.n2 B2.n1 30.672
R43 a_28_47.t0 a_28_47.n3 172.93
R44 a_28_47.t0 a_28_47.n4 170.961
R45 a_28_47.n2 a_28_47.n0 133.853
R46 a_28_47.n4 a_28_47.t1 131.164
R47 a_28_47.n2 a_28_47.n1 92.5
R48 a_28_47.n3 a_28_47.n2 44.307
R49 a_28_47.n1 a_28_47.t3 24.923
R50 a_28_47.n1 a_28_47.t5 24.923
R51 a_28_47.n0 a_28_47.t4 24.923
R52 a_28_47.n0 a_28_47.t2 24.923
R53 a_300_47.n4 a_300_47.t7 219.833
R54 a_300_47.n1 a_300_47.t1 128.218
R55 a_300_47.n5 a_300_47.n4 92.5
R56 a_300_47.n1 a_300_47.n0 52.624
R57 a_300_47.n4 a_300_47.n3 51.051
R58 a_300_47.n3 a_300_47.n1 48.238
R59 a_300_47.n3 a_300_47.n2 43.173
R60 a_300_47.n2 a_300_47.t6 33.23
R61 a_300_47.n2 a_300_47.t0 31.384
R62 a_300_47.n0 a_300_47.t2 24.923
R63 a_300_47.n0 a_300_47.t3 24.923
R64 a_300_47.n5 a_300_47.t4 24.923
R65 a_300_47.t5 a_300_47.n5 24.923
R66 VNB VNB.t2 6102.26
R67 VNB.t1 VNB.t9 4545.05
R68 VNB.t8 VNB.t0 2417.58
R69 VNB.t4 VNB.t3 2030.77
R70 VNB.t5 VNB.t4 2030.77
R71 VNB.t0 VNB.t5 2030.77
R72 VNB.t6 VNB.t8 2030.77
R73 VNB.t7 VNB.t6 2030.77
R74 VNB.t9 VNB.t7 2030.77
R75 VNB.t2 VNB.t1 2030.77
R76 C1.n0 C1.t3 212.079
R77 C1.n1 C1.t0 212.079
R78 C1.n0 C1.t1 139.779
R79 C1.n1 C1.t2 139.779
R80 C1 C1.n1 113.942
R81 C1.n1 C1.n0 61.345
R82 VPWR.n1 VPWR.n0 308.79
R83 VPWR.n14 VPWR.n13 292.5
R84 VPWR.n10 VPWR.n9 292.5
R85 VPWR.n2 VPWR.t1 169.602
R86 VPWR.n19 VPWR.t4 153.228
R87 VPWR.n0 VPWR.t0 42.355
R88 VPWR.n9 VPWR.t2 26.595
R89 VPWR.n13 VPWR.t3 26.595
R90 VPWR.n0 VPWR.t5 26.595
R91 VPWR.n4 VPWR.n3 4.65
R92 VPWR.n6 VPWR.n5 4.65
R93 VPWR.n8 VPWR.n7 4.65
R94 VPWR.n12 VPWR.n11 4.65
R95 VPWR.n16 VPWR.n15 4.65
R96 VPWR.n18 VPWR.n17 4.65
R97 VPWR.n20 VPWR.n19 4.65
R98 VPWR.n2 VPWR.n1 4.078
R99 VPWR.n15 VPWR.n14 0.847
R100 VPWR.n11 VPWR.n10 0.282
R101 VPWR.n4 VPWR.n2 0.138
R102 VPWR.n6 VPWR.n4 0.119
R103 VPWR.n8 VPWR.n6 0.119
R104 VPWR.n12 VPWR.n8 0.119
R105 VPWR.n16 VPWR.n12 0.119
R106 VPWR.n18 VPWR.n16 0.119
R107 VPWR.n20 VPWR.n18 0.119
R108 VPWR VPWR.n20 0.022
R109 B1.n1 B1.t3 241.534
R110 B1.n0 B1.t1 241.534
R111 B1.n1 B1.t2 169.234
R112 B1.n0 B1.t0 169.234
R113 B1.n2 B1.n0 162.479
R114 B1.n2 B1.n1 76
R115 B1 B1.n2 18.251
R116 VGND.n2 VGND.n0 125.963
R117 VGND.n2 VGND.n1 123.951
R118 VGND.n0 VGND.t1 24.923
R119 VGND.n0 VGND.t2 24.923
R120 VGND.n1 VGND.t3 24.923
R121 VGND.n1 VGND.t0 24.923
R122 VGND VGND.n2 1.099
R123 A1.n0 A1.t3 241.534
R124 A1.n1 A1.t1 241.534
R125 A1.n2 A1.n1 184.186
R126 A1.n0 A1.t0 169.234
R127 A1.n1 A1.t2 169.234
R128 A1.n2 A1.n0 76
R129 A1 A1.n2 23.68
R130 a_382_297.n1 a_382_297.n0 638.833
R131 a_382_297.n0 a_382_297.t0 26.595
R132 a_382_297.n0 a_382_297.t2 26.595
R133 a_382_297.n1 a_382_297.t3 26.595
R134 a_382_297.t1 a_382_297.n1 26.595
C0 VPWR VPB 0.12fF
C1 A1 VPWR 0.10fF
C2 VPWR VGND 0.12fF
C3 A1 Y 0.16fF
C4 B1 B2 0.33fF
C5 A1 A2 0.31fF
C6 B1 Y 0.65fF
C7 B1 A1 0.14fF
C8 VPWR Y 0.54fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__o221ai_4.ext - technology: sky130A

.subckt sky130_fd_sc_hd__o221ai_4 B1 B2 A2 C1 Y A1 VGND VPWR VNB VPB
X0 a_471_47.t9 A2.t0 VGND.t3 VNB.t13 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 a_471_47.t2 B2.t0 a_27_47.t5 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 a_471_47.t8 A2.t1 VGND.t2 VNB.t12 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 Y.t11 C1.t0 VPWR.t7 VPB.t11 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 VPWR.t8 A1.t0 a_1241_297.t3 VPB.t16 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 a_471_47.t3 B2.t1 a_27_47.t4 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 a_471_47.t12 A1.t1 VGND.t4 VNB.t16 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 Y.t7 C1.t1 a_27_47.t6 VNB.t6 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 VPWR.t6 C1.t2 Y.t10 VPB.t10 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 a_1241_297.t2 A1.t2 VPWR.t9 VPB.t17 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 a_27_47.t3 B2.t2 a_471_47.t4 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 VPWR.t0 B1.t0 a_553_297.t3 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 VGND.t1 A2.t2 a_471_47.t7 VNB.t11 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 a_553_297.t2 B1.t1 VPWR.t1 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14 a_27_47.t2 B2.t3 a_471_47.t5 VNB.t5 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X15 VGND.t0 A2.t3 a_471_47.t6 VNB.t10 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X16 a_27_47.t7 C1.t3 Y.t6 VNB.t7 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X17 VGND.t5 A1.t3 a_471_47.t13 VNB.t17 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X18 Y.t5 C1.t4 a_27_47.t8 VNB.t8 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X19 a_27_47.t9 C1.t5 Y.t4 VNB.t9 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X20 a_1241_297.t1 A1.t4 VPWR.t10 VPB.t18 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X21 VPWR.t2 B1.t2 a_553_297.t1 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X22 VPWR.t11 A1.t5 a_1241_297.t0 VPB.t19 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X23 Y.t1 B2.t4 a_553_297.t7 VPB.t7 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X24 a_1241_297.t7 A2.t4 Y.t15 VPB.t15 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X25 Y.t9 C1.t6 VPWR.t5 VPB.t9 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X26 a_553_297.t6 B2.t5 Y.t0 VPB.t6 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X27 a_471_47.t14 A1.t6 VGND.t6 VNB.t18 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X28 Y.t14 A2.t5 a_1241_297.t6 VPB.t14 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X29 a_553_297.t5 B2.t6 Y.t3 VPB.t5 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X30 a_27_47.t0 B1.t3 a_471_47.t0 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X31 VGND.t7 A1.t7 a_471_47.t15 VNB.t19 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X32 Y.t2 B2.t7 a_553_297.t4 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X33 a_1241_297.t5 A2.t6 Y.t13 VPB.t13 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X34 a_27_47.t1 B1.t4 a_471_47.t1 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X35 a_553_297.t0 B1.t5 VPWR.t3 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X36 Y.t12 A2.t7 a_1241_297.t4 VPB.t12 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X37 VPWR.t4 C1.t7 Y.t8 VPB.t8 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X38 a_471_47.t10 B1.t6 a_27_47.t10 VNB.t14 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X39 a_471_47.t11 B1.t7 a_27_47.t11 VNB.t15 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
R0 A2.n0 A2.t4 212.079
R1 A2.n2 A2.t5 212.079
R2 A2.n7 A2.t6 212.079
R3 A2.n5 A2.t7 212.079
R4 A2.n0 A2.t3 139.779
R5 A2.n2 A2.t1 139.779
R6 A2.n7 A2.t2 139.779
R7 A2.n5 A2.t0 139.779
R8 A2.n9 A2.n6 97.76
R9 A2.n4 A2.n1 97.76
R10 A2.n4 A2.n3 76
R11 A2.n9 A2.n8 76
R12 A2.n1 A2.n0 21.909
R13 A2 A2.n4 16
R14 A2.n6 A2.n5 13.145
R15 A2.n3 A2.n2 10.224
R16 A2 A2.n9 5.76
R17 A2.n8 A2.n7 1.46
R18 VGND.n3 VGND.n0 124.319
R19 VGND.n2 VGND.n1 115.464
R20 VGND.n7 VGND.n6 115.464
R21 VGND.n13 VGND.n12 115.464
R22 VGND.n0 VGND.t6 24.923
R23 VGND.n0 VGND.t5 24.923
R24 VGND.n1 VGND.t4 24.923
R25 VGND.n1 VGND.t0 24.923
R26 VGND.n6 VGND.t2 24.923
R27 VGND.n6 VGND.t1 24.923
R28 VGND.n12 VGND.t3 24.923
R29 VGND.n12 VGND.t7 24.923
R30 VGND.n14 VGND.n13 13.928
R31 VGND.n3 VGND.n2 6.256
R32 VGND.n5 VGND.n4 4.65
R33 VGND.n9 VGND.n8 4.65
R34 VGND.n11 VGND.n10 4.65
R35 VGND.n8 VGND.n7 3.764
R36 VGND VGND.n14 1.56
R37 VGND.n5 VGND.n3 0.275
R38 VGND.n14 VGND.n11 0.134
R39 VGND.n9 VGND.n5 0.119
R40 VGND.n11 VGND.n9 0.119
R41 a_471_47.n7 a_471_47.t0 232.401
R42 a_471_47.n1 a_471_47.t14 128.218
R43 a_471_47.n9 a_471_47.n4 92.5
R44 a_471_47.n8 a_471_47.n5 92.5
R45 a_471_47.n7 a_471_47.n6 92.5
R46 a_471_47.n9 a_471_47.n8 61.44
R47 a_471_47.n8 a_471_47.n7 61.44
R48 a_471_47.n1 a_471_47.n0 52.624
R49 a_471_47.n3 a_471_47.n2 52.624
R50 a_471_47.n13 a_471_47.n12 52.623
R51 a_471_47.n11 a_471_47.n10 51.073
R52 a_471_47.n11 a_471_47.n9 48.287
R53 a_471_47.n12 a_471_47.n11 40.338
R54 a_471_47.n10 a_471_47.t11 39.692
R55 a_471_47.n3 a_471_47.n1 38.786
R56 a_471_47.n12 a_471_47.n3 36.266
R57 a_471_47.n10 a_471_47.t15 24.923
R58 a_471_47.n6 a_471_47.t1 24.923
R59 a_471_47.n6 a_471_47.t10 24.923
R60 a_471_47.n5 a_471_47.t5 24.923
R61 a_471_47.n5 a_471_47.t2 24.923
R62 a_471_47.n4 a_471_47.t4 24.923
R63 a_471_47.n4 a_471_47.t3 24.923
R64 a_471_47.n2 a_471_47.t6 24.923
R65 a_471_47.n2 a_471_47.t8 24.923
R66 a_471_47.n0 a_471_47.t13 24.923
R67 a_471_47.n0 a_471_47.t12 24.923
R68 a_471_47.n13 a_471_47.t7 24.923
R69 a_471_47.t9 a_471_47.n13 24.923
R70 VNB VNB.t8 6150.61
R71 VNB.t9 VNB.t0 4545.05
R72 VNB.t15 VNB.t19 2417.58
R73 VNB.t17 VNB.t18 2030.77
R74 VNB.t16 VNB.t17 2030.77
R75 VNB.t10 VNB.t16 2030.77
R76 VNB.t12 VNB.t10 2030.77
R77 VNB.t11 VNB.t12 2030.77
R78 VNB.t13 VNB.t11 2030.77
R79 VNB.t19 VNB.t13 2030.77
R80 VNB.t4 VNB.t15 2030.77
R81 VNB.t3 VNB.t4 2030.77
R82 VNB.t5 VNB.t3 2030.77
R83 VNB.t2 VNB.t5 2030.77
R84 VNB.t1 VNB.t2 2030.77
R85 VNB.t14 VNB.t1 2030.77
R86 VNB.t0 VNB.t14 2030.77
R87 VNB.t6 VNB.t9 2030.77
R88 VNB.t7 VNB.t6 2030.77
R89 VNB.t8 VNB.t7 2030.77
R90 B2.n0 B2.t5 212.079
R91 B2.n3 B2.t4 212.079
R92 B2.n2 B2.t6 212.079
R93 B2.n1 B2.t7 212.079
R94 B2.n0 B2.t2 139.779
R95 B2.n3 B2.t1 139.779
R96 B2.n2 B2.t3 139.779
R97 B2.n1 B2.t0 139.779
R98 B2.n3 B2.n2 61.345
R99 B2.n2 B2.n1 61.345
R100 B2 B2.n4 33.101
R101 B2.n4 B2.n0 29.379
R102 B2.n4 B2.n3 20.489
R103 a_27_47.n6 a_27_47.t9 170.961
R104 a_27_47.n2 a_27_47.n0 141.372
R105 a_27_47.n5 a_27_47.t8 132.021
R106 a_27_47.n2 a_27_47.n1 92.5
R107 a_27_47.n7 a_27_47.n3 92.5
R108 a_27_47.n5 a_27_47.n4 92.5
R109 a_27_47.n9 a_27_47.n8 92.5
R110 a_27_47.n7 a_27_47.n6 54.69
R111 a_27_47.n8 a_27_47.n2 48.872
R112 a_27_47.n8 a_27_47.n7 48.872
R113 a_27_47.n6 a_27_47.n5 48.872
R114 a_27_47.n4 a_27_47.t6 24.923
R115 a_27_47.n4 a_27_47.t7 24.923
R116 a_27_47.n3 a_27_47.t10 24.923
R117 a_27_47.n3 a_27_47.t0 24.923
R118 a_27_47.n1 a_27_47.t4 24.923
R119 a_27_47.n1 a_27_47.t2 24.923
R120 a_27_47.n0 a_27_47.t11 24.923
R121 a_27_47.n0 a_27_47.t3 24.923
R122 a_27_47.t5 a_27_47.n9 24.923
R123 a_27_47.n9 a_27_47.t1 24.923
R124 C1.n5 C1.t6 212.079
R125 C1.n0 C1.t7 212.079
R126 C1.n2 C1.t0 212.079
R127 C1.n6 C1.t2 212.079
R128 C1.n5 C1.t4 139.779
R129 C1.n0 C1.t5 139.779
R130 C1.n2 C1.t1 139.779
R131 C1.n6 C1.t3 139.779
R132 C1.n4 C1.n1 97.76
R133 C1.n4 C1.n3 76
R134 C1 C1.n7 48.615
R135 C1.n1 C1.n0 35.054
R136 C1.n7 C1.n6 28.577
R137 C1.n3 C1.n2 23.369
R138 C1.n7 C1.n5 21.73
R139 C1 C1.n4 6.4
R140 VPWR.n26 VPWR.n25 314.004
R141 VPWR.n1 VPWR.n0 314.004
R142 VPWR.n14 VPWR.n13 311.444
R143 VPWR.n36 VPWR.n35 292.5
R144 VPWR.n32 VPWR.n31 292.5
R145 VPWR.n42 VPWR.n41 170.445
R146 VPWR.n2 VPWR.t8 159.576
R147 VPWR.n46 VPWR.t5 153.228
R148 VPWR.n13 VPWR.t9 34.475
R149 VPWR.n13 VPWR.t2 34.475
R150 VPWR.n31 VPWR.t1 26.595
R151 VPWR.n35 VPWR.t4 26.595
R152 VPWR.n41 VPWR.t7 26.595
R153 VPWR.n41 VPWR.t6 26.595
R154 VPWR.n25 VPWR.t3 26.595
R155 VPWR.n25 VPWR.t0 26.595
R156 VPWR.n0 VPWR.t10 26.595
R157 VPWR.n0 VPWR.t11 26.595
R158 VPWR.n4 VPWR.n3 4.65
R159 VPWR.n6 VPWR.n5 4.65
R160 VPWR.n8 VPWR.n7 4.65
R161 VPWR.n10 VPWR.n9 4.65
R162 VPWR.n12 VPWR.n11 4.65
R163 VPWR.n16 VPWR.n15 4.65
R164 VPWR.n18 VPWR.n17 4.65
R165 VPWR.n20 VPWR.n19 4.65
R166 VPWR.n22 VPWR.n21 4.65
R167 VPWR.n24 VPWR.n23 4.65
R168 VPWR.n28 VPWR.n27 4.65
R169 VPWR.n30 VPWR.n29 4.65
R170 VPWR.n34 VPWR.n33 4.65
R171 VPWR.n38 VPWR.n37 4.65
R172 VPWR.n40 VPWR.n39 4.65
R173 VPWR.n43 VPWR.n42 4.65
R174 VPWR.n45 VPWR.n44 4.65
R175 VPWR.n47 VPWR.n46 4.65
R176 VPWR.n2 VPWR.n1 3.937
R177 VPWR.n37 VPWR.n36 2.07
R178 VPWR.n33 VPWR.n32 0.941
R179 VPWR.n15 VPWR.n14 0.376
R180 VPWR.n27 VPWR.n26 0.376
R181 VPWR.n4 VPWR.n2 0.28
R182 VPWR.n6 VPWR.n4 0.119
R183 VPWR.n8 VPWR.n6 0.119
R184 VPWR.n10 VPWR.n8 0.119
R185 VPWR.n12 VPWR.n10 0.119
R186 VPWR.n16 VPWR.n12 0.119
R187 VPWR.n18 VPWR.n16 0.119
R188 VPWR.n20 VPWR.n18 0.119
R189 VPWR.n22 VPWR.n20 0.119
R190 VPWR.n24 VPWR.n22 0.119
R191 VPWR.n28 VPWR.n24 0.119
R192 VPWR.n30 VPWR.n28 0.119
R193 VPWR.n34 VPWR.n30 0.119
R194 VPWR.n38 VPWR.n34 0.119
R195 VPWR.n40 VPWR.n38 0.119
R196 VPWR.n43 VPWR.n40 0.119
R197 VPWR.n45 VPWR.n43 0.119
R198 VPWR.n47 VPWR.n45 0.119
R199 VPWR VPWR.n47 0.02
R200 Y.n2 Y.n0 348.9
R201 Y.n12 Y.n4 292.5
R202 Y.n13 Y.n3 292.5
R203 Y.n2 Y.n1 292.5
R204 Y.n12 Y.n11 169.93
R205 Y.n10 Y.n9 158.833
R206 Y.n7 Y.n6 141.372
R207 Y.n10 Y.n8 99.473
R208 Y.n7 Y.n5 92.5
R209 Y Y.n13 80.772
R210 Y.n11 Y.n7 64.141
R211 Y.n13 Y.n12 55.457
R212 Y Y.n2 35.49
R213 Y.n1 Y.t13 26.595
R214 Y.n1 Y.t12 26.595
R215 Y.n3 Y.t0 26.595
R216 Y.n3 Y.t1 26.595
R217 Y.n4 Y.t3 26.595
R218 Y.n4 Y.t2 26.595
R219 Y.n8 Y.t8 26.595
R220 Y.n8 Y.t11 26.595
R221 Y.n9 Y.t10 26.595
R222 Y.n9 Y.t9 26.595
R223 Y.n0 Y.t15 26.595
R224 Y.n0 Y.t14 26.595
R225 Y.n5 Y.t4 24.923
R226 Y.n5 Y.t7 24.923
R227 Y.n6 Y.t6 24.923
R228 Y.n6 Y.t5 24.923
R229 Y.n11 Y.n10 12.047
R230 VPB.t8 VPB.t1 556.386
R231 VPB.t2 VPB.t17 295.95
R232 VPB.t18 VPB.t16 248.598
R233 VPB.t19 VPB.t18 248.598
R234 VPB.t15 VPB.t19 248.598
R235 VPB.t14 VPB.t15 248.598
R236 VPB.t13 VPB.t14 248.598
R237 VPB.t12 VPB.t13 248.598
R238 VPB.t17 VPB.t12 248.598
R239 VPB.t6 VPB.t2 248.598
R240 VPB.t7 VPB.t6 248.598
R241 VPB.t5 VPB.t7 248.598
R242 VPB.t4 VPB.t5 248.598
R243 VPB.t3 VPB.t4 248.598
R244 VPB.t0 VPB.t3 248.598
R245 VPB.t1 VPB.t0 248.598
R246 VPB.t11 VPB.t8 248.598
R247 VPB.t10 VPB.t11 248.598
R248 VPB.t9 VPB.t10 248.598
R249 VPB VPB.t9 201.246
R250 A1.n6 A1.n3 247.545
R251 A1.n3 A1.t2 241.534
R252 A1.n0 A1.t0 212.079
R253 A1.n1 A1.t4 212.079
R254 A1.n4 A1.t5 212.079
R255 A1.n3 A1.t7 169.234
R256 A1.n0 A1.t6 139.779
R257 A1.n1 A1.t3 139.779
R258 A1.n4 A1.t1 139.779
R259 A1.n6 A1.n5 76.724
R260 A1 A1.n2 46.695
R261 A1.n2 A1.n0 31.954
R262 A1.n2 A1.n1 18.353
R263 A1.n5 A1.n4 13.145
R264 A1 A1.n6 1.92
R265 a_1241_297.n2 a_1241_297.n1 345.898
R266 a_1241_297.n2 a_1241_297.n0 292.5
R267 a_1241_297.n5 a_1241_297.n4 160.328
R268 a_1241_297.n4 a_1241_297.n3 142.024
R269 a_1241_297.n4 a_1241_297.n2 61.677
R270 a_1241_297.n3 a_1241_297.t0 26.595
R271 a_1241_297.n3 a_1241_297.t7 26.595
R272 a_1241_297.n0 a_1241_297.t6 26.595
R273 a_1241_297.n0 a_1241_297.t5 26.595
R274 a_1241_297.n1 a_1241_297.t4 26.595
R275 a_1241_297.n1 a_1241_297.t2 26.595
R276 a_1241_297.t3 a_1241_297.n5 26.595
R277 a_1241_297.n5 a_1241_297.t1 26.595
R278 B1.n3 B1.n0 251.856
R279 B1.n0 B1.t2 241.534
R280 B1.n1 B1.t5 212.079
R281 B1.n4 B1.t0 212.079
R282 B1.n7 B1.t1 212.079
R283 B1.n0 B1.t7 169.234
R284 B1.n1 B1.t4 139.779
R285 B1.n4 B1.t6 139.779
R286 B1.n7 B1.t3 139.779
R287 B1 B1.n8 88.48
R288 B1.n3 B1.n2 76
R289 B1.n6 B1.n5 76
R290 B1.n6 B1.n3 21.76
R291 B1.n2 B1.n1 16.796
R292 B1 B1.n6 9.28
R293 B1.n8 B1.n7 6.572
R294 B1.n5 B1.n4 5.112
R295 a_553_297.n2 a_553_297.n0 346.71
R296 a_553_297.n2 a_553_297.n1 292.5
R297 a_553_297.n5 a_553_297.n4 215.002
R298 a_553_297.n4 a_553_297.n3 141.247
R299 a_553_297.n4 a_553_297.n2 67.836
R300 a_553_297.n3 a_553_297.t4 26.595
R301 a_553_297.n3 a_553_297.t0 26.595
R302 a_553_297.n1 a_553_297.t7 26.595
R303 a_553_297.n1 a_553_297.t5 26.595
R304 a_553_297.n0 a_553_297.t1 26.595
R305 a_553_297.n0 a_553_297.t6 26.595
R306 a_553_297.t3 a_553_297.n5 26.595
R307 a_553_297.n5 a_553_297.t2 26.595
C0 A1 A2 0.53fF
C1 B1 Y 0.74fF
C2 VPB VPWR 0.19fF
C3 B1 A1 0.13fF
C4 VPWR Y 0.67fF
C5 VPWR VGND 0.20fF
C6 A1 Y 0.30fF
C7 C1 Y 0.43fF
C8 B1 B2 0.37fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__o311a_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__o311a_1 X A1 A2 A3 B1 C1 VGND VPWR VNB VPB
X0 a_585_47.t0 B1.t0 a_266_47.t0 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 VGND.t2 A2.t0 a_266_47.t2 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 VPWR.t3 a_81_21.t4 X.t0 VPB.t5 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 a_81_21.t3 C1.t0 a_585_47.t1 VNB.t5 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 VGND.t1 a_81_21.t5 X.t1 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 a_266_297.t0 A1.t0 VPWR.t2 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 a_368_297.t0 A2.t1 a_266_297.t1 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 a_266_47.t1 A3.t0 VGND.t0 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 a_266_47.t3 A1.t1 VGND.t3 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 a_81_21.t2 A3.t1 a_368_297.t1 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 a_81_21.t1 C1.t1 VPWR.t1 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 VPWR.t0 B1.t1 a_81_21.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
R0 B1.n0 B1.t1 238.154
R1 B1.n0 B1.t0 165.854
R2 B1 B1.n0 88.218
R3 a_266_47.n1 a_266_47.n0 207.613
R4 a_266_47.n1 a_266_47.t1 34.153
R5 a_266_47.n0 a_266_47.t2 33.23
R6 a_266_47.n0 a_266_47.t3 33.23
R7 a_266_47.t0 a_266_47.n1 33.23
R8 a_585_47.t0 a_585_47.t1 38.769
R9 VNB VNB.t2 6150.61
R10 VNB.t2 VNB.t4 3747.25
R11 VNB.t3 VNB.t1 2756.04
R12 VNB.t1 VNB.t0 2490.11
R13 VNB.t4 VNB.t3 2465.93
R14 VNB.t0 VNB.t5 1740.66
R15 A2.n0 A2.t1 241.534
R16 A2.n0 A2.t0 169.234
R17 A2.n1 A2.n0 76
R18 A2 A2.n1 11.899
R19 A2.n1 A2 2.07
R20 VGND.n2 VGND.n1 96.575
R21 VGND.n0 VGND.t3 59.076
R22 VGND.n0 VGND.t1 56.307
R23 VGND.n1 VGND.t0 38.769
R24 VGND.n1 VGND.t2 38.769
R25 VGND.n2 VGND.n0 3.517
R26 VGND VGND.n2 0.226
R27 a_81_21.n2 a_81_21.n0 289.676
R28 a_81_21.n1 a_81_21.t1 240.523
R29 a_81_21.n0 a_81_21.t4 231.014
R30 a_81_21.n0 a_81_21.t5 158.714
R31 a_81_21.n1 a_81_21.t3 139.645
R32 a_81_21.n3 a_81_21.n2 91.914
R33 a_81_21.n2 a_81_21.n1 45.109
R34 a_81_21.n3 a_81_21.t2 27.58
R35 a_81_21.t0 a_81_21.n3 26.595
R36 X.n2 X.n1 292.5
R37 X.n1 X.n0 147.056
R38 X.n3 X.t1 117.423
R39 X.n1 X.t0 26.595
R40 X.n0 X 10.1
R41 X X.n3 8.77
R42 X X.n2 7.862
R43 X.n3 X 7.348
R44 X.n2 X 4.571
R45 X.n0 X 2.299
R46 VPWR.n2 VPWR.n1 175.545
R47 VPWR.n2 VPWR.n0 163.422
R48 VPWR.n0 VPWR.t2 69.935
R49 VPWR.n0 VPWR.t3 53.19
R50 VPWR.n1 VPWR.t1 29.55
R51 VPWR.n1 VPWR.t0 29.55
R52 VPWR VPWR.n2 0.16
R53 VPB.t5 VPB.t2 458.722
R54 VPB.t3 VPB.t4 337.383
R55 VPB.t2 VPB.t3 301.869
R56 VPB.t0 VPB.t1 266.355
R57 VPB.t4 VPB.t0 251.557
R58 VPB VPB.t5 201.246
R59 C1.n0 C1.t1 230.154
R60 C1.n0 C1.t0 157.854
R61 C1 C1.n0 78.909
R62 A1.n0 A1.t0 241.534
R63 A1.n0 A1.t1 169.234
R64 A1 A1.n0 81.236
R65 a_266_297.t0 a_266_297.t1 70.92
R66 a_368_297.t0 a_368_297.t1 82.74
R67 A3.n0 A3.t1 234.17
R68 A3.n0 A3.t0 161.87
R69 A3.n1 A3.n0 76
R70 A3 A3.n1 13.818
R71 A3.n1 A3 2.427
C0 X VPWR 0.16fF
C1 A2 A3 0.21fF
C2 X VGND 0.12fF
C3 A1 A2 0.10fF
C4 A3 B1 0.11fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__o311a_2.ext - technology: sky130A

.subckt sky130_fd_sc_hd__o311a_2 X A2 A3 A1 B1 C1 VPWR VGND VNB VPB
X0 X.t1 a_91_21.t4 VPWR.t4 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_91_21.t1 C1.t0 VPWR.t1 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 a_360_47.t2 A3.t0 VGND.t1 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 VPWR.t0 B1.t0 a_91_21.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 a_360_297.t1 A1.t0 VPWR.t2 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 VGND.t2 A2.t0 a_360_47.t3 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 a_360_47.t1 A1.t1 VGND.t0 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 VPWR.t3 a_91_21.t5 X.t0 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 VGND.t4 a_91_21.t6 X.t3 VNB.t6 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 X.t2 a_91_21.t7 VGND.t3 VNB.t5 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 a_677_47.t0 B1.t1 a_360_47.t0 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 a_460_297.t0 A2.t1 a_360_297.t0 VPB.t5 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 a_91_21.t2 C1.t1 a_677_47.t1 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 a_91_21.t3 A3.t1 a_460_297.t1 VPB.t6 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
R0 a_91_21.n3 a_91_21.n1 319.595
R1 a_91_21.n2 a_91_21.t1 240.523
R2 a_91_21.n1 a_91_21.t5 212.079
R3 a_91_21.n0 a_91_21.t4 212.079
R4 a_91_21.n1 a_91_21.t6 139.779
R5 a_91_21.n0 a_91_21.t7 139.779
R6 a_91_21.n2 a_91_21.t2 139.645
R7 a_91_21.n4 a_91_21.n3 91.914
R8 a_91_21.n1 a_91_21.n0 61.345
R9 a_91_21.n3 a_91_21.n2 45.109
R10 a_91_21.n4 a_91_21.t3 27.58
R11 a_91_21.t0 a_91_21.n4 26.595
R12 VPWR.n3 VPWR.n0 175.528
R13 VPWR.n2 VPWR.n1 160.619
R14 VPWR.n6 VPWR.t4 160.233
R15 VPWR.n1 VPWR.t2 69.935
R16 VPWR.n1 VPWR.t3 53.19
R17 VPWR.n0 VPWR.t1 29.55
R18 VPWR.n0 VPWR.t0 29.55
R19 VPWR.n5 VPWR.n4 4.65
R20 VPWR.n7 VPWR.n6 4.65
R21 VPWR.n3 VPWR.n2 3.508
R22 VPWR.n5 VPWR.n3 0.152
R23 VPWR.n7 VPWR.n5 0.119
R24 VPWR VPWR.n7 0.02
R25 X.n2 X.n1 292.5
R26 X.n1 X.n0 147.045
R27 X.n5 X.n4 92.5
R28 X.n1 X.t0 26.595
R29 X.n1 X.t1 26.595
R30 X.n4 X.t3 24.923
R31 X.n4 X.t2 24.923
R32 X.n3 X 19.692
R33 X.n0 X 9.96
R34 X.n3 X 9.374
R35 X X.n5 8.61
R36 X X.n2 7.752
R37 X.n5 X 7.214
R38 X.n2 X 4.507
R39 X X.n3 2.884
R40 X.n0 X 2.266
R41 VPB.t3 VPB.t2 458.722
R42 VPB.t5 VPB.t6 337.383
R43 VPB.t2 VPB.t5 295.95
R44 VPB.t0 VPB.t1 266.355
R45 VPB.t6 VPB.t0 251.557
R46 VPB.t4 VPB.t3 248.598
R47 VPB VPB.t4 224.922
R48 C1.n0 C1.t0 230.154
R49 C1.n0 C1.t1 157.854
R50 C1 C1.n0 78.909
R51 A3.n0 A3.t1 234.17
R52 A3.n0 A3.t0 161.87
R53 A3.n1 A3.n0 76
R54 A3 A3.n1 13.818
R55 A3.n1 A3 2.427
R56 VGND.n7 VGND.t3 102.155
R57 VGND.n1 VGND.n0 96.447
R58 VGND.n2 VGND.t0 59.076
R59 VGND.n2 VGND.t4 56.307
R60 VGND.n0 VGND.t1 38.769
R61 VGND.n0 VGND.t2 38.769
R62 VGND.n8 VGND.n7 4.65
R63 VGND.n4 VGND.n3 4.65
R64 VGND.n6 VGND.n5 4.65
R65 VGND.n3 VGND.n2 2.531
R66 VGND.n4 VGND.n1 0.213
R67 VGND.n6 VGND.n4 0.119
R68 VGND.n8 VGND.n6 0.119
R69 VGND VGND.n8 0.02
R70 a_360_47.n1 a_360_47.n0 207.887
R71 a_360_47.n1 a_360_47.t2 34.153
R72 a_360_47.n0 a_360_47.t3 33.23
R73 a_360_47.t0 a_360_47.n1 33.23
R74 a_360_47.n0 a_360_47.t1 31.384
R75 VNB VNB.t5 6344.02
R76 VNB.t6 VNB.t1 3747.25
R77 VNB.t3 VNB.t2 2756.04
R78 VNB.t2 VNB.t0 2490.11
R79 VNB.t1 VNB.t3 2417.58
R80 VNB.t5 VNB.t6 2030.77
R81 VNB.t0 VNB.t4 1740.66
R82 B1.n0 B1.t0 238.154
R83 B1.n0 B1.t1 165.854
R84 B1 B1.n0 88.218
R85 A1.n0 A1.t0 241.534
R86 A1.n0 A1.t1 169.234
R87 A1 A1.n0 81.236
R88 a_360_297.t0 a_360_297.t1 68.95
R89 A2.n0 A2.t1 241.534
R90 A2.n0 A2.t0 169.234
R91 A2.n1 A2.n0 76
R92 A2 A2.n1 12.088
R93 A2.n1 A2 2.133
R94 a_677_47.t0 a_677_47.t1 38.769
R95 a_460_297.t0 a_460_297.t1 82.74
C0 VPWR X 0.38fF
C1 A3 B1 0.11fF
C2 A2 A3 0.21fF
C3 X VGND 0.26fF
C4 A1 A2 0.10fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__o311a_4.ext - technology: sky130A

.subckt sky130_fd_sc_hd__o311a_4 A1 A2 A3 B1 C1 X VPWR VGND VNB VPB
X0 a_79_21.t5 C1.t0 VPWR.t9 VPB.t13 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_467_47.t3 C1.t1 a_79_21.t7 VNB.t13 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 VGND.t4 A2.t0 a_717_47.t6 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 a_467_47.t0 B1.t0 a_717_47.t3 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 VGND.t5 A1.t0 a_717_47.t7 VNB.t7 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 VPWR.t1 a_79_21.t8 X.t3 VPB.t11 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 a_79_21.t6 C1.t2 a_467_47.t2 VNB.t12 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 X.t2 a_79_21.t9 VPWR.t2 VPB.t10 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 a_717_47.t4 B1.t1 a_467_47.t1 VNB.t5 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 VPWR.t5 a_79_21.t10 X.t1 VPB.t9 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 VGND.t9 a_79_21.t11 X.t7 VNB.t11 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 VGND.t8 a_79_21.t12 X.t6 VNB.t10 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 VGND.t0 A3.t0 a_717_47.t0 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 a_1147_297.t1 A1.t1 VPWR.t7 VPB.t7 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14 VPWR.t0 A1.t2 a_1147_297.t0 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 X.t5 a_79_21.t13 VGND.t7 VNB.t9 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X16 a_1147_297.t3 A2.t1 a_875_297.t3 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17 VPWR.t3 B1.t2 a_79_21.t2 VPB.t5 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X18 a_79_21.t0 A3.t1 a_875_297.t1 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X19 a_875_297.t0 A3.t2 a_79_21.t1 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X20 a_79_21.t3 B1.t3 VPWR.t4 VPB.t6 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X21 a_875_297.t2 A2.t2 a_1147_297.t2 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X22 a_717_47.t1 A3.t3 VGND.t1 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X23 a_717_47.t5 A2.t3 VGND.t3 VNB.t6 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X24 a_717_47.t2 A1.t3 VGND.t2 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X25 X.t0 a_79_21.t14 VPWR.t6 VPB.t8 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X26 VPWR.t8 C1.t3 a_79_21.t4 VPB.t12 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X27 X.t4 a_79_21.t15 VGND.t6 VNB.t8 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
R0 C1.n1 C1.t0 247.617
R1 C1.n0 C1.t3 221.719
R2 C1.n0 C1.t1 173.064
R3 C1.n1 C1.t2 128.533
R4 C1.n3 C1.n2 76
R5 C1.n2 C1.n1 21.582
R6 C1 C1.n3 18.215
R7 C1.n2 C1.n0 12.949
R8 C1.n3 C1 4.43
R9 VPWR.n1 VPWR.t3 363.558
R10 VPWR.n2 VPWR.n0 167.67
R11 VPWR.n16 VPWR.n15 163.438
R12 VPWR.n6 VPWR.n5 163.438
R13 VPWR.n20 VPWR.t6 145.234
R14 VPWR.n10 VPWR.t9 60.085
R15 VPWR.n10 VPWR.t1 60.085
R16 VPWR.n15 VPWR.t2 26.595
R17 VPWR.n15 VPWR.t5 26.595
R18 VPWR.n5 VPWR.t4 26.595
R19 VPWR.n5 VPWR.t8 26.595
R20 VPWR.n0 VPWR.t7 26.595
R21 VPWR.n0 VPWR.t0 26.595
R22 VPWR.n4 VPWR.n3 4.65
R23 VPWR.n7 VPWR.n6 4.65
R24 VPWR.n9 VPWR.n8 4.65
R25 VPWR.n12 VPWR.n11 4.65
R26 VPWR.n14 VPWR.n13 4.65
R27 VPWR.n17 VPWR.n16 4.65
R28 VPWR.n19 VPWR.n18 4.65
R29 VPWR.n21 VPWR.n20 4.65
R30 VPWR.n2 VPWR.n1 3.984
R31 VPWR.n11 VPWR.n10 0.562
R32 VPWR.n4 VPWR.n2 0.138
R33 VPWR.n7 VPWR.n4 0.119
R34 VPWR.n9 VPWR.n7 0.119
R35 VPWR.n12 VPWR.n9 0.119
R36 VPWR.n14 VPWR.n12 0.119
R37 VPWR.n17 VPWR.n14 0.119
R38 VPWR.n19 VPWR.n17 0.119
R39 VPWR.n21 VPWR.n19 0.119
R40 VPWR VPWR.n21 0.02
R41 a_79_21.n2 a_79_21.n1 372.876
R42 a_79_21.n10 a_79_21.t8 212.079
R43 a_79_21.n7 a_79_21.t9 212.079
R44 a_79_21.n5 a_79_21.t10 212.079
R45 a_79_21.n4 a_79_21.t14 212.079
R46 a_79_21.n12 a_79_21.n3 172.275
R47 a_79_21.n14 a_79_21.n13 159.159
R48 a_79_21.n2 a_79_21.n0 159.159
R49 a_79_21.n10 a_79_21.t12 139.779
R50 a_79_21.n7 a_79_21.t13 139.779
R51 a_79_21.n5 a_79_21.t11 139.779
R52 a_79_21.n4 a_79_21.t15 139.779
R53 a_79_21.n9 a_79_21.n6 92.738
R54 a_79_21.n11 a_79_21.n10 83.303
R55 a_79_21.n9 a_79_21.n8 76
R56 a_79_21.n5 a_79_21.n4 61.345
R57 a_79_21.n13 a_79_21.n12 57.6
R58 a_79_21.n13 a_79_21.n2 44.8
R59 a_79_21.n6 a_79_21.n5 30.672
R60 a_79_21.n1 a_79_21.t1 26.595
R61 a_79_21.n1 a_79_21.t0 26.595
R62 a_79_21.n0 a_79_21.t2 26.595
R63 a_79_21.n0 a_79_21.t3 26.595
R64 a_79_21.n14 a_79_21.t4 26.595
R65 a_79_21.t5 a_79_21.n14 26.595
R66 a_79_21.n3 a_79_21.t7 24.923
R67 a_79_21.n3 a_79_21.t6 24.923
R68 a_79_21.n8 a_79_21.n7 18.987
R69 a_79_21.n11 a_79_21.n9 16.738
R70 a_79_21.n12 a_79_21.n11 3.938
R71 VPB.t5 VPB.t0 568.224
R72 VPB.t1 VPB.t3 556.386
R73 VPB.t11 VPB.t13 449.844
R74 VPB.t4 VPB.t7 248.598
R75 VPB.t2 VPB.t4 248.598
R76 VPB.t3 VPB.t2 248.598
R77 VPB.t0 VPB.t1 248.598
R78 VPB.t6 VPB.t5 248.598
R79 VPB.t12 VPB.t6 248.598
R80 VPB.t13 VPB.t12 248.598
R81 VPB.t10 VPB.t11 248.598
R82 VPB.t9 VPB.t10 248.598
R83 VPB.t8 VPB.t9 248.598
R84 VPB VPB.t8 189.408
R85 a_467_47.n1 a_467_47.t0 218.584
R86 a_467_47.t2 a_467_47.n1 218.584
R87 a_467_47.n1 a_467_47.n0 49.651
R88 a_467_47.n0 a_467_47.t1 24.923
R89 a_467_47.n0 a_467_47.t3 24.923
R90 VNB VNB.t8 6053.91
R91 VNB.t4 VNB.t0 4593.41
R92 VNB.t10 VNB.t12 4545.05
R93 VNB.t0 VNB.t1 3723.08
R94 VNB.t7 VNB.t3 2030.77
R95 VNB.t6 VNB.t7 2030.77
R96 VNB.t2 VNB.t6 2030.77
R97 VNB.t1 VNB.t2 2030.77
R98 VNB.t5 VNB.t4 2030.77
R99 VNB.t13 VNB.t5 2030.77
R100 VNB.t12 VNB.t13 2030.77
R101 VNB.t9 VNB.t10 2030.77
R102 VNB.t11 VNB.t9 2030.77
R103 VNB.t8 VNB.t11 2030.77
R104 A2.n0 A2.t1 221.719
R105 A2.n1 A2.t2 221.719
R106 A2.n0 A2.t3 149.419
R107 A2.n1 A2.t0 149.419
R108 A2.n3 A2.n2 76
R109 A2.n2 A2.n0 51.77
R110 A2.n2 A2.n1 23.207
R111 A2.n3 A2 19.2
R112 A2 A2.n3 3.446
R113 a_717_47.n1 a_717_47.t2 214.091
R114 a_717_47.t0 a_717_47.n5 166.346
R115 a_717_47.n5 a_717_47.n4 142.886
R116 a_717_47.n1 a_717_47.n0 92.5
R117 a_717_47.n3 a_717_47.n2 92.5
R118 a_717_47.n5 a_717_47.n3 69.078
R119 a_717_47.n3 a_717_47.n1 51.2
R120 a_717_47.n4 a_717_47.t3 24.923
R121 a_717_47.n4 a_717_47.t4 24.923
R122 a_717_47.n2 a_717_47.t6 24.923
R123 a_717_47.n2 a_717_47.t1 24.923
R124 a_717_47.n0 a_717_47.t7 24.923
R125 a_717_47.n0 a_717_47.t5 24.923
R126 VGND.n24 VGND.t8 195.032
R127 VGND.n3 VGND.n0 109.971
R128 VGND.n2 VGND.n1 106.463
R129 VGND.n30 VGND.n29 106.463
R130 VGND.n34 VGND.t6 102.978
R131 VGND.n7 VGND.n6 92.5
R132 VGND.n9 VGND.n8 92.5
R133 VGND.n6 VGND.t1 25.846
R134 VGND.n8 VGND.t0 25.846
R135 VGND.n0 VGND.t2 24.923
R136 VGND.n0 VGND.t5 24.923
R137 VGND.n1 VGND.t3 24.923
R138 VGND.n1 VGND.t4 24.923
R139 VGND.n29 VGND.t7 24.923
R140 VGND.n29 VGND.t9 24.923
R141 VGND.n35 VGND.n34 4.65
R142 VGND.n5 VGND.n4 4.65
R143 VGND.n11 VGND.n10 4.65
R144 VGND.n13 VGND.n12 4.65
R145 VGND.n15 VGND.n14 4.65
R146 VGND.n17 VGND.n16 4.65
R147 VGND.n19 VGND.n18 4.65
R148 VGND.n21 VGND.n20 4.65
R149 VGND.n23 VGND.n22 4.65
R150 VGND.n26 VGND.n25 4.65
R151 VGND.n28 VGND.n27 4.65
R152 VGND.n31 VGND.n30 4.65
R153 VGND.n33 VGND.n32 4.65
R154 VGND.n10 VGND.n9 4.23
R155 VGND.n3 VGND.n2 3.671
R156 VGND.n25 VGND.n24 3.388
R157 VGND.n10 VGND.n7 3.145
R158 VGND.n5 VGND.n3 0.256
R159 VGND.n11 VGND.n5 0.119
R160 VGND.n13 VGND.n11 0.119
R161 VGND.n15 VGND.n13 0.119
R162 VGND.n17 VGND.n15 0.119
R163 VGND.n19 VGND.n17 0.119
R164 VGND.n21 VGND.n19 0.119
R165 VGND.n23 VGND.n21 0.119
R166 VGND.n26 VGND.n23 0.119
R167 VGND.n28 VGND.n26 0.119
R168 VGND.n31 VGND.n28 0.119
R169 VGND.n33 VGND.n31 0.119
R170 VGND.n35 VGND.n33 0.119
R171 VGND VGND.n35 0.02
R172 B1.n1 B1.t3 229.905
R173 B1.n0 B1.t2 184.766
R174 B1.n0 B1.t0 180.658
R175 B1.n1 B1.t1 139.779
R176 B1.n3 B1.n2 76
R177 B1.n2 B1.n1 22.067
R178 B1 B1.n3 16.246
R179 B1.n3 B1 6.4
R180 B1.n2 B1.n0 5.807
R181 A1.n0 A1.t1 237.653
R182 A1.n2 A1.t2 221.719
R183 A1.n0 A1.t3 165.353
R184 A1.n2 A1.t0 149.419
R185 A1.n1 A1.n0 76
R186 A1.n4 A1.n3 76
R187 A1.n3 A1.n2 36.596
R188 A1.n4 A1.n1 16.738
R189 A1 A1.n4 3.2
R190 A1.n1 A1 2.707
R191 X.n2 X.n1 203.959
R192 X.n2 X.n0 159.159
R193 X.n5 X.n3 155.747
R194 X.n5 X.n4 92.5
R195 X.n0 X.t1 26.595
R196 X.n0 X.t0 26.595
R197 X.n1 X.t3 26.595
R198 X.n1 X.t2 26.595
R199 X X.n6 26.092
R200 X.n3 X.t6 24.923
R201 X.n3 X.t5 24.923
R202 X.n4 X.t7 24.923
R203 X.n4 X.t4 24.923
R204 X.n6 X.n2 12.8
R205 X.n6 X.n5 12.8
R206 A3.n6 A3.t1 241.356
R207 A3.n2 A3.t2 221.719
R208 A3.n1 A3.t3 176.196
R209 A3.n5 A3.t0 149.419
R210 A3.n1 A3.n0 76
R211 A3.n4 A3.n3 76
R212 A3.n7 A3.n6 76
R213 A3.n3 A3.n1 60.696
R214 A3.n7 A3.n4 16.738
R215 A3.n0 A3 14.276
R216 A3.n6 A3.n5 10.711
R217 A3.n0 A3 8.369
R218 A3.n3 A3.n2 5.355
R219 A3 A3.n7 3.446
R220 A3.n4 A3 2.461
R221 a_1147_297.n1 a_1147_297.t2 472.325
R222 a_1147_297.n1 a_1147_297.n0 299.276
R223 a_1147_297.t1 a_1147_297.n1 264.336
R224 a_1147_297.n0 a_1147_297.t0 26.595
R225 a_1147_297.n0 a_1147_297.t3 26.595
R226 a_875_297.n1 a_875_297.t0 456.143
R227 a_875_297.t1 a_875_297.n1 375.93
R228 a_875_297.n1 a_875_297.n0 194.673
R229 a_875_297.n0 a_875_297.t3 26.595
R230 a_875_297.n0 a_875_297.t2 26.595
C0 X VGND 0.43fF
C1 VPB VPWR 0.16fF
C2 VPWR X 0.52fF
C3 VPWR VGND 0.17fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__o311ai_0.ext - technology: sky130A

.subckt sky130_fd_sc_hd__o311ai_0 A2 C1 A1 Y A3 B1 VGND VPWR VNB VPB
X0 VGND.t2 A2.t0 a_138_47.t3 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1 a_138_369.t0 A1.t0 VPWR.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X2 a_138_47.t0 A1.t1 VGND.t0 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3 a_138_47.t1 A3.t0 VGND.t1 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 Y.t1 C1.t0 a_458_47.t0 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 Y.t2 C1.t1 VPWR.t1 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X6 Y.t0 A3.t1 a_222_369.t0 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X7 a_222_369.t1 A2.t1 a_138_369.t1 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X8 a_458_47.t1 B1.t0 a_138_47.t2 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9 VPWR.t2 B1.t1 Y.t3 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
R0 A2.n0 A2.t1 299.374
R1 A2.n0 A2.t0 206.188
R2 A2.n1 A2.n0 76
R3 A2.n1 A2 11.767
R4 A2 A2.n1 2.27
R5 a_138_47.n1 a_138_47.n0 279.869
R6 a_138_47.n0 a_138_47.t2 135.714
R7 a_138_47.n0 a_138_47.t1 38.571
R8 a_138_47.n1 a_138_47.t3 38.571
R9 a_138_47.t0 a_138_47.n1 38.571
R10 VGND.n1 VGND.t0 136.222
R11 VGND.n1 VGND.n0 109.848
R12 VGND.n0 VGND.t1 38.571
R13 VGND.n0 VGND.t2 38.571
R14 VGND VGND.n1 0.217
R15 VNB VNB.t0 7408.82
R16 VNB.t2 VNB.t3 4917.65
R17 VNB.t4 VNB.t2 2717.65
R18 VNB.t0 VNB.t4 2717.65
R19 VNB.t3 VNB.t1 2329.41
R20 A1.n0 A1.t0 288.854
R21 A1.n0 A1.t1 195.668
R22 A1.n1 A1.n0 76
R23 A1.n2 A1 6.07
R24 A1.n1 A1 4.063
R25 A1 A1.n2 3.657
R26 A1.n2 A1.n1 1.625
R27 VPWR.n1 VPWR.t0 216.827
R28 VPWR.n1 VPWR.n0 169.294
R29 VPWR.n0 VPWR.t1 56.945
R30 VPWR.n0 VPWR.t2 56.945
R31 VPWR VPWR.n1 0.096
R32 a_138_369.t0 a_138_369.t1 83.109
R33 VPB.t1 VPB.t4 355.14
R34 VPB.t4 VPB.t3 307.788
R35 VPB VPB.t0 278.193
R36 VPB.t2 VPB.t1 248.598
R37 VPB.t0 VPB.t2 248.598
R38 A3.n0 A3.t1 299.374
R39 A3.n0 A3.t0 206.188
R40 A3 A3.n0 78.011
R41 C1.n0 C1.t1 269.919
R42 C1.n0 C1.t0 176.733
R43 C1 C1.n0 127.968
R44 a_458_47.t0 a_458_47.t1 60
R45 Y.n0 Y.t2 200.789
R46 Y.n2 Y.n1 146.71
R47 Y.n4 Y.t1 131.071
R48 Y.n1 Y.t3 69.257
R49 Y.n1 Y.t0 69.257
R50 Y.n3 Y 28.767
R51 Y Y.n5 10.12
R52 Y.n5 Y.n4 8.847
R53 Y.n3 Y 7.905
R54 Y Y.n0 7.239
R55 Y Y.n2 6.38
R56 Y.n4 Y 4.517
R57 Y.n5 Y 3.952
R58 Y Y.n3 2.976
R59 Y.n0 Y 1.72
R60 Y.n2 Y 1.518
R61 a_222_369.t0 a_222_369.t1 83.109
R62 B1.n0 B1.t1 295.573
R63 B1.n0 B1.t0 202.387
R64 B1 B1.n0 77.562
C0 Y VGND 0.13fF
C1 C1 Y 0.22fF
C2 A2 Y 0.16fF
C3 A1 A2 0.20fF
C4 VPWR Y 0.48fF
C5 A3 B1 0.10fF
C6 A1 VPWR 0.14fF
C7 B1 Y 0.16fF
C8 A2 VPWR 0.12fF
C9 A2 A3 0.15fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__o311ai_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__o311ai_1 Y A1 A2 A3 B1 C1 VGND VPWR VNB VPB
X0 VGND.t0 A2.t0 a_138_47.t1 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 a_138_47.t3 A1.t0 VGND.t2 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 Y.t3 C1.t0 VPWR.t2 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 a_138_47.t2 A3.t0 VGND.t1 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 Y.t1 A3.t1 a_222_297.t1 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 Y.t2 C1.t1 a_458_47.t1 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 a_222_297.t0 A2.t1 a_138_297.t0 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 VPWR.t0 B1.t0 Y.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 a_458_47.t0 B1.t1 a_138_47.t0 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 a_138_297.t1 A1.t1 VPWR.t1 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
R0 A2.n0 A2.t1 241.534
R1 A2.n0 A2.t0 169.234
R2 A2 A2.n0 78.27
R3 a_138_47.n1 a_138_47.n0 264.811
R4 a_138_47.t0 a_138_47.n1 87.692
R5 a_138_47.n0 a_138_47.t1 24.923
R6 a_138_47.n0 a_138_47.t3 24.923
R7 a_138_47.n1 a_138_47.t2 24.923
R8 VGND.n1 VGND.n0 109.883
R9 VGND.n1 VGND.t2 97.504
R10 VGND.n0 VGND.t1 24.923
R11 VGND.n0 VGND.t0 24.923
R12 VGND VGND.n1 0.177
R13 VNB VNB.t4 6779.19
R14 VNB.t3 VNB.t0 3674.73
R15 VNB.t1 VNB.t3 2030.77
R16 VNB.t4 VNB.t1 2030.77
R17 VNB.t0 VNB.t2 1740.66
R18 A1.n0 A1.t1 231.014
R19 A1.n0 A1.t0 158.714
R20 A1.n1 A1.n0 76
R21 A1.n1 A1 10.084
R22 A1 A1.n1 7.757
R23 C1.n0 C1.t0 212.079
R24 C1.n0 C1.t1 139.779
R25 C1 C1.n0 127.968
R26 VPWR.n1 VPWR.n0 170.651
R27 VPWR.n1 VPWR.t1 137.371
R28 VPWR.n0 VPWR.t2 36.445
R29 VPWR.n0 VPWR.t0 36.445
R30 VPWR VPWR.n1 0.096
R31 Y.n6 Y.n5 292.5
R32 Y.n3 Y.n2 292.5
R33 Y.n2 Y.n1 146.315
R34 Y.n5 Y.n4 146.308
R35 Y.n0 Y.t2 81.187
R36 Y.n5 Y.t0 44.325
R37 Y.n5 Y.t1 44.325
R38 Y Y.n6 35.941
R39 Y.n2 Y.t3 32.505
R40 Y.n7 Y.n3 19.952
R41 Y.n8 Y 16.669
R42 Y.n3 Y 8.814
R43 Y.n7 Y 7.905
R44 Y.n1 Y 6.763
R45 Y.n4 Y 5.967
R46 Y.n6 Y 3.84
R47 Y Y.n8 3.572
R48 Y Y.n0 3.514
R49 Y Y.n7 2.976
R50 Y.n0 Y 2.716
R51 Y.n1 Y 2.178
R52 Y.n4 Y 1.921
R53 Y.n8 Y 1.113
R54 VPB.t2 VPB.t0 355.14
R55 VPB.t0 VPB.t4 307.788
R56 VPB VPB.t3 278.193
R57 VPB.t1 VPB.t2 248.598
R58 VPB.t3 VPB.t1 248.598
R59 A3.n0 A3.t1 241.534
R60 A3.n0 A3.t0 169.234
R61 A3 A3.n0 78.011
R62 a_222_297.t0 a_222_297.t1 53.19
R63 a_458_47.t0 a_458_47.t1 38.769
R64 a_138_297.t0 a_138_297.t1 53.19
R65 B1.n0 B1.t0 237.733
R66 B1.n0 B1.t1 165.433
R67 B1 B1.n0 77.655
C0 A2 Y 0.16fF
C1 A1 A2 0.11fF
C2 VPWR Y 0.49fF
C3 A1 VPWR 0.14fF
C4 B1 Y 0.16fF
C5 A2 VPWR 0.14fF
C6 A2 A3 0.11fF
C7 Y VGND 0.14fF
C8 C1 Y 0.18fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__o311ai_2.ext - technology: sky130A

.subckt sky130_fd_sc_hd__o311ai_2 A1 Y C1 B1 A3 A2 VGND VPWR VNB VPB
X0 VPWR.t5 A1.t0 a_51_297.t3 VPB.t9 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_55_47.t7 A1.t1 VGND.t5 VNB.t9 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 Y.t5 C1.t0 a_729_47.t3 VNB.t6 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 VPWR.t2 C1.t1 Y.t7 VPB.t6 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 Y.t6 C1.t2 VPWR.t3 VPB.t7 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 a_55_47.t0 A3.t0 VGND.t0 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 VGND.t4 A1.t2 a_55_47.t6 VNB.t8 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 a_55_47.t3 B1.t0 a_729_47.t0 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 VGND.t3 A2.t0 a_55_47.t5 VNB.t5 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 Y.t2 B1.t1 VPWR.t0 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 VGND.t1 A3.t1 a_55_47.t1 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 a_729_47.t2 C1.t3 Y.t4 VNB.t7 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 a_51_297.t0 A2.t1 a_301_297.t3 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13 a_729_47.t1 B1.t2 a_55_47.t4 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14 a_301_297.t2 A2.t2 a_51_297.t1 VPB.t5 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 a_55_47.t2 A2.t3 VGND.t2 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X16 VPWR.t1 B1.t3 Y.t3 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17 a_51_297.t2 A1.t3 VPWR.t4 VPB.t8 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X18 Y.t0 A3.t2 a_301_297.t1 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X19 a_301_297.t0 A3.t3 Y.t1 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
R0 A1.n3 A1.t0 223.504
R1 A1.n0 A1.t3 221.719
R2 A1.n0 A1.t1 152.989
R3 A1.n2 A1.t2 149.419
R4 A1 A1.n1 92.492
R5 A1.n4 A1.n3 76
R6 A1.n4 A1 22.4
R7 A1.n1 A1.n0 12.496
R8 A1.n3 A1.n2 1.785
R9 A1 A1.n4 0.246
R10 a_51_297.t0 a_51_297.n1 472.325
R11 a_51_297.n1 a_51_297.t3 260.818
R12 a_51_297.n1 a_51_297.n0 159.159
R13 a_51_297.n0 a_51_297.t1 26.595
R14 a_51_297.n0 a_51_297.t2 26.595
R15 VPWR.n1 VPWR.n0 166.823
R16 VPWR.n18 VPWR.n17 163.438
R17 VPWR.n2 VPWR.t0 60.085
R18 VPWR.n2 VPWR.t1 60.085
R19 VPWR.n0 VPWR.t3 26.595
R20 VPWR.n0 VPWR.t2 26.595
R21 VPWR.n17 VPWR.t4 26.595
R22 VPWR.n17 VPWR.t5 26.595
R23 VPWR.n4 VPWR.n3 4.65
R24 VPWR.n6 VPWR.n5 4.65
R25 VPWR.n8 VPWR.n7 4.65
R26 VPWR.n10 VPWR.n9 4.65
R27 VPWR.n12 VPWR.n11 4.65
R28 VPWR.n14 VPWR.n13 4.65
R29 VPWR.n16 VPWR.n15 4.65
R30 VPWR.n19 VPWR.n18 4.095
R31 VPWR.n3 VPWR.n2 1.406
R32 VPWR.n4 VPWR.n1 0.233
R33 VPWR.n19 VPWR.n16 0.133
R34 VPWR VPWR.n19 0.127
R35 VPWR.n6 VPWR.n4 0.119
R36 VPWR.n8 VPWR.n6 0.119
R37 VPWR.n10 VPWR.n8 0.119
R38 VPWR.n12 VPWR.n10 0.119
R39 VPWR.n14 VPWR.n12 0.119
R40 VPWR.n16 VPWR.n14 0.119
R41 VPB.t4 VPB.t1 556.386
R42 VPB.t3 VPB.t2 449.844
R43 VPB.t2 VPB.t6 331.464
R44 VPB VPB.t9 263.395
R45 VPB.t6 VPB.t7 248.598
R46 VPB.t0 VPB.t3 248.598
R47 VPB.t1 VPB.t0 248.598
R48 VPB.t5 VPB.t4 248.598
R49 VPB.t8 VPB.t5 248.598
R50 VPB.t9 VPB.t8 248.598
R51 VGND.n9 VGND.n8 106.463
R52 VGND.n14 VGND.n13 106.463
R53 VGND.n1 VGND.n0 92.5
R54 VGND.n3 VGND.n2 92.5
R55 VGND.n0 VGND.t0 34.153
R56 VGND.n2 VGND.t1 34.153
R57 VGND.n8 VGND.t2 24.923
R58 VGND.n8 VGND.t3 24.923
R59 VGND.n13 VGND.t5 24.923
R60 VGND.n13 VGND.t4 24.923
R61 VGND.n5 VGND.n1 6.437
R62 VGND.n5 VGND.n4 4.65
R63 VGND.n7 VGND.n6 4.65
R64 VGND.n10 VGND.n9 4.65
R65 VGND.n12 VGND.n11 4.65
R66 VGND.n15 VGND.n14 4.115
R67 VGND.n4 VGND.n3 0.449
R68 VGND.n15 VGND.n12 0.133
R69 VGND VGND.n15 0.128
R70 VGND.n7 VGND.n5 0.119
R71 VGND.n10 VGND.n7 0.119
R72 VGND.n12 VGND.n10 0.119
R73 a_55_47.n3 a_55_47.t3 224.961
R74 a_55_47.t6 a_55_47.n5 166.16
R75 a_55_47.n5 a_55_47.n0 99.652
R76 a_55_47.n4 a_55_47.n1 99.652
R77 a_55_47.n3 a_55_47.n2 99.652
R78 a_55_47.n4 a_55_47.n3 71.234
R79 a_55_47.n5 a_55_47.n4 46.747
R80 a_55_47.n0 a_55_47.t5 24.923
R81 a_55_47.n0 a_55_47.t7 24.923
R82 a_55_47.n1 a_55_47.t1 24.923
R83 a_55_47.n1 a_55_47.t2 24.923
R84 a_55_47.n2 a_55_47.t4 24.923
R85 a_55_47.n2 a_55_47.t0 24.923
R86 VNB VNB.t8 6755.01
R87 VNB.t3 VNB.t7 4738.46
R88 VNB.t1 VNB.t0 4158.24
R89 VNB.t7 VNB.t6 2030.77
R90 VNB.t4 VNB.t3 2030.77
R91 VNB.t0 VNB.t4 2030.77
R92 VNB.t2 VNB.t1 2030.77
R93 VNB.t5 VNB.t2 2030.77
R94 VNB.t9 VNB.t5 2030.77
R95 VNB.t8 VNB.t9 2030.77
R96 C1.n3 C1.t1 225.289
R97 C1.n2 C1.t2 221.719
R98 C1.n3 C1.t3 149.419
R99 C1.n1 C1.t0 149.419
R100 C1.n5 C1.n4 76
R101 C1.n4 C1.n3 49.985
R102 C1.n4 C1.n2 21.422
R103 C1.n5 C1.n0 16.738
R104 C1.n0 C1 3.692
R105 C1.n2 C1.n1 3.57
R106 C1 C1.n5 2.215
R107 a_729_47.n1 a_729_47.n0 262.913
R108 a_729_47.n0 a_729_47.t3 24.923
R109 a_729_47.n0 a_729_47.t2 24.923
R110 a_729_47.t0 a_729_47.n1 24.923
R111 a_729_47.n1 a_729_47.t1 24.923
R112 Y.n4 Y.t1 421.307
R113 Y.n1 Y.t6 208.443
R114 Y Y.t4 178.391
R115 Y.n5 Y.n3 159.159
R116 Y.n6 Y.n2 153.394
R117 Y.n0 Y.t5 117.423
R118 Y.n6 Y.n5 66.666
R119 Y.n5 Y.n4 41.966
R120 Y.n8 Y.n0 40.464
R121 Y.n2 Y.t7 40.385
R122 Y.n2 Y.t2 40.385
R123 Y.n3 Y.t3 26.595
R124 Y.n3 Y.t0 26.595
R125 Y.n8 Y 11.911
R126 Y Y.n1 5.857
R127 Y.n1 Y 4.908
R128 Y.n0 Y 4.547
R129 Y.n7 Y.n6 3.466
R130 Y.n4 Y 2.7
R131 Y Y.n7 1.422
R132 Y.n7 Y 0.533
R133 Y Y.n8 0.177
R134 A3.n0 A3.t2 232.43
R135 A3.n1 A3.t3 221.719
R136 A3.n4 A3.t1 185.122
R137 A3.n0 A3.t0 149.419
R138 A3.n3 A3.n2 76
R139 A3.n5 A3.n4 76
R140 A3.n2 A3.n0 57.125
R141 A3.n5 A3.n3 16.738
R142 A3.n2 A3.n1 7.14
R143 A3.n3 A3 3.692
R144 A3 A3.n5 2.215
R145 B1.n0 B1.t1 291.341
R146 B1.n2 B1.t3 221.719
R147 B1.n2 B1.t2 160.13
R148 B1.n1 B1.t0 149.419
R149 B1.n0 B1 84.615
R150 B1.n4 B1.n3 76
R151 B1.n3 B1.n1 58.911
R152 B1 B1.n4 14.523
R153 B1.n4 B1 8.123
R154 B1.n3 B1.n2 5.355
R155 B1.n1 B1.n0 1.785
R156 A2.n3 A2.t2 225.289
R157 A2.n0 A2.t1 221.719
R158 A2.n0 A2.t3 152.989
R159 A2.n3 A2.t0 149.419
R160 A2 A2.n4 78.215
R161 A2.n2 A2.n1 76
R162 A2 A2.n2 14.523
R163 A2.n2 A2 8.123
R164 A2.n1 A2.n0 5.355
R165 A2.n4 A2.n3 5.355
R166 a_301_297.n1 a_301_297.n0 378.051
R167 a_301_297.n0 a_301_297.t3 26.595
R168 a_301_297.n0 a_301_297.t2 26.595
R169 a_301_297.t1 a_301_297.n1 26.595
R170 a_301_297.n1 a_301_297.t0 26.595
C0 VPB VPWR 0.12fF
C1 A1 A2 0.10fF
C2 VPWR Y 0.74fF
C3 A3 Y 0.12fF
C4 VPWR VGND 0.13fF
C5 B1 Y 0.29fF
C6 C1 Y 0.33fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__o311ai_4.ext - technology: sky130A

.subckt sky130_fd_sc_hd__o311ai_4 Y C1 B1 A3 A2 A1 VGND VPWR VNB VPB
X0 a_39_297.t3 A1.t0 VPWR.t3 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 Y.t11 C1.t0 VPWR.t7 VPB.t11 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 VPWR.t2 A1.t1 a_39_297.t2 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 VPWR.t11 B1.t0 Y.t7 VPB.t19 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 a_125_47.t3 A3.t0 VGND.t3 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 a_125_47.t7 A1.t2 VGND.t7 VNB.t7 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 a_125_47.t8 A2.t0 VGND.t8 VNB.t8 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 a_1163_47.t3 B1.t1 a_125_47.t12 VNB.t15 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 a_39_297.t1 A1.t3 VPWR.t1 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 a_1163_47.t2 B1.t2 a_125_47.t15 VNB.t14 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 VGND.t2 A3.t1 a_125_47.t2 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 VPWR.t8 C1.t1 Y.t10 VPB.t12 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 VGND.t6 A1.t4 a_125_47.t6 VNB.t6 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 VGND.t1 A3.t2 a_125_47.t1 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14 a_39_297.t6 A2.t1 a_461_297.t7 VPB.t6 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 VGND.t5 A1.t5 a_125_47.t5 VNB.t5 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X16 a_125_47.t14 B1.t3 a_1163_47.t1 VNB.t13 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X17 Y.t9 C1.t2 VPWR.t9 VPB.t13 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X18 a_125_47.t4 A1.t6 VGND.t4 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X19 VGND.t9 A2.t2 a_125_47.t9 VNB.t9 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X20 a_125_47.t13 B1.t4 a_1163_47.t0 VNB.t12 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X21 VGND.t10 A2.t3 a_125_47.t10 VNB.t10 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X22 Y.t15 C1.t3 a_1163_47.t7 VNB.t19 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X23 Y.t14 C1.t4 a_1163_47.t6 VNB.t18 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X24 a_461_297.t6 A2.t4 a_39_297.t7 VPB.t7 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X25 Y.t5 A3.t3 a_461_297.t3 VPB.t17 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X26 VPWR.t10 C1.t5 Y.t8 VPB.t14 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X27 Y.t6 A3.t4 a_461_297.t2 VPB.t18 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X28 Y.t0 B1.t5 VPWR.t4 VPB.t8 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X29 a_125_47.t0 A3.t5 VGND.t0 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X30 VPWR.t0 A1.t7 a_39_297.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X31 a_461_297.t1 A3.t6 Y.t4 VPB.t16 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X32 a_461_297.t0 A3.t7 Y.t3 VPB.t15 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X33 VPWR.t5 B1.t6 Y.t1 VPB.t9 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X34 a_125_47.t11 A2.t5 VGND.t11 VNB.t11 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X35 a_1163_47.t5 C1.t6 Y.t13 VNB.t17 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X36 a_1163_47.t4 C1.t7 Y.t12 VNB.t16 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X37 Y.t2 B1.t7 VPWR.t6 VPB.t10 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X38 a_39_297.t4 A2.t6 a_461_297.t5 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X39 a_461_297.t4 A2.t7 a_39_297.t5 VPB.t5 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
R0 A1.n1 A1.t0 221.719
R1 A1.n3 A1.t1 221.719
R2 A1.n0 A1.t3 221.719
R3 A1.n8 A1.t7 221.719
R4 A1.n1 A1.t5 149.419
R5 A1.n3 A1.t2 149.419
R6 A1.n0 A1.t4 149.419
R7 A1.n8 A1.t6 149.419
R8 A1.n2 A1 80.43
R9 A1.n5 A1.n4 76
R10 A1.n7 A1.n6 76
R11 A1.n10 A1.n9 76
R12 A1.n9 A1.n7 60.696
R13 A1.n4 A1.n0 50.877
R14 A1.n2 A1.n1 38.381
R15 A1.n3 A1.n2 36.596
R16 A1.n4 A1.n3 24.1
R17 A1 A1.n10 22.153
R18 A1.n6 A1 16.246
R19 A1.n5 A1 12.307
R20 A1 A1.n5 10.338
R21 A1.n7 A1.n0 9.818
R22 A1.n6 A1 6.4
R23 A1.n9 A1.n8 4.462
R24 A1.n10 A1 0.492
R25 VPWR.n3 VPWR.n2 166.835
R26 VPWR.n1 VPWR.n0 163.438
R27 VPWR.n7 VPWR.n6 163.438
R28 VPWR.n12 VPWR.n11 163.438
R29 VPWR.n33 VPWR.n32 163.438
R30 VPWR.n38 VPWR.n37 163.438
R31 VPWR.n2 VPWR.t7 26.595
R32 VPWR.n2 VPWR.t8 26.595
R33 VPWR.n0 VPWR.t9 26.595
R34 VPWR.n0 VPWR.t10 26.595
R35 VPWR.n6 VPWR.t4 26.595
R36 VPWR.n6 VPWR.t5 26.595
R37 VPWR.n11 VPWR.t6 26.595
R38 VPWR.n11 VPWR.t11 26.595
R39 VPWR.n32 VPWR.t3 26.595
R40 VPWR.n32 VPWR.t2 26.595
R41 VPWR.n37 VPWR.t1 26.595
R42 VPWR.n37 VPWR.t0 26.595
R43 VPWR.n5 VPWR.n4 4.65
R44 VPWR.n8 VPWR.n7 4.65
R45 VPWR.n10 VPWR.n9 4.65
R46 VPWR.n13 VPWR.n12 4.65
R47 VPWR.n15 VPWR.n14 4.65
R48 VPWR.n17 VPWR.n16 4.65
R49 VPWR.n19 VPWR.n18 4.65
R50 VPWR.n21 VPWR.n20 4.65
R51 VPWR.n23 VPWR.n22 4.65
R52 VPWR.n25 VPWR.n24 4.65
R53 VPWR.n27 VPWR.n26 4.65
R54 VPWR.n29 VPWR.n28 4.65
R55 VPWR.n31 VPWR.n30 4.65
R56 VPWR.n34 VPWR.n33 4.65
R57 VPWR.n36 VPWR.n35 4.65
R58 VPWR.n39 VPWR.n38 4.05
R59 VPWR.n3 VPWR.n1 3.856
R60 VPWR.n5 VPWR.n3 0.258
R61 VPWR.n39 VPWR.n36 0.134
R62 VPWR VPWR.n39 0.131
R63 VPWR.n8 VPWR.n5 0.119
R64 VPWR.n10 VPWR.n8 0.119
R65 VPWR.n13 VPWR.n10 0.119
R66 VPWR.n15 VPWR.n13 0.119
R67 VPWR.n17 VPWR.n15 0.119
R68 VPWR.n19 VPWR.n17 0.119
R69 VPWR.n21 VPWR.n19 0.119
R70 VPWR.n23 VPWR.n21 0.119
R71 VPWR.n25 VPWR.n23 0.119
R72 VPWR.n27 VPWR.n25 0.119
R73 VPWR.n29 VPWR.n27 0.119
R74 VPWR.n31 VPWR.n29 0.119
R75 VPWR.n34 VPWR.n31 0.119
R76 VPWR.n36 VPWR.n34 0.119
R77 a_39_297.n1 a_39_297.t6 472.325
R78 a_39_297.n1 a_39_297.n0 299.276
R79 a_39_297.n3 a_39_297.t0 259.132
R80 a_39_297.n3 a_39_297.n2 159.159
R81 a_39_297.n5 a_39_297.n4 159.158
R82 a_39_297.n4 a_39_297.n1 44.8
R83 a_39_297.n4 a_39_297.n3 44.8
R84 a_39_297.n0 a_39_297.t7 26.595
R85 a_39_297.n0 a_39_297.t4 26.595
R86 a_39_297.n2 a_39_297.t2 26.595
R87 a_39_297.n2 a_39_297.t1 26.595
R88 a_39_297.n5 a_39_297.t5 26.595
R89 a_39_297.t3 a_39_297.n5 26.595
R90 VPB.t6 VPB.t15 556.386
R91 VPB.t17 VPB.t19 260.436
R92 VPB VPB.t0 251.557
R93 VPB.t12 VPB.t11 248.598
R94 VPB.t13 VPB.t12 248.598
R95 VPB.t14 VPB.t13 248.598
R96 VPB.t8 VPB.t14 248.598
R97 VPB.t9 VPB.t8 248.598
R98 VPB.t10 VPB.t9 248.598
R99 VPB.t19 VPB.t10 248.598
R100 VPB.t16 VPB.t17 248.598
R101 VPB.t18 VPB.t16 248.598
R102 VPB.t15 VPB.t18 248.598
R103 VPB.t7 VPB.t6 248.598
R104 VPB.t4 VPB.t7 248.598
R105 VPB.t5 VPB.t4 248.598
R106 VPB.t3 VPB.t5 248.598
R107 VPB.t2 VPB.t3 248.598
R108 VPB.t1 VPB.t2 248.598
R109 VPB.t0 VPB.t1 248.598
R110 C1.n9 C1.t5 228.859
R111 C1.n0 C1.t0 221.719
R112 C1.n4 C1.t1 221.719
R113 C1.n8 C1.t2 221.719
R114 C1.n0 C1.t7 156.559
R115 C1.n9 C1.t3 149.419
R116 C1.n5 C1.t6 149.419
R117 C1.n3 C1.t4 149.419
R118 C1.n2 C1.n1 76
R119 C1.n7 C1.n6 76
R120 C1.n11 C1.n10 76
R121 C1.n2 C1.n0 64.266
R122 C1.n6 C1.n4 49.985
R123 C1.n10 C1.n8 35.703
R124 C1.n10 C1.n9 32.133
R125 C1.n6 C1.n5 17.851
R126 C1.n11 C1.n7 16.738
R127 C1.n1 C1 13.046
R128 C1.n1 C1 9.6
R129 C1.n4 C1.n3 7.14
R130 C1.n7 C1 3.692
R131 C1.n3 C1.n2 3.57
R132 C1 C1.n11 2.215
R133 Y.n9 Y.t3 472.325
R134 Y.n9 Y.n8 299.276
R135 Y.n14 Y.t11 208.328
R136 Y.n13 Y.n4 159.159
R137 Y.n12 Y.n5 159.159
R138 Y.n11 Y.n6 159.159
R139 Y.n10 Y.n7 157.824
R140 Y.n2 Y.n1 139.247
R141 Y.n2 Y.n0 92.5
R142 Y.n11 Y.n10 45.333
R143 Y.n10 Y.n9 45.333
R144 Y.n13 Y.n12 44.8
R145 Y.n12 Y.n11 44.8
R146 Y.n15 Y.n13 40.266
R147 Y.n7 Y.t7 30.535
R148 Y.n4 Y.t10 26.595
R149 Y.n4 Y.t9 26.595
R150 Y.n5 Y.t8 26.595
R151 Y.n5 Y.t0 26.595
R152 Y.n6 Y.t1 26.595
R153 Y.n6 Y.t2 26.595
R154 Y.n7 Y.t5 26.595
R155 Y.n8 Y.t4 26.595
R156 Y.n8 Y.t6 26.595
R157 Y.n0 Y.t12 24.923
R158 Y.n0 Y.t14 24.923
R159 Y.n1 Y.t13 24.923
R160 Y.n1 Y.t15 24.923
R161 Y.n3 Y.n2 20.034
R162 Y Y.n3 13.612
R163 Y Y.n14 6.161
R164 Y.n15 Y 6.063
R165 Y.n14 Y 5.164
R166 Y.n16 Y.n15 4.042
R167 Y.n16 Y 1.625
R168 Y Y.n16 1.347
R169 Y.n3 Y 0.203
R170 B1.n11 B1.t0 228.859
R171 B1.n1 B1.t5 221.719
R172 B1.n2 B1.t6 221.719
R173 B1.n10 B1.t7 221.719
R174 B1.n1 B1.t2 156.559
R175 B1.n11 B1.t3 149.419
R176 B1.n9 B1.t1 149.419
R177 B1.n3 B1.t4 149.419
R178 B1.n5 B1.n4 76
R179 B1.n8 B1.n7 76
R180 B1.n13 B1.n12 76
R181 B1.n8 B1.n0 60.696
R182 B1.n4 B1.n3 50.877
R183 B1.n12 B1.n10 49.092
R184 B1.n12 B1.n11 18.744
R185 B1.n4 B1.n1 16.959
R186 B1.n7 B1.n6 16.738
R187 B1.n13 B1 16.246
R188 B1.n5 B1 11.323
R189 B1 B1.n5 11.323
R190 B1.n3 B1.n2 7.14
R191 B1.n10 B1.n9 7.14
R192 B1 B1.n13 6.4
R193 B1.n6 B1 5.415
R194 B1.n9 B1.n8 4.462
R195 B1.n2 B1.n0 2.677
R196 B1.n7 B1 0.492
R197 A3.n2 A3.t3 277.059
R198 A3.n3 A3.t6 221.719
R199 A3.n7 A3.t4 221.719
R200 A3.n0 A3.t7 221.719
R201 A3.n14 A3.t0 165.485
R202 A3.n13 A3.t2 149.419
R203 A3.n6 A3.t5 149.419
R204 A3.n4 A3.t1 149.419
R205 A3.n2 A3.n1 76
R206 A3.n9 A3.n8 76
R207 A3.n12 A3.n11 76
R208 A3.n15 A3.n14 76
R209 A3.n14 A3.n13 58.911
R210 A3.n5 A3.n0 48.2
R211 A3.n8 A3.n7 33.918
R212 A3.n8 A3.n4 26.777
R213 A3.n3 A3.n2 19.637
R214 A3.n11 A3.n10 16.738
R215 A3 A3.n9 14.523
R216 A3.n4 A3.n3 14.281
R217 A3.n7 A3.n6 14.281
R218 A3.n1 A3 14.03
R219 A3.n15 A3 13.046
R220 A3.n6 A3.n5 12.496
R221 A3.n12 A3.n0 12.496
R222 A3 A3.n15 9.6
R223 A3.n1 A3 8.615
R224 A3.n9 A3 8.123
R225 A3.n11 A3 3.692
R226 A3.n10 A3 2.215
R227 A3.n13 A3.n12 1.785
R228 VGND.n0 VGND.t2 194.325
R229 VGND.n2 VGND.n1 106.463
R230 VGND.n12 VGND.n11 106.463
R231 VGND.n17 VGND.n16 106.463
R232 VGND.n22 VGND.n21 106.463
R233 VGND.n6 VGND.n5 105.665
R234 VGND.n26 VGND.t4 96.068
R235 VGND.n5 VGND.t10 28.615
R236 VGND.n1 VGND.t0 24.923
R237 VGND.n1 VGND.t1 24.923
R238 VGND.n5 VGND.t3 24.923
R239 VGND.n11 VGND.t11 24.923
R240 VGND.n11 VGND.t9 24.923
R241 VGND.n16 VGND.t8 24.923
R242 VGND.n16 VGND.t5 24.923
R243 VGND.n21 VGND.t7 24.923
R244 VGND.n21 VGND.t6 24.923
R245 VGND.n27 VGND.n26 4.65
R246 VGND.n4 VGND.n3 4.65
R247 VGND.n8 VGND.n7 4.65
R248 VGND.n10 VGND.n9 4.65
R249 VGND.n13 VGND.n12 4.65
R250 VGND.n15 VGND.n14 4.65
R251 VGND.n18 VGND.n17 4.65
R252 VGND.n20 VGND.n19 4.65
R253 VGND.n23 VGND.n22 4.65
R254 VGND.n25 VGND.n24 4.65
R255 VGND.n3 VGND.n2 1.882
R256 VGND.n7 VGND.n6 1.882
R257 VGND.n4 VGND.n0 0.569
R258 VGND.n8 VGND.n4 0.119
R259 VGND.n10 VGND.n8 0.119
R260 VGND.n13 VGND.n10 0.119
R261 VGND.n15 VGND.n13 0.119
R262 VGND.n18 VGND.n15 0.119
R263 VGND.n20 VGND.n18 0.119
R264 VGND.n23 VGND.n20 0.119
R265 VGND.n25 VGND.n23 0.119
R266 VGND.n27 VGND.n25 0.119
R267 VGND VGND.n27 0.027
R268 a_125_47.n9 a_125_47.n8 146.399
R269 a_125_47.n3 a_125_47.n1 139.247
R270 a_125_47.n9 a_125_47.n7 99.652
R271 a_125_47.n10 a_125_47.n6 99.652
R272 a_125_47.n11 a_125_47.n5 99.652
R273 a_125_47.n4 a_125_47.n0 99.652
R274 a_125_47.n13 a_125_47.n12 99.652
R275 a_125_47.n3 a_125_47.n2 92.5
R276 a_125_47.n4 a_125_47.n3 77.913
R277 a_125_47.n12 a_125_47.n11 47.86
R278 a_125_47.n12 a_125_47.n4 46.747
R279 a_125_47.n11 a_125_47.n10 46.747
R280 a_125_47.n10 a_125_47.n9 46.747
R281 a_125_47.n2 a_125_47.t12 24.923
R282 a_125_47.n2 a_125_47.t14 24.923
R283 a_125_47.n1 a_125_47.t15 24.923
R284 a_125_47.n1 a_125_47.t13 24.923
R285 a_125_47.n8 a_125_47.t6 24.923
R286 a_125_47.n8 a_125_47.t4 24.923
R287 a_125_47.n7 a_125_47.t5 24.923
R288 a_125_47.n7 a_125_47.t7 24.923
R289 a_125_47.n6 a_125_47.t9 24.923
R290 a_125_47.n6 a_125_47.t8 24.923
R291 a_125_47.n5 a_125_47.t10 24.923
R292 a_125_47.n5 a_125_47.t11 24.923
R293 a_125_47.n0 a_125_47.t2 24.923
R294 a_125_47.n0 a_125_47.t0 24.923
R295 a_125_47.n13 a_125_47.t1 24.923
R296 a_125_47.t3 a_125_47.n13 24.923
R297 VNB VNB.t4 6561.6
R298 VNB.t2 VNB.t13 4738.46
R299 VNB.t10 VNB.t3 2127.47
R300 VNB.t18 VNB.t16 2030.77
R301 VNB.t17 VNB.t18 2030.77
R302 VNB.t19 VNB.t17 2030.77
R303 VNB.t14 VNB.t19 2030.77
R304 VNB.t12 VNB.t14 2030.77
R305 VNB.t15 VNB.t12 2030.77
R306 VNB.t13 VNB.t15 2030.77
R307 VNB.t0 VNB.t2 2030.77
R308 VNB.t1 VNB.t0 2030.77
R309 VNB.t3 VNB.t1 2030.77
R310 VNB.t11 VNB.t10 2030.77
R311 VNB.t9 VNB.t11 2030.77
R312 VNB.t8 VNB.t9 2030.77
R313 VNB.t5 VNB.t8 2030.77
R314 VNB.t7 VNB.t5 2030.77
R315 VNB.t6 VNB.t7 2030.77
R316 VNB.t4 VNB.t6 2030.77
R317 A2.n0 A2.t1 221.719
R318 A2.n2 A2.t4 221.719
R319 A2.n8 A2.t6 221.719
R320 A2.n9 A2.t7 221.719
R321 A2.n0 A2.t3 149.419
R322 A2.n2 A2.t5 149.419
R323 A2.n8 A2.t2 149.419
R324 A2.n9 A2.t0 149.419
R325 A2.n5 A2.n3 76
R326 A2.n7 A2.n6 76
R327 A2.n11 A2.n10 76
R328 A2.n7 A2.n3 60.696
R329 A2.n10 A2.n8 58.911
R330 A2.n2 A2.n1 48.2
R331 A2.n1 A2.n0 26.777
R332 A2 A2.n11 17.476
R333 A2.n5 A2.n4 16.738
R334 A2.n10 A2.n9 16.066
R335 A2.n3 A2.n2 12.496
R336 A2.n6 A2 11.569
R337 A2.n6 A2 11.076
R338 A2 A2.n5 5.661
R339 A2.n11 A2 5.169
R340 A2.n8 A2.n7 1.785
R341 A2.n4 A2 0.246
R342 a_1163_47.n1 a_1163_47.t4 224.961
R343 a_1163_47.n4 a_1163_47.t1 224.961
R344 a_1163_47.n1 a_1163_47.n0 92.5
R345 a_1163_47.n5 a_1163_47.n4 92.5
R346 a_1163_47.n3 a_1163_47.n2 49.971
R347 a_1163_47.n3 a_1163_47.n1 46.747
R348 a_1163_47.n4 a_1163_47.n3 46.747
R349 a_1163_47.n2 a_1163_47.t7 24.923
R350 a_1163_47.n2 a_1163_47.t2 24.923
R351 a_1163_47.n0 a_1163_47.t6 24.923
R352 a_1163_47.n0 a_1163_47.t5 24.923
R353 a_1163_47.n5 a_1163_47.t0 24.923
R354 a_1163_47.t3 a_1163_47.n5 24.923
R355 a_461_297.n2 a_461_297.n0 188.65
R356 a_461_297.n5 a_461_297.n4 188.649
R357 a_461_297.n2 a_461_297.n1 150.25
R358 a_461_297.n4 a_461_297.n3 150.25
R359 a_461_297.n4 a_461_297.n2 77.552
R360 a_461_297.n0 a_461_297.t5 26.595
R361 a_461_297.n0 a_461_297.t4 26.595
R362 a_461_297.n1 a_461_297.t7 26.595
R363 a_461_297.n1 a_461_297.t6 26.595
R364 a_461_297.n3 a_461_297.t2 26.595
R365 a_461_297.n3 a_461_297.t0 26.595
R366 a_461_297.t3 a_461_297.n5 26.595
R367 a_461_297.n5 a_461_297.t1 26.595
C0 C1 Y 0.56fF
C1 C1 B1 0.10fF
C2 VGND A1 0.10fF
C3 VPWR VPB 0.18fF
C4 VPWR Y 1.16fF
C5 Y A3 0.33fF
C6 VPWR VGND 0.20fF
C7 Y B1 0.43fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__o2111a_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__o2111a_1 X D1 C1 B1 A2 A1 VPWR VGND VNB VPB
X0 a_676_297.t1 A2.t0 a_79_21.t4 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_512_47.t0 B1.t0 a_409_47.t1 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 a_306_47.t1 D1.t0 a_79_21.t0 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 VGND.t1 A2.t1 a_512_47.t2 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 VPWR.t4 C1.t0 a_79_21.t1 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 a_79_21.t3 B1.t1 VPWR.t0 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 VPWR.t2 A1.t0 a_676_297.t0 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 a_512_47.t1 A1.t1 VGND.t0 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 a_409_47.t0 C1.t1 a_306_47.t0 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 VPWR.t3 a_79_21.t5 X.t1 VPB.t5 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 a_79_21.t2 D1.t1 VPWR.t1 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 VGND.t2 a_79_21.t6 X.t0 VNB.t5 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
R0 A2.n0 A2.t0 241.437
R1 A2.n0 A2.t1 169.137
R2 A2 A2.n0 83.68
R3  A2 12.142
R4 a_79_21.n3 a_79_21.n2 240.551
R5 a_79_21.n0 a_79_21.t5 234.801
R6 a_79_21.n4 a_79_21.n3 164.215
R7 a_79_21.n0 a_79_21.t6 162.501
R8 a_79_21.n1 a_79_21.t0 117.672
R9 a_79_21.n1 a_79_21.n0 76
R10 a_79_21.n3 a_79_21.n1 73.599
R11 a_79_21.n2 a_79_21.t3 57.13
R12 a_79_21.t1 a_79_21.n4 44.325
R13 a_79_21.n4 a_79_21.t2 41.37
R14 a_79_21.n2 a_79_21.t4 26.595
R15 a_676_297.t0 a_676_297.t1 41.37
R16 VPB.t5 VPB.t1 541.588
R17 VPB.t0 VPB.t2 449.844
R18 VPB.t1 VPB.t0 346.261
R19 VPB.t2 VPB.t4 340.342
R20 VPB.t4 VPB.t3 213.084
R21 VPB VPB.t5 192.367
R22 B1.n0 B1.t1 238.192
R23 B1.n0 B1.t0 165.892
R24 B1.n1 B1.n0 78.133
R25  B1.n1 12.016
R26 B1.n1 B1 4.654
R27 a_409_47.t0 a_409_47.t1 67.384
R28 a_512_47.n0 a_512_47.t1 272.246
R29 a_512_47.t0 a_512_47.n0 87.692
R30 a_512_47.n0 a_512_47.t2 24.923
R31 VNB VNB.t5 6078.09
R32 VNB.t5 VNB.t0 4762.64
R33 VNB.t2 VNB.t4 3674.73
R34 VNB.t1 VNB.t2 2490.11
R35 VNB.t0 VNB.t1 2490.11
R36 VNB.t4 VNB.t3 2030.77
R37 D1.n0 D1.t1 241.437
R38 D1.n0 D1.t0 169.137
R39 D1 D1.n0 80.864
R40  D1 24.783
R41 a_306_47.t0 a_306_47.t1 67.384
R42 VGND.n1 VGND.t2 194.709
R43 VGND.n1 VGND.n0 113.011
R44 VGND.n0 VGND.t0 24.923
R45 VGND.n0 VGND.t1 24.923
R46 VGND VGND.n1 0.144
R47 C1.n0 C1.t0 241.437
R48 C1.n0 C1.t1 169.137
R49 C1 C1.n0 78.607
R50 VPWR.n1 VPWR.t2 195.3
R51 VPWR.n11 VPWR.n10 146.25
R52 VPWR.n7 VPWR.n6 146.25
R53 VPWR.n0 VPWR.t0 60.085
R54 VPWR.n0 VPWR.t4 60.085
R55 VPWR.n10 VPWR.t3 28.565
R56 VPWR.n6 VPWR.t1 27.58
R57 VPWR.n1 VPWR.n0 6.253
R58 VPWR.n9 VPWR.n8 4.65
R59 VPWR.n3 VPWR.n2 4.65
R60 VPWR.n5 VPWR.n4 4.65
R61 VPWR.n12 VPWR.n11 3.995
R62 VPWR.n8 VPWR.n7 0.263
R63 VPWR.n3 VPWR.n1 0.153
R64 VPWR.n12 VPWR.n9 0.136
R65 VPWR VPWR.n12 0.125
R66 VPWR.n5 VPWR.n3 0.119
R67 VPWR.n9 VPWR.n5 0.119
R68 A1.n0 A1.t0 234.211
R69 A1.n0 A1.t1 161.911
R70 A1.n1 A1.n0 76
R71 A1.n1 A1 11.054
R72 A1 A1.n1 2.133
R73 X.n0 X.t1 172.965
R74 X X.t0 157.361
R75 X X.n0 12.564
R76 X.n0 X 4.065
C0 A2 A1 0.13fF
C1 D1 C1 0.19fF
C2 X VPWR 0.14fF
C3 A2 VPWR 0.12fF
C4 C1 B1 0.15fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__o2111a_2.ext - technology: sky130A

.subckt sky130_fd_sc_hd__o2111a_2 D1 C1 A2 A1 B1 X VGND VPWR VNB VPB
X0 VPWR.t2 a_80_21.t5 X.t1 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 X.t0 a_80_21.t6 VPWR.t1 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 a_80_21.t1 D1.t0 VPWR.t4 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 VGND.t2 a_80_21.t7 X.t3 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 VPWR.t3 C1.t0 a_80_21.t0 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 X.t2 a_80_21.t8 VGND.t1 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 a_80_21.t4 B1.t0 VPWR.t5 VPB.t6 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 a_674_297.t0 A2.t0 a_80_21.t3 VPB.t5 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 a_386_47.t1 D1.t1 a_80_21.t2 VNB.t6 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 VPWR.t0 A1.t0 a_674_297.t1 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 a_566_47.t1 B1.t1 a_458_47.t0 VNB.t5 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 VGND.t3 A2.t1 a_566_47.t0 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 a_566_47.t2 A1.t1 VGND.t0 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 a_458_47.t1 C1.t1 a_386_47.t0 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
R0 a_80_21.n1 a_80_21.t5 212.079
R1 a_80_21.n0 a_80_21.t6 212.079
R2 a_80_21.n4 a_80_21.n3 189.221
R3 a_80_21.n5 a_80_21.n4 150.872
R4 a_80_21.n1 a_80_21.t7 139.779
R5 a_80_21.n0 a_80_21.t8 139.779
R6 a_80_21.n2 a_80_21.t2 119.909
R7 a_80_21.n2 a_80_21.n1 106.672
R8 a_80_21.n4 a_80_21.n2 64.276
R9 a_80_21.n1 a_80_21.n0 62.806
R10 a_80_21.n3 a_80_21.t4 39.4
R11 a_80_21.n3 a_80_21.t3 37.43
R12 a_80_21.t0 a_80_21.n5 27.58
R13 a_80_21.n5 a_80_21.t1 27.58
R14 X.n2 X.n1 94.618
R15 X.n3 X.n2 49.497
R16 X.n3 X.n0 43.346
R17 X.n1 X.t1 27.58
R18 X.n1 X.t0 27.58
R19 X.n0 X.t3 25.846
R20 X.n0 X.t2 25.846
R21 X.n2 X 7.252
R22 X X.n3 5.91
R23 VPWR.n1 VPWR.n0 307.239
R24 VPWR.n10 VPWR.n9 292.5
R25 VPWR.n6 VPWR.n5 292.5
R26 VPWR.n15 VPWR.t1 159.042
R27 VPWR.n2 VPWR.t0 156.939
R28 VPWR.n0 VPWR.t3 39.4
R29 VPWR.n0 VPWR.t5 37.43
R30 VPWR.n5 VPWR.t4 27.58
R31 VPWR.n9 VPWR.t2 27.58
R32 VPWR.n4 VPWR.n3 4.65
R33 VPWR.n8 VPWR.n7 4.65
R34 VPWR.n12 VPWR.n11 4.65
R35 VPWR.n14 VPWR.n13 4.65
R36 VPWR.n16 VPWR.n15 4.65
R37 VPWR.n2 VPWR.n1 3.993
R38 VPWR.n7 VPWR.n6 0.839
R39 VPWR.n11 VPWR.n10 0.629
R40 VPWR.n4 VPWR.n2 0.144
R41 VPWR.n8 VPWR.n4 0.119
R42 VPWR.n12 VPWR.n8 0.119
R43 VPWR.n14 VPWR.n12 0.119
R44 VPWR.n16 VPWR.n14 0.119
R45 VPWR VPWR.n16 0.02
R46 VPB.t2 VPB.t4 520.872
R47 VPB.t5 VPB.t0 319.626
R48 VPB.t6 VPB.t5 319.626
R49 VPB.t3 VPB.t6 319.626
R50 VPB.t4 VPB.t3 254.517
R51 VPB.t1 VPB.t2 254.517
R52 VPB VPB.t1 192.367
R53 D1.n0 D1.t0 230.791
R54 D1.n0 D1.t1 158.491
R55 D1.n1 D1.n0 76
R56  D1.n1 11.054
R57 D1.n1 D1 2.133
R58 VGND.n1 VGND.t2 193.465
R59 VGND.n5 VGND.t1 112.988
R60 VGND.n2 VGND.n0 110.769
R61 VGND.n0 VGND.t0 38.769
R62 VGND.n0 VGND.t3 33.23
R63 VGND.n6 VGND.n5 4.65
R64 VGND.n4 VGND.n3 4.65
R65 VGND.n2 VGND.n1 3.984
R66 VGND.n4 VGND.n2 0.138
R67 VGND.n6 VGND.n4 0.119
R68 VGND VGND.n6 0.02
R69 VNB VNB.t1 6078.09
R70 VNB.t2 VNB.t6 4593.41
R71 VNB.t4 VNB.t0 2610.99
R72 VNB.t5 VNB.t4 2610.99
R73 VNB.t3 VNB.t5 2610.99
R74 VNB.t1 VNB.t2 2079.12
R75 VNB.t6 VNB.t3 1740.66
R76 C1.n0 C1.t0 241.437
R77 C1.n0 C1.t1 169.137
R78 C1.n1 C1.n0 76
R79  C1 11.303
R80 C1.n1  9.475
R81  C1.n1 1.828
R82 B1.n0 B1.t0 241.437
R83 B1.n0 B1.t1 169.137
R84 B1.n1 B1.n0 76
R85  B1.n1 8.685
R86 B1.n1 B1 1.676
R87 A2.n0 A2.t0 241.437
R88 A2.n0 A2.t1 169.137
R89 A2.n1 A2.n0 76
R90 A2.n1 A2 41.176
R91 A2 A2.n1 1.955
R92 a_674_297.t0 a_674_297.t1 76.83
R93 a_386_47.t0 a_386_47.t1 38.769
R94 A1.n0 A1.t0 236.02
R95 A1.n0 A1.t1 163.72
R96 A1.n1 A1.n0 76
R97 A1  12.246
R98 A1 A1.n1 10.735
R99 A1.n1 A1 8.258
R100 a_458_47.t0 a_458_47.t1 72
R101 a_566_47.n0 a_566_47.t2 181.557
R102 a_566_47.n0 a_566_47.t1 36.923
R103 a_566_47.t0 a_566_47.n0 35.076
C0 X VGND 0.18fF
C1 A2 A1 0.10fF
C2 D1 C1 0.15fF
C3 VPWR X 0.26fF
C4 A2 VPWR 0.15fF
C5 B1 A2 0.11fF
C6 VPWR VGND 0.12fF
C7 A1 VPWR 0.18fF
C8 C1 B1 0.10fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__o2111a_4.ext - technology: sky130A

.subckt sky130_fd_sc_hd__o2111a_4 X A1 A2 C1 B1 D1 VPWR VGND VNB VPB
X0 VGND.t7 A1.t0 a_361_47.t5 VNB.t13 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 X.t7 a_27_297.t10 VPWR.t3 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 a_27_297.t1 A2.t0 a_852_297.t0 VPB.t5 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 VPWR.t2 a_27_297.t11 X.t6 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 VGND.t2 a_27_297.t12 X.t3 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 VPWR.t6 B1.t0 a_27_297.t4 VPB.t8 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 a_852_297.t1 A1.t1 VPWR.t11 VPB.t13 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 a_27_297.t5 B1.t1 VPWR.t7 VPB.t9 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 a_361_47.t4 A1.t2 VGND.t6 VNB.t12 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 VPWR.t4 C1.t0 a_27_297.t2 VPB.t6 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 VGND.t0 A2.t1 a_361_47.t0 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 a_27_297.t6 D1.t0 VPWR.t8 VPB.t10 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 X.t2 a_27_297.t13 VGND.t3 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 X.t5 a_27_297.t14 VPWR.t1 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14 a_27_47.t3 D1.t1 a_27_297.t7 VNB.t10 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X15 a_361_47.t2 B1.t2 a_277_47.t0 VNB.t8 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X16 a_361_47.t1 A2.t2 VGND.t1 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X17 a_277_47.t1 C1.t1 a_27_47.t1 VNB.t6 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X18 a_445_47.t0 B1.t3 a_361_47.t3 VNB.t9 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X19 X.t1 a_27_297.t15 VGND.t4 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X20 a_27_297.t3 C1.t2 VPWR.t5 VPB.t7 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X21 a_681_297.t0 A2.t3 a_27_297.t0 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X22 a_27_47.t0 C1.t3 a_445_47.t1 VNB.t7 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X23 VGND.t5 a_27_297.t16 X.t0 VNB.t5 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X24 VPWR.t9 D1.t2 a_27_297.t8 VPB.t11 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X25 VPWR.t0 a_27_297.t17 X.t4 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X26 VPWR.t10 A1.t3 a_681_297.t1 VPB.t12 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X27 a_27_297.t9 D1.t3 a_27_47.t2 VNB.t11 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
R0 A1.n0 A1.t3 218.076
R1 A1.n0 A1.t1 194.781
R2 A1.n1 A1.t2 171.912
R3 A1.n1 A1.t0 145.955
R4 A1 A1.n2 89.744
R5 A1.n2 A1.n0 21.283
R6 A1.n2 A1.n1 12.519
R7 a_361_47.n2 a_361_47.n1 192.022
R8 a_361_47.n3 a_361_47.n2 95.465
R9 a_361_47.n2 a_361_47.n0 49.159
R10 a_361_47.t0 a_361_47.n3 34.153
R11 a_361_47.n3 a_361_47.t4 34.153
R12 a_361_47.n0 a_361_47.t1 33.23
R13 a_361_47.n1 a_361_47.t3 24.923
R14 a_361_47.n1 a_361_47.t2 24.923
R15 a_361_47.n0 a_361_47.t5 24.923
R16 VGND.n16 VGND.t1 190.315
R17 VGND.n2 VGND.t5 187.062
R18 VGND.n6 VGND.n5 110.854
R19 VGND.n1 VGND.n0 107.86
R20 VGND.n11 VGND.n10 105.645
R21 VGND.n5 VGND.t3 48
R22 VGND.n5 VGND.t0 34.153
R23 VGND.n0 VGND.t2 26.769
R24 VGND.n0 VGND.t4 25.846
R25 VGND.n10 VGND.t6 24.923
R26 VGND.n10 VGND.t7 24.923
R27 VGND.n4 VGND.n3 4.65
R28 VGND.n7 VGND.n6 4.65
R29 VGND.n9 VGND.n8 4.65
R30 VGND.n13 VGND.n12 4.65
R31 VGND.n15 VGND.n14 4.65
R32 VGND.n18 VGND.n17 4.65
R33 VGND.n2 VGND.n1 3.812
R34 VGND.n17 VGND.n16 0.752
R35 VGND VGND.n19 0.725
R36 VGND.n12 VGND.n11 0.376
R37 VGND.n4 VGND.n2 0.257
R38 VGND.n19 VGND.n18 0.134
R39 VGND.n7 VGND.n4 0.119
R40 VGND.n9 VGND.n7 0.119
R41 VGND.n13 VGND.n9 0.119
R42 VGND.n15 VGND.n13 0.119
R43 VGND.n18 VGND.n15 0.119
R44 VNB VNB.t11 6078.09
R45 VNB.t7 VNB.t1 4714.29
R46 VNB.t0 VNB.t3 2876.92
R47 VNB.t12 VNB.t0 2514.28
R48 VNB.t3 VNB.t2 2441.76
R49 VNB.t1 VNB.t13 2248.35
R50 VNB.t4 VNB.t5 2151.65
R51 VNB.t2 VNB.t4 2103.3
R52 VNB.t13 VNB.t12 2030.77
R53 VNB.t8 VNB.t9 2030.77
R54 VNB.t6 VNB.t8 2030.77
R55 VNB.t10 VNB.t6 2030.77
R56 VNB.t11 VNB.t10 2030.77
R57 VNB.t9 VNB.t7 1740.66
R58 a_27_297.n19 a_27_297.n18 313.926
R59 a_27_297.n0 a_27_297.t17 225.289
R60 a_27_297.n2 a_27_297.t10 221.719
R61 a_27_297.n6 a_27_297.t11 221.719
R62 a_27_297.n10 a_27_297.t14 221.719
R63 a_27_297.n15 a_27_297.t8 191.984
R64 a_27_297.n13 a_27_297.t1 178.49
R65 a_27_297.n11 a_27_297.t13 165.485
R66 a_27_297.n17 a_27_297.n16 153.821
R67 a_27_297.n7 a_27_297.t12 149.419
R68 a_27_297.n3 a_27_297.t15 149.419
R69 a_27_297.n0 a_27_297.t16 149.419
R70 a_27_297.n23 a_27_297.n21 146.25
R71 a_27_297.n15 a_27_297.n14 135.352
R72 a_27_297.n21 a_27_297.n13 112.307
R73 a_27_297.n5 a_27_297.n1 93.763
R74 a_27_297.n12 a_27_297.n11 76
R75 a_27_297.n5 a_27_297.n4 76
R76 a_27_297.n9 a_27_297.n8 76
R77 a_27_297.n13 a_27_297.n12 74.263
R78 a_27_297.n23 a_27_297.n22 66.98
R79 a_27_297.n20 a_27_297.n19 50.718
R80 a_27_297.n1 a_27_297.n0 49.092
R81 a_27_297.n19 a_27_297.n17 41.325
R82 a_27_297.n4 a_27_297.n3 30.348
R83 a_27_297.n16 a_27_297.t2 26.595
R84 a_27_297.n16 a_27_297.t6 26.595
R85 a_27_297.n18 a_27_297.t4 26.595
R86 a_27_297.n18 a_27_297.t5 26.595
R87 a_27_297.t0 a_27_297.n23 26.595
R88 a_27_297.n22 a_27_297.t3 26.595
R89 a_27_297.n14 a_27_297.t7 24.923
R90 a_27_297.n14 a_27_297.t9 24.923
R91 a_27_297.n9 a_27_297.n5 17.763
R92 a_27_297.n12 a_27_297.n9 17.763
R93 a_27_297.n8 a_27_297.n7 13.388
R94 a_27_297.n17 a_27_297.n15 11.337
R95 a_27_297.n7 a_27_297.n6 10.711
R96 a_27_297.n11 a_27_297.n10 9.818
R97 a_27_297.n3 a_27_297.n2 8.033
R98 a_27_297.n21 a_27_297.n20 6.853
R99 VPWR.n5 VPWR.t1 575.785
R100 VPWR.n25 VPWR.n24 312.98
R101 VPWR.n30 VPWR.n29 307.239
R102 VPWR.n12 VPWR.n11 306.463
R103 VPWR.n19 VPWR.n18 306.463
R104 VPWR.n2 VPWR.t0 195.051
R105 VPWR.n1 VPWR.n0 164.774
R106 VPWR.n11 VPWR.t11 27.58
R107 VPWR.n11 VPWR.t10 27.58
R108 VPWR.n0 VPWR.t3 26.595
R109 VPWR.n0 VPWR.t2 26.595
R110 VPWR.n18 VPWR.t5 26.595
R111 VPWR.n18 VPWR.t6 26.595
R112 VPWR.n24 VPWR.t7 26.595
R113 VPWR.n24 VPWR.t4 26.595
R114 VPWR.n29 VPWR.t8 26.595
R115 VPWR.n29 VPWR.t9 26.595
R116 VPWR.n4 VPWR.n3 4.65
R117 VPWR.n6 VPWR.n5 4.65
R118 VPWR.n8 VPWR.n7 4.65
R119 VPWR.n10 VPWR.n9 4.65
R120 VPWR.n13 VPWR.n12 4.65
R121 VPWR.n15 VPWR.n14 4.65
R122 VPWR.n17 VPWR.n16 4.65
R123 VPWR.n21 VPWR.n20 4.65
R124 VPWR.n23 VPWR.n22 4.65
R125 VPWR.n26 VPWR.n25 4.65
R126 VPWR.n28 VPWR.n27 4.65
R127 VPWR.n31 VPWR.n30 3.932
R128 VPWR.n2 VPWR.n1 3.733
R129 VPWR.n20 VPWR.n19 0.376
R130 VPWR.n4 VPWR.n2 0.262
R131 VPWR.n31 VPWR.n28 0.137
R132 VPWR VPWR.n31 0.123
R133 VPWR.n6 VPWR.n4 0.119
R134 VPWR.n8 VPWR.n6 0.119
R135 VPWR.n10 VPWR.n8 0.119
R136 VPWR.n13 VPWR.n10 0.119
R137 VPWR.n15 VPWR.n13 0.119
R138 VPWR.n17 VPWR.n15 0.119
R139 VPWR.n21 VPWR.n17 0.119
R140 VPWR.n23 VPWR.n21 0.119
R141 VPWR.n26 VPWR.n23 0.119
R142 VPWR.n28 VPWR.n26 0.119
R143 X.n5 X.n3 230.688
R144 X.n5 X.n4 177.361
R145 X.n2 X.n0 163.427
R146 X.n2 X.n1 115.54
R147 X.n0 X.t2 40.615
R148 X.n1 X.t0 28.615
R149 X.n3 X.t6 26.595
R150 X.n3 X.t5 26.595
R151 X.n4 X.t4 26.595
R152 X.n4 X.t7 26.595
R153 X.n1 X.t1 25.846
R154 X.n0 X.t3 24.923
R155 X X.n5 23.717
R156 X.n6 X.n2 19.576
R157 X.n6 X 15.407
R158 X X.n6 0.711
R159 VPB.t5 VPB.t1 556.386
R160 VPB.t7 VPB.t4 449.844
R161 VPB.t13 VPB.t5 298.909
R162 VPB.t12 VPB.t13 254.517
R163 VPB.t4 VPB.t12 251.557
R164 VPB.t3 VPB.t0 248.598
R165 VPB.t2 VPB.t3 248.598
R166 VPB.t1 VPB.t2 248.598
R167 VPB.t8 VPB.t7 248.598
R168 VPB.t9 VPB.t8 248.598
R169 VPB.t6 VPB.t9 248.598
R170 VPB.t10 VPB.t6 248.598
R171 VPB.t11 VPB.t10 248.598
R172 VPB VPB.t11 192.367
R173 A2.n1 A2.t3 242.053
R174 A2.n0 A2.t0 234.009
R175  A2.n0 186.481
R176 A2.n0 A2.t1 169.137
R177 A2.n1 A2.t2 160.355
R178 A2.n2 A2.n1 76.261
R179  A2.n2 10.847
R180 A2.n2 A2 3.905
R181 a_852_297.t0 a_852_297.t1 69.935
R182 B1.n0 B1.t0 221.719
R183 B1.n1 B1.t1 221.719
R184 B1.n0 B1.t3 149.419
R185 B1.n1 B1.t2 149.419
R186 B1 B1.n2 77.6
R187 B1.n2 B1.n0 37.488
R188 B1.n2 B1.n1 37.488
R189 C1.n1 C1.t2 645.107
R190 C1.n0 C1.t0 241.534
R191  C1.n0 184.478
R192 C1.n0 C1.t1 169.234
R193 C1.n1 C1.t3 164.359
R194 C1.n2 C1.n1 76
R195  C1.n2 12.902
R196 C1.n2 C1 1.877
R197 D1.n1 D1.t2 230.791
R198 D1.n0 D1.t0 221.719
R199 D1.n1 D1.t3 158.491
R200 D1.n0 D1.t1 149.419
R201 D1.n2 D1.n1 76
R202 D1.n1 D1.n0 61.588
R203  D1.n2 16.581
R204 D1.n2 D1 3.2
R205 a_27_47.n1 a_27_47.t0 265.732
R206 a_27_47.t2 a_27_47.n1 201.04
R207 a_27_47.n1 a_27_47.n0 92.5
R208 a_27_47.n0 a_27_47.t1 24.923
R209 a_27_47.n0 a_27_47.t3 24.923
R210 a_277_47.t0 a_277_47.t1 49.846
R211 a_445_47.t0 a_445_47.t1 38.769
R212 a_681_297.t0 a_681_297.t1 54.175
C0 X VGND 0.36fF
C1 A2 A1 0.27fF
C2 VPB VPWR 0.15fF
C3 VPWR X 0.54fF
C4 VPWR VGND 0.16fF
C5 C1 B1 0.29fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__o2111ai_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__o2111ai_1 D1 C1 A2 A1 B1 Y VGND VPWR VNB VPB
X0 VPWR.t3 C1.t0 Y.t4 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_235_47.t1 C1.t1 a_163_47.t1 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 a_343_47.t1 B1.t0 a_235_47.t0 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 Y.t0 B1.t1 VPWR.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 a_454_297.t0 A2.t0 Y.t2 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 Y.t1 D1.t0 VPWR.t1 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 VPWR.t2 A1.t0 a_454_297.t1 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 a_163_47.t0 D1.t1 Y.t3 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 VGND.t0 A2.t1 a_343_47.t0 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 a_343_47.t2 A1.t1 VGND.t1 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
R0 C1.n0 C1.t0 241.437
R1 C1.n0 C1.t1 169.137
R2 C1.n1 C1.n0 76
R3 C1.n1 C1 28.509
R4  C1.n1 11.054
R5 Y.n2 Y.n0 195.985
R6 Y.n2 Y.n1 149.636
R7 Y.n3 Y.t3 83.186
R8 Y.n4 Y.n3 56.504
R9 Y.n0 Y.t0 42.355
R10 Y.n0 Y.t2 37.43
R11 Y.n4 Y.n2 37.052
R12 Y.n1 Y.t4 27.58
R13 Y.n1 Y.t1 27.58
R14 Y.n3 Y 3.186
R15  Y.n4 2.933
R16 VPWR.n7 VPWR.t1 571.144
R17 VPWR.n2 VPWR.n1 307.239
R18 VPWR.n0 VPWR.t2 197.073
R19 VPWR.n1 VPWR.t3 39.4
R20 VPWR.n1 VPWR.t0 37.43
R21 VPWR.n8 VPWR.n7 9.167
R22 VPWR.n6 VPWR.n5 4.65
R23 VPWR.n4 VPWR.n3 4.65
R24 VPWR.n3 VPWR.n2 4.517
R25 VPWR.n4 VPWR.n0 0.143
R26 VPWR.n6 VPWR.n4 0.119
R27 VPWR.n8 VPWR.n6 0.119
R28 VPWR VPWR.n8 0.022
R29 VPB.t0 VPB.t2 328.504
R30 VPB.t2 VPB.t3 319.626
R31 VPB.t4 VPB.t0 319.626
R32 VPB VPB.t1 310.747
R33 VPB.t1 VPB.t4 254.517
R34 a_163_47.t0 a_163_47.t1 38.769
R35 a_235_47.t0 a_235_47.t1 72
R36 VNB VNB.t2 8531.38
R37 VNB.t0 VNB.t1 2683.52
R38 VNB.t1 VNB.t3 2610.99
R39 VNB.t4 VNB.t0 2610.99
R40 VNB.t2 VNB.t4 1740.66
R41 B1.n0 B1.t1 241.437
R42 B1.n0 B1.t0 169.137
R43 B1.n1 B1.n0 76
R44  B1.n1 12.579
R45 B1.n1 B1 2.427
R46 a_343_47.n0 a_343_47.t2 181.428
R47 a_343_47.n0 a_343_47.t1 39.692
R48 a_343_47.t0 a_343_47.n0 35.076
R49 A2.n0 A2.t0 241.437
R50 A2.n0 A2.t1 169.137
R51 A2.n1 A2.n0 76
R52  A2.n1 5.79
R53 A2.n1 A2 1.117
R54 a_454_297.t0 a_454_297.t1 76.83
R55 D1.n0 D1.t0 241.437
R56 D1.n0 D1.t1 169.137
R57 D1.n1 D1.n0 76
R58  D1.n1 11.054
R59 D1.n1 D1 2.133
R60 A1.n0 A1.t0 233.866
R61 A1.n0 A1.t1 161.566
R62 A1 A1.n0 78.133
R63 VGND VGND.n0 110.826
R64 VGND.n0 VGND.t1 38.769
R65 VGND.n0 VGND.t0 33.23
C0 C1 B1 0.15fF
C1 Y C1 0.12fF
C2 A2 A1 0.15fF
C3 Y VPWR 0.39fF
C4 D1 C1 0.14fF
C5 A2 VPWR 0.15fF
C6 B1 A2 0.15fF
C7 Y D1 0.21fF
C8 Y VGND 0.12fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__o2111ai_2.ext - technology: sky130A

.subckt sky130_fd_sc_hd__o2111ai_2 A1 A2 B1 C1 D1 Y VPWR VGND VNB VPB
X0 Y.t8 C1.t0 VPWR.t6 VPB.t8 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_298_47.t1 C1.t1 a_27_47.t3 VNB.t5 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 VGND.t1 A1.t0 a_497_47.t1 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 a_664_297.t3 A1.t1 VPWR.t2 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 VGND.t2 A2.t0 a_497_47.t4 VNB.t8 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 VPWR.t5 C1.t2 Y.t7 VPB.t7 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 a_298_47.t2 B1.t0 a_497_47.t2 VNB.t6 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 a_497_47.t5 A2.t1 VGND.t3 VNB.t9 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 Y.t0 D1.t0 a_27_47.t0 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 a_497_47.t3 B1.t1 a_298_47.t3 VNB.t7 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 Y.t5 B1.t2 VPWR.t3 VPB.t5 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 Y.t3 A2.t2 a_664_297.t0 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 a_27_47.t2 C1.t3 a_298_47.t0 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 VPWR.t0 D1.t1 Y.t1 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14 VPWR.t4 B1.t3 Y.t6 VPB.t6 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 a_27_47.t1 D1.t2 Y.t2 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X16 a_497_47.t0 A1.t2 VGND.t0 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X17 Y.t9 D1.t3 VPWR.t7 VPB.t9 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X18 VPWR.t1 A1.t3 a_664_297.t2 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X19 a_664_297.t1 A2.t3 Y.t4 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
R0 C1.n0 C1.t2 221.719
R1 C1.n1 C1.t0 221.719
R2 C1.n0 C1.t3 149.419
R3 C1.n1 C1.t1 149.419
R4 C1 C1.n2 81.12
R5 C1.n2 C1.n0 39.274
R6 C1.n2 C1.n1 37.488
R7  C1 23.552
R8 VPWR.n15 VPWR.t7 200.936
R9 VPWR.n1 VPWR.t4 191.794
R10 VPWR.n2 VPWR.n0 171.994
R11 VPWR.n11 VPWR.n10 164.214
R12 VPWR.n6 VPWR.n5 164.214
R13 VPWR.n10 VPWR.t6 27.58
R14 VPWR.n10 VPWR.t0 27.58
R15 VPWR.n5 VPWR.t3 27.58
R16 VPWR.n5 VPWR.t5 27.58
R17 VPWR.n0 VPWR.t2 27.58
R18 VPWR.n0 VPWR.t1 27.58
R19 VPWR.n4 VPWR.n3 4.65
R20 VPWR.n7 VPWR.n6 4.65
R21 VPWR.n9 VPWR.n8 4.65
R22 VPWR.n12 VPWR.n11 4.65
R23 VPWR.n14 VPWR.n13 4.65
R24 VPWR.n16 VPWR.n15 4.65
R25 VPWR.n2 VPWR.n1 4.039
R26 VPWR.n4 VPWR.n2 0.137
R27 VPWR.n7 VPWR.n4 0.119
R28 VPWR.n9 VPWR.n7 0.119
R29 VPWR.n12 VPWR.n9 0.119
R30 VPWR.n14 VPWR.n12 0.119
R31 VPWR.n16 VPWR.n14 0.119
R32 VPWR VPWR.n16 0.022
R33 Y.n4 Y.n2 407.421
R34 Y.n4 Y.n3 172.76
R35 Y.n6 Y.n5 171.384
R36 Y.n1 Y.n0 144.889
R37 Y Y.n7 95.699
R38 Y.n6 Y.n4 50.447
R39 Y.n8 Y.n6 50.447
R40 Y.n0 Y.t1 27.58
R41 Y.n0 Y.t9 27.58
R42 Y.n2 Y.t4 27.58
R43 Y.n2 Y.t3 27.58
R44 Y.n3 Y.t6 27.58
R45 Y.n3 Y.t5 27.58
R46 Y.n5 Y.t7 27.58
R47 Y.n5 Y.t8 27.58
R48 Y.n7 Y.t2 25.846
R49 Y.n7 Y.t0 25.846
R50 Y Y.n8 10.092
R51 Y Y.n1 9.331
R52 Y.n1 Y 7.072
R53 Y.n8 Y 6.646
R54 VPB.t6 VPB.t1 583.021
R55 VPB.t3 VPB.t4 254.517
R56 VPB.t2 VPB.t3 254.517
R57 VPB.t1 VPB.t2 254.517
R58 VPB.t5 VPB.t6 254.517
R59 VPB.t7 VPB.t5 254.517
R60 VPB.t8 VPB.t7 254.517
R61 VPB.t0 VPB.t8 254.517
R62 VPB.t9 VPB.t0 254.517
R63 VPB VPB.t9 242.679
R64 a_27_47.n1 a_27_47.t2 192.189
R65 a_27_47.t0 a_27_47.n1 141.81
R66 a_27_47.n1 a_27_47.n0 92.5
R67 a_27_47.n0 a_27_47.t1 26.769
R68 a_27_47.n0 a_27_47.t3 24.923
R69 a_298_47.n1 a_298_47.n0 307.918
R70 a_298_47.t1 a_298_47.n1 26.769
R71 a_298_47.n0 a_298_47.t3 25.846
R72 a_298_47.n0 a_298_47.t2 25.846
R73 a_298_47.n1 a_298_47.t0 24.923
R74 VNB VNB.t0 6489.08
R75 VNB.t4 VNB.t6 4762.64
R76 VNB.t2 VNB.t3 2079.12
R77 VNB.t9 VNB.t2 2079.12
R78 VNB.t8 VNB.t9 2079.12
R79 VNB.t7 VNB.t8 2079.12
R80 VNB.t6 VNB.t7 2079.12
R81 VNB.t5 VNB.t4 2079.12
R82 VNB.t1 VNB.t5 2079.12
R83 VNB.t0 VNB.t1 2079.12
R84 A1.n0 A1.t1 221.719
R85 A1.n1 A1.t3 221.719
R86 A1.n0 A1.t2 149.419
R87 A1.n1 A1.t0 149.419
R88 A1.n3 A1.n2 76
R89 A1.n2 A1.n1 44.629
R90 A1.n2 A1.n0 32.133
R91 A1.n3 A1 20.736
R92 A1 A1.n3 2.816
R93 a_497_47.n2 a_497_47.t2 227.854
R94 a_497_47.t0 a_497_47.n3 187.263
R95 a_497_47.n3 a_497_47.n0 97.552
R96 a_497_47.n2 a_497_47.n1 92.5
R97 a_497_47.n3 a_497_47.n2 55.45
R98 a_497_47.n1 a_497_47.t4 26.769
R99 a_497_47.n0 a_497_47.t1 25.846
R100 a_497_47.n0 a_497_47.t5 25.846
R101 a_497_47.n1 a_497_47.t3 24.923
R102 VGND.n2 VGND.n0 110.945
R103 VGND.n2 VGND.n1 110.741
R104 VGND.n0 VGND.t0 25.846
R105 VGND.n0 VGND.t1 25.846
R106 VGND.n1 VGND.t3 25.846
R107 VGND.n1 VGND.t2 25.846
R108 VGND VGND.n2 1.072
R109 a_664_297.n0 a_664_297.t3 296.74
R110 a_664_297.n0 a_664_297.t0 240.086
R111 a_664_297.n1 a_664_297.n0 90.497
R112 a_664_297.t2 a_664_297.n1 27.58
R113 a_664_297.n1 a_664_297.t1 27.58
R114 A2.n0 A2.t3 221.719
R115 A2.n1 A2.t2 221.719
R116 A2.n0 A2.t1 149.419
R117 A2.n1 A2.t0 149.419
R118 A2.n3 A2.n2 76
R119 A2.n2 A2.n1 40.166
R120 A2.n2 A2.n0 36.596
R121 A2  23.552
R122  A2.n3 18.944
R123 A2.n3 A2 4.608
R124 B1.n3 B1.t2 237.785
R125 B1.n2 B1.t3 221.719
R126 B1.n0 B1.t1 192.263
R127 B1.n1 B1.t0 149.419
R128 B1 B1.n0 81.888
R129 B1 B1.n3 80.096
R130 B1.n3 B1.n2 60.696
R131 B1.n1 B1.n0 33.918
R132 B1.n2 B1.n1 22.314
R133 D1.n0 D1.t1 212.079
R134 D1.n1 D1.t3 212.079
R135 D1.n0 D1.t2 139.779
R136 D1.n1 D1.t0 139.779
R137 D1 D1.n1 124.344
R138 D1.n1 D1.n0 62.806
C0 B1 Y 0.25fF
C1 VPWR VGND 0.12fF
C2 A2 Y 0.11fF
C3 C1 Y 0.23fF
C4 VPB VPWR 0.11fF
C5 VPWR Y 0.92fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__o2111ai_4.ext - technology: sky130A

.subckt sky130_fd_sc_hd__o2111ai_4 A1 A2 B1 C1 D1 Y VGND VPWR VNB VPB
X0 a_27_47.t3 C1.t0 a_445_47.t3 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 a_803_47.t7 A2.t0 VGND.t6 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 a_27_47.t2 C1.t1 a_445_47.t2 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 VGND.t5 A2.t1 a_803_47.t6 VNB.t5 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 a_1163_297.t7 A2.t2 Y.t13 VPB.t15 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 VPWR.t3 C1.t2 Y.t3 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 VGND.t4 A2.t3 a_803_47.t5 VNB.t6 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 Y.t4 D1.t0 VPWR.t8 VPB.t8 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 Y.t12 A2.t4 a_1163_297.t6 VPB.t14 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 a_1163_297.t5 A2.t5 Y.t15 VPB.t13 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 a_445_47.t4 B1.t0 a_803_47.t8 VNB.t16 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 VPWR.t9 D1.t1 Y.t5 VPB.t9 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 a_445_47.t5 B1.t1 a_803_47.t9 VNB.t17 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 Y.t6 D1.t2 VPWR.t10 VPB.t10 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14 VPWR.t6 A1.t0 a_1163_297.t2 VPB.t6 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 a_27_47.t4 D1.t3 Y.t7 VNB.t12 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X16 a_27_47.t5 D1.t4 Y.t8 VNB.t13 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X17 VGND.t3 A1.t1 a_803_47.t3 VNB.t11 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X18 VPWR.t12 B1.t2 Y.t16 VPB.t16 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X19 Y.t17 B1.t3 VPWR.t13 VPB.t17 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X20 a_1163_297.t3 A1.t2 VPWR.t7 VPB.t7 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X21 a_803_47.t10 B1.t4 a_445_47.t6 VNB.t18 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X22 Y.t18 B1.t5 VPWR.t14 VPB.t18 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X23 Y.t2 C1.t3 VPWR.t2 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X24 VPWR.t4 A1.t3 a_1163_297.t0 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X25 a_803_47.t11 B1.t6 a_445_47.t7 VNB.t19 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X26 Y.t9 D1.t5 a_27_47.t6 VNB.t14 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X27 VPWR.t15 B1.t7 Y.t19 VPB.t19 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X28 a_445_47.t1 C1.t4 a_27_47.t1 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X29 a_803_47.t0 A1.t4 VGND.t0 VNB.t8 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X30 VPWR.t1 C1.t5 Y.t1 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X31 a_1163_297.t1 A1.t5 VPWR.t5 VPB.t5 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X32 Y.t14 A2.t6 a_1163_297.t4 VPB.t12 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X33 a_445_47.t0 C1.t6 a_27_47.t0 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X34 a_803_47.t1 A1.t6 VGND.t1 VNB.t9 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X35 Y.t0 C1.t7 VPWR.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X36 a_803_47.t4 A2.t7 VGND.t7 VNB.t7 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X37 VPWR.t11 D1.t6 Y.t10 VPB.t11 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X38 Y.t11 D1.t7 a_27_47.t7 VNB.t15 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X39 VGND.t2 A1.t7 a_803_47.t2 VNB.t10 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
R0 C1.n0 C1.t3 221.719
R1 C1.n2 C1.t5 221.719
R2 C1.n8 C1.t7 221.719
R3 C1.n9 C1.t2 221.719
R4 C1.n0 C1.t1 149.419
R5 C1.n2 C1.t6 149.419
R6 C1.n8 C1.t0 149.419
R7 C1.n9 C1.t4 149.419
R8 C1.n5 C1.n3 76
R9 C1.n7 C1.n6 76
R10 C1.n11 C1.n10 76
R11 C1.n7 C1.n3 60.696
R12 C1.n10 C1.n8 58.911
R13 C1.n2 C1.n1 48.2
R14 C1.n1 C1.n0 26.777
R15 C1.n5 C1.n4 16.118
R16 C1.n10 C1.n9 16.066
R17 C1.n6 C1 15.644
R18 C1.n3 C1.n2 12.496
R19 C1 C1.n11 11.851
R20 C1.n11 C1 9.955
R21 C1.n6 C1 6.162
R22 C1.n4 C1 5.214
R23 C1.n8 C1.n7 1.785
R24 C1 C1.n5 0.474
R25 a_445_47.n4 a_445_47.n3 149.089
R26 a_445_47.n2 a_445_47.n0 149.089
R27 a_445_47.n2 a_445_47.n1 92.5
R28 a_445_47.n5 a_445_47.n4 92.5
R29 a_445_47.n4 a_445_47.n2 91.621
R30 a_445_47.n3 a_445_47.t3 24.923
R31 a_445_47.n3 a_445_47.t1 24.923
R32 a_445_47.n1 a_445_47.t7 24.923
R33 a_445_47.n1 a_445_47.t5 24.923
R34 a_445_47.n0 a_445_47.t6 24.923
R35 a_445_47.n0 a_445_47.t4 24.923
R36 a_445_47.n5 a_445_47.t2 24.923
R37 a_445_47.t0 a_445_47.n5 24.923
R38 a_27_47.n2 a_27_47.t7 227.55
R39 a_27_47.n4 a_27_47.t2 208.315
R40 a_27_47.n2 a_27_47.n1 92.5
R41 a_27_47.n3 a_27_47.n0 92.5
R42 a_27_47.n5 a_27_47.n4 92.5
R43 a_27_47.n3 a_27_47.n2 62.989
R44 a_27_47.n4 a_27_47.n3 55.341
R45 a_27_47.n0 a_27_47.t1 24.923
R46 a_27_47.n0 a_27_47.t5 24.923
R47 a_27_47.n1 a_27_47.t6 24.923
R48 a_27_47.n1 a_27_47.t4 24.923
R49 a_27_47.n5 a_27_47.t0 24.923
R50 a_27_47.t3 a_27_47.n5 24.923
R51 VNB VNB.t15 6053.91
R52 VNB.t2 VNB.t17 4545.05
R53 VNB.t7 VNB.t11 2151.65
R54 VNB.t18 VNB.t6 2151.65
R55 VNB.t4 VNB.t5 2127.47
R56 VNB.t10 VNB.t9 2030.77
R57 VNB.t8 VNB.t10 2030.77
R58 VNB.t11 VNB.t8 2030.77
R59 VNB.t5 VNB.t7 2030.77
R60 VNB.t6 VNB.t4 2030.77
R61 VNB.t16 VNB.t18 2030.77
R62 VNB.t19 VNB.t16 2030.77
R63 VNB.t17 VNB.t19 2030.77
R64 VNB.t0 VNB.t2 2030.77
R65 VNB.t3 VNB.t0 2030.77
R66 VNB.t1 VNB.t3 2030.77
R67 VNB.t13 VNB.t1 2030.77
R68 VNB.t14 VNB.t13 2030.77
R69 VNB.t12 VNB.t14 2030.77
R70 VNB.t15 VNB.t12 2030.77
R71 A2.n8 A2.t5 278.005
R72 A2.n0 A2.t6 221.719
R73 A2.n6 A2.t2 221.719
R74 A2.n0 A2.t7 209.222
R75 A2.n8 A2.t4 198.942
R76 A2.n9 A2.t3 174.936
R77 A2.n7 A2.t0 149.419
R78 A2.n2 A2.t1 149.419
R79 A2.n5 A2.n4 76
R80 A2.n11 A2.n10 76
R81 A2.n5 A2.n2 46.414
R82 A2.n9 A2.n8 33.078
R83 A2.n10 A2.n7 28.562
R84 A2.n7 A2.n6 18.744
R85 A2.n4 A2.n3 16.118
R86 A2.n2 A2.n1 14.281
R87 A2.n10 A2.n9 14.281
R88 A2.n6 A2.n5 13.388
R89 A2.n11 A2 12.8
R90 A2 A2.n11 9.007
R91 A2.n4 A2 3.318
R92 A2.n3 A2 2.37
R93 A2.n1 A2.n0 0.892
R94 VGND.n3 VGND.n0 109.784
R95 VGND.n12 VGND.n11 107.239
R96 VGND.n7 VGND.n6 106.657
R97 VGND.n2 VGND.n1 106.463
R98 VGND.n0 VGND.t1 24.923
R99 VGND.n0 VGND.t2 24.923
R100 VGND.n1 VGND.t0 24.923
R101 VGND.n1 VGND.t3 24.923
R102 VGND.n6 VGND.t7 24.923
R103 VGND.n6 VGND.t5 24.923
R104 VGND.n11 VGND.t6 24.923
R105 VGND.n11 VGND.t4 24.923
R106 VGND.n5 VGND.n4 4.65
R107 VGND.n8 VGND.n7 4.65
R108 VGND.n10 VGND.n9 4.65
R109 VGND.n13 VGND.n12 4.02
R110 VGND.n3 VGND.n2 3.891
R111 VGND VGND.n13 1.557
R112 VGND.n5 VGND.n3 0.263
R113 VGND.n13 VGND.n10 0.137
R114 VGND.n8 VGND.n5 0.119
R115 VGND.n10 VGND.n8 0.119
R116 a_803_47.n6 a_803_47.t9 218.584
R117 a_803_47.n1 a_803_47.t1 211.297
R118 a_803_47.n1 a_803_47.n0 92.5
R119 a_803_47.n3 a_803_47.n2 92.5
R120 a_803_47.n7 a_803_47.n4 92.5
R121 a_803_47.n6 a_803_47.n5 92.5
R122 a_803_47.n9 a_803_47.n8 92.5
R123 a_803_47.n8 a_803_47.n3 45.312
R124 a_803_47.n7 a_803_47.n6 44.288
R125 a_803_47.n3 a_803_47.n1 43.008
R126 a_803_47.n8 a_803_47.n7 43.008
R127 a_803_47.n4 a_803_47.t10 29.538
R128 a_803_47.n2 a_803_47.t4 29.538
R129 a_803_47.n9 a_803_47.t6 28.615
R130 a_803_47.n5 a_803_47.t8 24.923
R131 a_803_47.n5 a_803_47.t11 24.923
R132 a_803_47.n4 a_803_47.t5 24.923
R133 a_803_47.n2 a_803_47.t3 24.923
R134 a_803_47.n0 a_803_47.t2 24.923
R135 a_803_47.n0 a_803_47.t0 24.923
R136 a_803_47.t7 a_803_47.n9 24.923
R137 Y.n1 Y.t14 553.039
R138 Y.n1 Y.n0 314.489
R139 Y.n13 Y.n12 177.655
R140 Y.n3 Y.n2 176.013
R141 Y.n5 Y.n4 176.013
R142 Y.n7 Y.n6 176.013
R143 Y.n9 Y.n8 176.013
R144 Y.n11 Y.n10 176.013
R145 Y.n18 Y.t10 172.959
R146 Y.n16 Y.n14 155.747
R147 Y.n16 Y.n15 92.5
R148 Y.n6 Y.t19 66.98
R149 Y.n7 Y.n5 64.376
R150 Y.n3 Y.n1 51.576
R151 Y.n5 Y.n3 48.941
R152 Y.n9 Y.n7 48.941
R153 Y.n11 Y.n9 48.941
R154 Y.n13 Y.n11 48.941
R155 Y.n17 Y.n13 48.188
R156 Y.n2 Y.t15 31.52
R157 Y.n0 Y.t13 26.595
R158 Y.n0 Y.t12 26.595
R159 Y.n2 Y.t17 26.595
R160 Y.n4 Y.t16 26.595
R161 Y.n4 Y.t18 26.595
R162 Y.n6 Y.t2 26.595
R163 Y.n8 Y.t1 26.595
R164 Y.n8 Y.t0 26.595
R165 Y.n10 Y.t3 26.595
R166 Y.n10 Y.t4 26.595
R167 Y.n12 Y.t5 26.595
R168 Y.n12 Y.t6 26.595
R169 Y.n15 Y.t7 24.923
R170 Y.n15 Y.t11 24.923
R171 Y.n14 Y.t8 24.923
R172 Y.n14 Y.t9 24.923
R173 Y Y.n16 24.508
R174 Y.n18 Y 11.884
R175 Y Y.n17 8.405
R176 Y.n17 Y 6.841
R177 Y Y.n18 3.843
R178 a_1163_297.n4 a_1163_297.n0 292.5
R179 a_1163_297.n3 a_1163_297.n1 250.068
R180 a_1163_297.n5 a_1163_297.n4 198.421
R181 a_1163_297.n3 a_1163_297.n2 151.483
R182 a_1163_297.n4 a_1163_297.n3 85.442
R183 a_1163_297.n0 a_1163_297.t4 26.595
R184 a_1163_297.n0 a_1163_297.t7 26.595
R185 a_1163_297.n1 a_1163_297.t2 26.595
R186 a_1163_297.n1 a_1163_297.t3 26.595
R187 a_1163_297.n2 a_1163_297.t0 26.595
R188 a_1163_297.n2 a_1163_297.t1 26.595
R189 a_1163_297.t6 a_1163_297.n5 26.595
R190 a_1163_297.n5 a_1163_297.t5 26.595
R191 VPB.t12 VPB.t5 550.467
R192 VPB.t2 VPB.t19 369.937
R193 VPB.t17 VPB.t13 263.395
R194 VPB.t7 VPB.t6 248.598
R195 VPB.t4 VPB.t7 248.598
R196 VPB.t5 VPB.t4 248.598
R197 VPB.t15 VPB.t12 248.598
R198 VPB.t14 VPB.t15 248.598
R199 VPB.t13 VPB.t14 248.598
R200 VPB.t16 VPB.t17 248.598
R201 VPB.t18 VPB.t16 248.598
R202 VPB.t19 VPB.t18 248.598
R203 VPB.t1 VPB.t2 248.598
R204 VPB.t0 VPB.t1 248.598
R205 VPB.t3 VPB.t0 248.598
R206 VPB.t8 VPB.t3 248.598
R207 VPB.t9 VPB.t8 248.598
R208 VPB.t10 VPB.t9 248.598
R209 VPB.t11 VPB.t10 248.598
R210 VPB VPB.t11 189.408
R211 VPWR.n5 VPWR.t5 496.364
R212 VPWR.n2 VPWR.t6 195.972
R213 VPWR.n39 VPWR.n38 166.139
R214 VPWR.n16 VPWR.n15 165.798
R215 VPWR.n1 VPWR.n0 164.542
R216 VPWR.n29 VPWR.n28 164.542
R217 VPWR.n33 VPWR.n32 164.542
R218 VPWR.n44 VPWR.n43 164.253
R219 VPWR.n22 VPWR.n21 163.702
R220 VPWR.n0 VPWR.t7 26.595
R221 VPWR.n0 VPWR.t4 26.595
R222 VPWR.n15 VPWR.t13 26.595
R223 VPWR.n15 VPWR.t12 26.595
R224 VPWR.n21 VPWR.t14 26.595
R225 VPWR.n21 VPWR.t15 26.595
R226 VPWR.n28 VPWR.t2 26.595
R227 VPWR.n28 VPWR.t1 26.595
R228 VPWR.n32 VPWR.t0 26.595
R229 VPWR.n32 VPWR.t3 26.595
R230 VPWR.n38 VPWR.t8 26.595
R231 VPWR.n38 VPWR.t9 26.595
R232 VPWR.n43 VPWR.t10 26.595
R233 VPWR.n43 VPWR.t11 26.595
R234 VPWR.n17 VPWR.n16 5.27
R235 VPWR.n4 VPWR.n3 4.65
R236 VPWR.n6 VPWR.n5 4.65
R237 VPWR.n8 VPWR.n7 4.65
R238 VPWR.n10 VPWR.n9 4.65
R239 VPWR.n12 VPWR.n11 4.65
R240 VPWR.n14 VPWR.n13 4.65
R241 VPWR.n18 VPWR.n17 4.65
R242 VPWR.n20 VPWR.n19 4.65
R243 VPWR.n23 VPWR.n22 4.65
R244 VPWR.n25 VPWR.n24 4.65
R245 VPWR.n27 VPWR.n26 4.65
R246 VPWR.n31 VPWR.n30 4.65
R247 VPWR.n35 VPWR.n34 4.65
R248 VPWR.n37 VPWR.n36 4.65
R249 VPWR.n40 VPWR.n39 4.65
R250 VPWR.n42 VPWR.n41 4.65
R251 VPWR.n30 VPWR.n29 4.141
R252 VPWR.n45 VPWR.n44 3.958
R253 VPWR.n2 VPWR.n1 3.727
R254 VPWR.n34 VPWR.n33 1.129
R255 VPWR.n4 VPWR.n2 0.258
R256 VPWR.n45 VPWR.n42 0.137
R257 VPWR VPWR.n45 0.122
R258 VPWR.n6 VPWR.n4 0.119
R259 VPWR.n8 VPWR.n6 0.119
R260 VPWR.n10 VPWR.n8 0.119
R261 VPWR.n12 VPWR.n10 0.119
R262 VPWR.n14 VPWR.n12 0.119
R263 VPWR.n18 VPWR.n14 0.119
R264 VPWR.n20 VPWR.n18 0.119
R265 VPWR.n23 VPWR.n20 0.119
R266 VPWR.n25 VPWR.n23 0.119
R267 VPWR.n27 VPWR.n25 0.119
R268 VPWR.n31 VPWR.n27 0.119
R269 VPWR.n35 VPWR.n31 0.119
R270 VPWR.n37 VPWR.n35 0.119
R271 VPWR.n40 VPWR.n37 0.119
R272 VPWR.n42 VPWR.n40 0.119
R273 D1.n1 D1.t0 192.799
R274 D1.n0 D1.t1 192.799
R275 D1.n5 D1.t2 192.799
R276 D1.n6 D1.t6 192.799
R277 D1.n1 D1.t4 149.419
R278 D1.n0 D1.t5 149.419
R279 D1.n5 D1.t3 149.419
R280 D1.n6 D1.t7 149.419
R281 D1 D1.n2 77.659
R282 D1.n4 D1.n3 76
R283 D1.n8 D1.n7 76
R284 D1.n2 D1.n0 34.141
R285 D1.n7 D1.n6 32.133
R286 D1.n5 D1.n4 30.794
R287 D1.n4 D1.n0 25.438
R288 D1.n7 D1.n5 24.1
R289 D1.n2 D1.n1 22.091
R290 D1.n3 D1 19.437
R291 D1.n8 D1 17.066
R292 D1 D1.n8 4.74
R293 D1.n3 D1 2.37
R294 B1.n10 B1.t7 260.279
R295 B1.n1 B1.t4 233.839
R296 B1.n1 B1.t3 222.716
R297 B1.n3 B1.t2 221.719
R298 B1.n8 B1.t5 221.719
R299 B1.n2 B1.t0 168.699
R300 B1.n9 B1.t1 147.813
R301 B1.n0 B1.t6 147.813
R302 B1.n5 B1.n4 76
R303 B1.n7 B1.n6 76
R304 B1.n11 B1.n10 76
R305 B1.n4 B1.n2 53.458
R306 B1.n7 B1.n0 30.672
R307 B1.n8 B1.n7 24.538
R308 B1 B1.n11 20.385
R309 B1.n3 B1.n0 18.403
R310 B1.n9 B1.n8 18.403
R311 B1.n10 B1.n9 16.65
R312 B1.n6 B1 14.696
R313 B1.n5 B1 12.8
R314 B1.n4 B1.n3 10.516
R315 B1 B1.n5 9.007
R316 B1.n2 B1.n1 7.914
R317 B1.n6 B1 7.111
R318 B1.n11 B1 1.422
R319 A1.n1 A1.t0 248.496
R320 A1.n0 A1.t2 221.719
R321 A1.n7 A1.t3 221.719
R322 A1.n11 A1.t5 221.719
R323 A1.n11 A1.t1 176.196
R324 A1.n10 A1.t4 149.419
R325 A1.n6 A1.t7 149.419
R326 A1.n1 A1.t6 149.419
R327 A1.n3 A1.n2 76
R328 A1.n5 A1.n4 76
R329 A1.n9 A1.n8 76
R330 A1.n13 A1.n12 76
R331 A1.n7 A1.n6 48.2
R332 A1.n2 A1.n0 42.844
R333 A1.n12 A1.n10 37.488
R334 A1.n5 A1.n0 17.851
R335 A1.n13 A1.n9 16.422
R336 A1.n3 A1 16.181
R337 A1.n4 A1 11.833
R338 A1.n12 A1.n11 10.711
R339 A1.n4 A1 10.384
R340 A1.n6 A1.n5 8.925
R341 A1 A1.n3 6.037
R342 A1.n2 A1.n1 5.355
R343 A1.n9 A1 4.588
R344 A1.n8 A1.n7 3.57
R345 A1 A1.n13 1.207
C0 C1 Y 0.42fF
C1 VPWR VGND 0.21fF
C2 B1 Y 0.43fF
C3 Y VPWR 1.70fF
C4 A2 Y 0.32fF
C5 VPB VPWR 0.19fF
C6 D1 Y 0.50fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__or2_0.ext - technology: sky130A

.subckt sky130_fd_sc_hd__or2_0 A X B VGND VPWR VNB VPB
X0 VGND.t0 A.t0 a_68_355.t0 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1 a_150_355.t1 B.t0 a_68_355.t1 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 a_68_355.t2 B.t1 VGND.t1 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3 X.t1 a_68_355.t3 VGND.t2 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 VPWR.t0 A.t1 a_150_355.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 X.t0 a_68_355.t4 VPWR.t1 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
R0 A.n0 A.t1 241.535
R1 A.n0 A.t0 132.281
R2 A.n1 A.n0 76
R3  A.n1 11.224
R4 A.n1 A 2.166
R5 a_68_355.n1 a_68_355.t1 370.207
R6 a_68_355.n0 a_68_355.t4 271.526
R7 a_68_355.n1 a_68_355.n0 187.434
R8 a_68_355.n2 a_68_355.n1 172.324
R9 a_68_355.n0 a_68_355.t3 126.926
R10 a_68_355.t0 a_68_355.n2 38.571
R11 a_68_355.n2 a_68_355.t2 38.571
R12 VGND.n1 VGND.t1 170.818
R13 VGND.n1 VGND.n0 136.769
R14 VGND.n0 VGND.t0 55.714
R15 VGND.n0 VGND.t2 40
R16 VGND VGND.n1 0.145
R17 VNB VNB.t1 13557.8
R18 VNB.t0 VNB.t2 3138.24
R19 VNB.t1 VNB.t0 2717.65
R20 B.n0 B.t0 227.986
R21 B.n0 B.t1 118.732
R22 B B.n0 81.574
R23 a_150_355.t0 a_150_355.t1 98.5
R24 VPB VPB.t2 313.707
R25 VPB.t0 VPB.t1 287.071
R26 VPB.t2 VPB.t0 213.084
R27 X X.t0 381.046
R28 X X.t1 181.935
R29 VPWR VPWR.n0 320.22
R30 VPWR.n0 VPWR.t0 96.154
R31 VPWR.n0 VPWR.t1 40.016
C0 VPWR X 0.15fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__or2_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__or2_1 A X B VGND VPWR VNB VPB
X0 VGND.t1 A.t0 a_68_297.t2 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1 a_68_297.t1 B.t0 VGND.t0 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 X.t1 a_68_297.t3 VGND.t2 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 VPWR.t0 A.t1 a_150_297.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 X.t0 a_68_297.t4 VPWR.t1 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 a_150_297.t1 B.t1 a_68_297.t0 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
R0 A.n0 A.t0 206.188
R1 A.n0 A.t1 148.348
R2 A A.n0 78.656
R3  A 16.422
R4 a_68_297.t0 a_68_297.n2 370.207
R5 a_68_297.n1 a_68_297.t4 236.179
R6 a_68_297.n2 a_68_297.n0 167.806
R7 a_68_297.n2 a_68_297.n1 165.599
R8 a_68_297.n1 a_68_297.t3 163.879
R9 a_68_297.n0 a_68_297.t2 38.571
R10 a_68_297.n0 a_68_297.t1 38.571
R11 VGND.n1 VGND.t0 158.551
R12 VGND.n1 VGND.n0 123.076
R13 VGND.n0 VGND.t1 55.714
R14 VGND.n0 VGND.t2 26.857
R15 VGND VGND.n1 0.145
R16 VNB VNB.t0 7424.51
R17 VNB.t0 VNB.t1 2717.65
R18 VNB.t1 VNB.t2 2303.7
R19 B.n0 B.t0 192.639
R20 B.n0 B.t1 134.799
R21 B B.n0 77.983
R22  B 12.259
R23 X.n0 X.t0 194.32
R24 X X.t1 128.201
R25 X.n0 X 2.438
R26 X X.n0 1.435
R27 a_150_297.t0 a_150_297.t1 98.5
R28 VPWR VPWR.n0 172.477
R29 VPWR.n0 VPWR.t0 96.154
R30 VPWR.n0 VPWR.t1 25.61
R31 VPB VPB.t2 313.707
R32 VPB.t0 VPB.t1 287.071
R33 VPB.t2 VPB.t0 213.084
C0 VPWR X 0.18fF
C1 X VGND 0.15fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__or2_2.ext - technology: sky130A

.subckt sky130_fd_sc_hd__or2_2 B X A VPWR VGND VNB VPB
X0 a_121_297.t1 B.t0 a_39_297.t2 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1 X.t1 a_39_297.t3 VGND.t2 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 VPWR.t2 a_39_297.t4 X.t3 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 X.t2 a_39_297.t5 VPWR.t1 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 VGND.t1 a_39_297.t6 X.t0 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 VPWR.t0 A.t0 a_121_297.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 VGND.t0 A.t1 a_39_297.t0 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7 a_39_297.t1 B.t1 VGND.t3 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
R0 B.n0 B.t1 193.301
R1 B.n0 B.t0 135.461
R2 B B.n0 79.61
R3  B 22.317
R4 a_39_297.n3 a_39_297.t2 363.055
R5 a_39_297.n0 a_39_297.t4 212.079
R6 a_39_297.n1 a_39_297.t5 212.079
R7 a_39_297.n4 a_39_297.n3 169.826
R8 a_39_297.n3 a_39_297.n2 164.093
R9 a_39_297.n0 a_39_297.t6 139.779
R10 a_39_297.n1 a_39_297.t3 139.779
R11 a_39_297.n2 a_39_297.n0 41.627
R12 a_39_297.t0 a_39_297.n4 38.571
R13 a_39_297.n4 a_39_297.t1 38.571
R14 a_39_297.n2 a_39_297.n1 19.718
R15 a_121_297.t0 a_121_297.t1 98.5
R16 VPB.t0 VPB.t1 298.909
R17 VPB.t1 VPB.t2 248.598
R18 VPB VPB.t3 224.922
R19 VPB.t3 VPB.t0 213.084
R20 VGND.n2 VGND.t1 189.995
R21 VGND.n5 VGND.t3 154.004
R22 VGND.n1 VGND.n0 109.973
R23 VGND.n0 VGND.t0 61.428
R24 VGND.n0 VGND.t2 25.846
R25 VGND.n6 VGND.n5 4.65
R26 VGND.n4 VGND.n3 4.65
R27 VGND.n2 VGND.n1 3.736
R28 VGND.n4 VGND.n2 0.269
R29 VGND.n6 VGND.n4 0.119
R30 VGND VGND.n6 0.02
R31 X X.n0 157.725
R32 X X.n1 143.934
R33 X.n0 X.t3 26.595
R34 X.n0 X.t2 26.595
R35 X.n1 X.t0 24.923
R36 X.n1 X.t1 24.923
R37 VNB VNB.t3 6438.23
R38 VNB.t3 VNB.t0 2717.65
R39 VNB.t0 VNB.t2 2400.4
R40 VNB.t2 VNB.t1 2030.77
R41 VPWR.n1 VPWR.t2 590.294
R42 VPWR.n1 VPWR.n0 180.082
R43 VPWR.n0 VPWR.t0 101.83
R44 VPWR.n0 VPWR.t1 26.595
R45 VPWR VPWR.n1 0.402
R46 A.n0 A.t1 206.188
R47 A.n0 A.t0 148.348
R48 A A.n0 77.717
R49  A 10.614
C0 VPWR X 0.23fF
C1 X VGND 0.16fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__or2_4.ext - technology: sky130A

.subckt sky130_fd_sc_hd__or2_4 X A B VGND VPWR VNB VPB
X0 a_121_297.t1 B.t0 a_35_297.t2 VPB.t5 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 VPWR.t3 a_35_297.t3 X.t7 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 X.t6 a_35_297.t4 VPWR.t2 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 X.t3 a_35_297.t5 VGND.t3 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 X.t2 a_35_297.t6 VGND.t2 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 VPWR.t1 a_35_297.t7 X.t5 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 X.t4 a_35_297.t8 VPWR.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 VGND.t1 a_35_297.t9 X.t1 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 VPWR.t4 A.t0 a_121_297.t0 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 VGND.t0 a_35_297.t10 X.t0 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 VGND.t4 A.t1 a_35_297.t0 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 a_35_297.t1 B.t1 VGND.t5 VNB.t5 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
R0 B.n0 B.t0 228.647
R1 B.n0 B.t1 156.347
R2 B B.n0 78.76
R3  B 17.066
R4 a_35_297.n0 a_35_297.t3 212.079
R5 a_35_297.n1 a_35_297.t4 212.079
R6 a_35_297.n5 a_35_297.t7 212.079
R7 a_35_297.n6 a_35_297.t8 212.079
R8 a_35_297.n0 a_35_297.t10 139.779
R9 a_35_297.n1 a_35_297.t6 139.779
R10 a_35_297.n5 a_35_297.t9 139.779
R11 a_35_297.n6 a_35_297.t5 139.779
R12 a_35_297.t2 a_35_297.n10 131.986
R13 a_35_297.n10 a_35_297.n9 106.312
R14 a_35_297.n4 a_35_297.n2 101.6
R15 a_35_297.n10 a_35_297.n8 80.059
R16 a_35_297.n4 a_35_297.n3 76
R17 a_35_297.n8 a_35_297.n7 76
R18 a_35_297.n2 a_35_297.n0 58.424
R19 a_35_297.n7 a_35_297.n5 35.054
R20 a_35_297.n7 a_35_297.n6 26.29
R21 a_35_297.n9 a_35_297.t0 24.923
R22 a_35_297.n9 a_35_297.t1 24.923
R23 a_35_297.n8 a_35_297.n4 22.588
R24 a_35_297.n2 a_35_297.n1 2.921
R25 a_121_297.t0 a_121_297.t1 41.37
R26 VPB.t4 VPB.t0 298.909
R27 VPB.t2 VPB.t3 248.598
R28 VPB.t1 VPB.t2 248.598
R29 VPB.t0 VPB.t1 248.598
R30 VPB VPB.t5 224.922
R31 VPB.t5 VPB.t4 213.084
R32 X.n2 X.n0 194.359
R33 X.n2 X.n1 98.052
R34 X.n5 X.n3 90.831
R35 X.n5 X.n4 52.431
R36 X X.n5 36.74
R37 X X.n2 28.144
R38 X.n1 X.t7 26.595
R39 X.n1 X.t6 26.595
R40 X.n0 X.t5 26.595
R41 X.n0 X.t4 26.595
R42 X.n3 X.t1 24.923
R43 X.n3 X.t3 24.923
R44 X.n4 X.t0 24.923
R45 X.n4 X.t2 24.923
R46 VPWR.n1 VPWR.n0 314.711
R47 VPWR.n2 VPWR.t3 210.693
R48 VPWR.n6 VPWR.n5 173.841
R49 VPWR.n5 VPWR.t4 35.46
R50 VPWR.n5 VPWR.t0 34.475
R51 VPWR.n0 VPWR.t2 26.595
R52 VPWR.n0 VPWR.t1 26.595
R53 VPWR.n2 VPWR.n1 7.37
R54 VPWR.n8 VPWR.n7 4.65
R55 VPWR.n4 VPWR.n3 4.65
R56 VPWR.n7 VPWR.n6 0.376
R57 VPWR.n4 VPWR.n2 0.292
R58 VPWR.n9 VPWR.n8 0.132
R59 VPWR VPWR.n9 0.127
R60 VPWR.n8 VPWR.n4 0.119
R61 VGND.n2 VGND.t0 199.568
R62 VGND.n11 VGND.t5 183.596
R63 VGND.n6 VGND.n5 129.394
R64 VGND.n1 VGND.n0 116.217
R65 VGND.n5 VGND.t4 33.23
R66 VGND.n5 VGND.t3 32.307
R67 VGND.n0 VGND.t2 24.923
R68 VGND.n0 VGND.t1 24.923
R69 VGND.n2 VGND.n1 7.37
R70 VGND.n12 VGND.n11 4.65
R71 VGND.n4 VGND.n3 4.65
R72 VGND.n8 VGND.n7 4.65
R73 VGND.n10 VGND.n9 4.65
R74 VGND.n7 VGND.n6 0.376
R75 VGND.n4 VGND.n2 0.292
R76 VGND.n8 VGND.n4 0.119
R77 VGND.n10 VGND.n8 0.119
R78 VGND.n12 VGND.n10 0.119
R79 VGND VGND.n12 0.02
R80 VNB VNB.t5 6053.91
R81 VNB.t4 VNB.t3 2441.76
R82 VNB.t2 VNB.t0 2030.77
R83 VNB.t1 VNB.t2 2030.77
R84 VNB.t3 VNB.t1 2030.77
R85 VNB.t5 VNB.t4 2030.77
R86 A.n0 A.t0 241.534
R87 A.n0 A.t1 169.234
R88 A A.n0 80.654
C0 X VGND 0.44fF
C1 VPWR X 0.49fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__or2b_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__or2b_1 A B_N X VGND VPWR VNB VPB
X0 a_219_297.t1 a_27_53.t2 VGND.t0 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1 VGND.t1 B_N.t0 a_27_53.t0 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 VPWR.t1 A.t0 a_301_297.t1 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3 X.t1 a_219_297.t3 VGND.t3 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 a_301_297.t0 a_27_53.t3 a_219_297.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 X.t0 a_219_297.t4 VPWR.t0 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 a_27_53.t1 B_N.t1 VPWR.t2 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7 VGND.t2 A.t1 a_219_297.t2 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
R0 a_27_53.n1 a_27_53.t1 379.583
R1 a_27_53.n0 a_27_53.t2 186.028
R2 a_27_53.t0 a_27_53.n1 168.69
R3 a_27_53.n0 a_27_53.t3 137.828
R4 a_27_53.n1 a_27_53.n0 95.393
R5 VGND.n1 VGND.n0 108.687
R6 VGND.n3 VGND.n2 92.5
R7 VGND.n7 VGND.n6 92.5
R8 VGND.n0 VGND.t2 52.857
R9 VGND.n2 VGND.t0 38.571
R10 VGND.n6 VGND.t1 38.571
R11 VGND.n0 VGND.t3 27.568
R12 VGND.n9 VGND.n8 4.65
R13 VGND.n5 VGND.n4 4.65
R14 VGND.n5 VGND.n1 0.864
R15 VGND.n4 VGND.n3 0.196
R16 VGND.n8 VGND.n7 0.196
R17 VGND.n9 VGND.n5 0.119
R18 VGND.n10 VGND.n9 0.119
R19 VGND VGND.n10 0.02
R20 a_219_297.t0 a_219_297.n2 439.31
R21 a_219_297.n0 a_219_297.t4 240.482
R22 a_219_297.n2 a_219_297.n1 171.328
R23 a_219_297.n0 a_219_297.t3 168.182
R24 a_219_297.n2 a_219_297.n0 76
R25 a_219_297.n1 a_219_297.t2 38.571
R26 a_219_297.n1 a_219_297.t1 38.571
R27 VNB VNB.t1 7214.71
R28 VNB.t1 VNB.t0 5823.53
R29 VNB.t0 VNB.t3 2717.65
R30 VNB.t3 VNB.t2 2327.87
R31 B_N.n0 B_N.t0 185.375
R32 B_N.n0 B_N.t1 137.175
R33 B_N B_N.n0 81.632
R34 A A.t0 487.895
R35 A.t0 A.t1 392.026
R36 a_301_297.t0 a_301_297.t1 98.5
R37 VPWR.n1 VPWR.t2 413.04
R38 VPWR.n1 VPWR.n0 173.038
R39 VPWR.n0 VPWR.t1 96.154
R40 VPWR.n0 VPWR.t0 26.595
R41 VPWR VPWR.n1 0.039
R42 VPB.t3 VPB.t0 568.224
R43 VPB.t2 VPB.t1 290.031
R44 VPB.t0 VPB.t2 213.084
R45 VPB VPB.t3 189.408
R46 X X.t0 214.087
R47 X X.t1 194.571
C0 VPWR X 0.13fF
C1 VPWR A 0.25fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__or2b_2.ext - technology: sky130A

.subckt sky130_fd_sc_hd__or2b_2 A B_N X VPWR VGND VNB VPB
X0 VPWR.t3 A.t0 a_300_297.t1 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1 a_218_297.t1 a_27_53.t2 VGND.t4 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 VGND.t0 B_N.t0 a_27_53.t0 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3 a_300_297.t0 a_27_53.t3 a_218_297.t2 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 X.t1 a_218_297.t3 VGND.t1 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 VPWR.t1 a_218_297.t4 X.t3 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 X.t2 a_218_297.t5 VPWR.t2 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 VGND.t2 a_218_297.t6 X.t0 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 a_27_53.t1 B_N.t1 VPWR.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9 VGND.t3 A.t1 a_218_297.t0 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
R0 A A.t0 487.902
R1 A.t0 A.t1 392.026
R2 a_300_297.t0 a_300_297.t1 98.5
R3 VPWR.n9 VPWR.t0 408.005
R4 VPWR.n1 VPWR.n0 169.105
R5 VPWR.n2 VPWR.t1 156.652
R6 VPWR.n0 VPWR.t3 96.154
R7 VPWR.n0 VPWR.t2 26.595
R8 VPWR.n6 VPWR.n5 4.65
R9 VPWR.n8 VPWR.n7 4.65
R10 VPWR.n10 VPWR.n9 4.65
R11 VPWR.n4 VPWR.n3 4.65
R12 VPWR.n2 VPWR.n1 3.903
R13 VPWR.n4 VPWR.n2 0.237
R14 VPWR.n6 VPWR.n4 0.119
R15 VPWR.n8 VPWR.n6 0.119
R16 VPWR.n10 VPWR.n8 0.119
R17 VPWR VPWR.n10 0.02
R18 VPB.t0 VPB.t1 565.264
R19 VPB.t4 VPB.t3 290.031
R20 VPB.t3 VPB.t2 248.598
R21 VPB.t1 VPB.t4 213.084
R22 VPB VPB.t0 189.408
R23 a_27_53.n1 a_27_53.t1 380.142
R24 a_27_53.n0 a_27_53.t2 186.028
R25 a_27_53.t0 a_27_53.n1 168.627
R26 a_27_53.n0 a_27_53.t3 137.828
R27 a_27_53.n1 a_27_53.n0 95.393
R28 VGND.n2 VGND.t2 106.595
R29 VGND.n1 VGND.n0 105.973
R30 VGND.n6 VGND.n5 92.5
R31 VGND.n10 VGND.n9 92.5
R32 VGND.n0 VGND.t3 52.857
R33 VGND.n5 VGND.t4 38.571
R34 VGND.n9 VGND.t0 38.571
R35 VGND.n0 VGND.t1 27.568
R36 VGND.n12 VGND.n11 4.65
R37 VGND.n8 VGND.n7 4.65
R38 VGND.n4 VGND.n3 4.65
R39 VGND.n2 VGND.n1 3.868
R40 VGND.n4 VGND.n2 0.242
R41 VGND.n11 VGND.n10 0.196
R42 VGND.n8 VGND.n4 0.119
R43 VGND.n12 VGND.n8 0.119
R44 VGND.n13 VGND.n12 0.119
R45 VGND.n7 VGND.n6 0.098
R46 VGND VGND.n13 0.022
R47 a_218_297.n2 a_218_297.t2 439.31
R48 a_218_297.n0 a_218_297.t4 212.079
R49 a_218_297.n1 a_218_297.t5 212.079
R50 a_218_297.n3 a_218_297.n2 171.328
R51 a_218_297.n0 a_218_297.t6 139.779
R52 a_218_297.n1 a_218_297.t3 139.779
R53 a_218_297.n2 a_218_297.n1 86.224
R54 a_218_297.n1 a_218_297.n0 61.345
R55 a_218_297.t0 a_218_297.n3 38.571
R56 a_218_297.n3 a_218_297.t1 38.571
R57 VNB VNB.t0 7247.06
R58 VNB.t0 VNB.t4 5791.18
R59 VNB.t4 VNB.t3 2717.65
R60 VNB.t3 VNB.t2 2327.87
R61 VNB.t2 VNB.t1 2030.77
R62 B_N.n0 B_N.t0 185.168
R63 B_N.n0 B_N.t1 136.968
R64 B_N B_N.n0 81.632
R65 X X.n1 173.44
R66 X X.n0 154.172
R67 X.n0 X.t3 26.595
R68 X.n0 X.t2 26.595
R69 X.n1 X.t0 24.923
R70 X.n1 X.t1 24.923
C0 VPWR A 0.25fF
C1 VPWR X 0.23fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__or2b_4.ext - technology: sky130A

.subckt sky130_fd_sc_hd__or2b_4 A B_N X VGND VPWR VNB VPB
X0 VPWR.t5 a_219_297.t3 X.t7 VPB.t6 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 VGND.t6 B_N.t0 a_27_53.t0 VNB.t6 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 VPWR.t1 A.t0 a_301_297.t1 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 a_27_53.t1 B_N.t1 VPWR.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 X.t3 a_219_297.t4 VGND.t4 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 a_301_297.t0 a_27_53.t2 a_219_297.t2 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 X.t6 a_219_297.t5 VPWR.t4 VPB.t5 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 VGND.t0 A.t1 a_219_297.t0 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 VPWR.t3 a_219_297.t6 X.t5 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 VGND.t3 a_219_297.t7 X.t2 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 X.t4 a_219_297.t8 VPWR.t2 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 VGND.t2 a_219_297.t9 X.t1 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 a_219_297.t1 a_27_53.t3 VGND.t5 VNB.t5 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 X.t0 a_219_297.t10 VGND.t1 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
R0 a_219_297.n0 a_219_297.t3 212.079
R1 a_219_297.n2 a_219_297.t5 212.079
R2 a_219_297.n5 a_219_297.t6 212.079
R3 a_219_297.n6 a_219_297.t8 212.079
R4 a_219_297.t2 a_219_297.n10 161.295
R5 a_219_297.n0 a_219_297.t9 139.779
R6 a_219_297.n2 a_219_297.t10 139.779
R7 a_219_297.n5 a_219_297.t7 139.779
R8 a_219_297.n6 a_219_297.t4 139.779
R9 a_219_297.n10 a_219_297.n9 106.002
R10 a_219_297.n10 a_219_297.n8 105.033
R11 a_219_297.n4 a_219_297.n1 101.6
R12 a_219_297.n4 a_219_297.n3 76
R13 a_219_297.n8 a_219_297.n7 76
R14 a_219_297.n7 a_219_297.n6 54.772
R15 a_219_297.n1 a_219_297.n0 29.942
R16 a_219_297.n8 a_219_297.n4 25.6
R17 a_219_297.n9 a_219_297.t0 24.923
R18 a_219_297.n9 a_219_297.t1 24.923
R19 a_219_297.n3 a_219_297.n2 18.257
R20 a_219_297.n7 a_219_297.n5 6.572
R21 X.n2 X.n1 183.822
R22 X.n2 X.n0 99.472
R23 X.n5 X.n3 90.831
R24 X.n5 X.n4 52.431
R25 X X.n5 33.955
R26 X.n0 X.t7 26.595
R27 X.n0 X.t6 26.595
R28 X.n1 X.t5 26.595
R29 X.n1 X.t4 26.595
R30 X.n3 X.t2 24.923
R31 X.n3 X.t3 24.923
R32 X.n4 X.t1 24.923
R33 X.n4 X.t0 24.923
R34 X X.n2 22.15
R35 VPWR.n14 VPWR.t0 377.405
R36 VPWR.n1 VPWR.n0 314.004
R37 VPWR.n2 VPWR.t5 203.7
R38 VPWR.n6 VPWR.n5 167.407
R39 VPWR.n5 VPWR.t1 39.4
R40 VPWR.n5 VPWR.t2 27.58
R41 VPWR.n0 VPWR.t4 26.595
R42 VPWR.n0 VPWR.t3 26.595
R43 VPWR.n4 VPWR.n3 4.65
R44 VPWR.n7 VPWR.n6 4.65
R45 VPWR.n9 VPWR.n8 4.65
R46 VPWR.n11 VPWR.n10 4.65
R47 VPWR.n13 VPWR.n12 4.65
R48 VPWR.n15 VPWR.n14 4.65
R49 VPWR.n2 VPWR.n1 3.934
R50 VPWR.n4 VPWR.n2 0.293
R51 VPWR.n7 VPWR.n4 0.119
R52 VPWR.n9 VPWR.n7 0.119
R53 VPWR.n11 VPWR.n9 0.119
R54 VPWR.n13 VPWR.n11 0.119
R55 VPWR.n15 VPWR.n13 0.119
R56 VPWR VPWR.n15 0.022
R57 VPB.t0 VPB.t2 568.224
R58 VPB.t1 VPB.t3 290.031
R59 VPB.t5 VPB.t6 248.598
R60 VPB.t4 VPB.t5 248.598
R61 VPB.t3 VPB.t4 248.598
R62 VPB.t2 VPB.t1 213.084
R63 VPB VPB.t0 192.367
R64 B_N.n0 B_N.t1 323.548
R65 B_N.n0 B_N.t0 185.375
R66 B_N.n1 B_N.n0 76
R67  B_N.n1 10.889
R68 B_N.n1 B_N 2.101
R69 a_27_53.n1 a_27_53.t1 425.725
R70 a_27_53.n0 a_27_53.t2 220.842
R71 a_27_53.t0 a_27_53.n1 172.712
R72 a_27_53.n0 a_27_53.t3 139.779
R73 a_27_53.n1 a_27_53.n0 129.312
R74 VGND.n2 VGND.t2 188.958
R75 VGND.n1 VGND.n0 115.088
R76 VGND.n11 VGND.n10 98.668
R77 VGND.n15 VGND.n14 92.5
R78 VGND.n6 VGND.n5 80.988
R79 VGND.n14 VGND.t6 38.571
R80 VGND.n5 VGND.t0 37.846
R81 VGND.n0 VGND.t1 24.923
R82 VGND.n0 VGND.t3 24.923
R83 VGND.n5 VGND.t4 24.923
R84 VGND.n10 VGND.t5 18.526
R85 VGND.n2 VGND.n1 9.975
R86 VGND.n17 VGND.n16 4.65
R87 VGND.n13 VGND.n12 4.65
R88 VGND.n4 VGND.n3 4.65
R89 VGND.n7 VGND.n6 4.65
R90 VGND.n9 VGND.n8 4.65
R91 VGND.n4 VGND.n2 0.322
R92 VGND.n12 VGND.n11 0.196
R93 VGND.n16 VGND.n15 0.196
R94 VGND.n7 VGND.n4 0.119
R95 VGND.n9 VGND.n7 0.119
R96 VGND.n13 VGND.n9 0.119
R97 VGND.n17 VGND.n13 0.119
R98 VGND.n18 VGND.n17 0.119
R99 VGND VGND.n18 0.022
R100 VNB VNB.t6 6404.97
R101 VNB.t6 VNB.t5 4773.87
R102 VNB.t0 VNB.t4 2369.23
R103 VNB.t1 VNB.t2 2030.77
R104 VNB.t3 VNB.t1 2030.77
R105 VNB.t4 VNB.t3 2030.77
R106 VNB.t5 VNB.t0 2030.77
R107 A.n0 A.t0 241.534
R108 A.n0 A.t1 169.234
R109 A A.n0 84.64
R110 a_301_297.t0 a_301_297.t1 41.37
C0 VPWR X 0.53fF
C1 X VGND 0.41fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__or3_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__or3_1 A X B C VPWR VGND VNB VPB
X0 X.t1 a_29_53.t4 VPWR.t1 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_111_297.t1 C.t0 a_29_53.t2 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 X.t0 a_29_53.t5 VGND.t3 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 a_183_297.t0 B.t0 a_111_297.t0 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 VPWR.t0 A.t0 a_183_297.t1 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 a_29_53.t0 B.t1 VGND.t0 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 VGND.t2 C.t1 a_29_53.t3 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7 VGND.t1 A.t1 a_29_53.t1 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
R0 a_29_53.n1 a_29_53.t2 486.739
R1 a_29_53.n0 a_29_53.t4 241.534
R2 a_29_53.n2 a_29_53.t3 201.47
R3 a_29_53.n0 a_29_53.t5 169.234
R4 a_29_53.n3 a_29_53.n2 106.429
R5 a_29_53.n1 a_29_53.n0 76
R6 a_29_53.n2 a_29_53.n1 63.397
R7 a_29_53.n3 a_29_53.t1 38.571
R8 a_29_53.t0 a_29_53.n3 38.571
R9 VPWR VPWR.n0 172.957
R10 VPWR.n0 VPWR.t0 96.154
R11 VPWR.n0 VPWR.t1 26.595
R12 X X.t1 211.8
R13 X X.t0 194.174
R14 VPB.t0 VPB.t3 290.031
R15 VPB.t1 VPB.t0 284.112
R16 VPB.t2 VPB.t1 213.084
R17 VPB VPB.t2 201.246
R18 C.n0 C.t1 185.375
R19 C.n0 C.t0 137.175
R20 C C.n0 80.46
R21 a_111_297.t0 a_111_297.t1 98.5
R22 VGND.n2 VGND.n1 111.327
R23 VGND.n2 VGND.n0 109.414
R24 VGND.n0 VGND.t1 52.857
R25 VGND.n1 VGND.t0 38.571
R26 VGND.n1 VGND.t2 38.571
R27 VGND.n0 VGND.t3 27.568
R28 VGND VGND.n2 0.244
R29 VNB VNB.t2 7344.12
R30 VNB.t0 VNB.t1 2717.65
R31 VNB.t2 VNB.t0 2717.65
R32 VNB.t1 VNB.t3 2327.87
R33 B.t0 B.t1 378.254
R34 B B.t0 253.559
R35 a_183_297.t0 a_183_297.t1 154.785
R36 A.n0 A.t1 196.548
R37 A.n0 A.t0 148.348
R38 A A.n0 85.503
R39 A A.n1 14.157
R40 A.n1 A 7.876
R41 A.n1 A 3.684
C0 VPWR X 0.13fF
C1 VPWR B 0.20fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__or3_2.ext - technology: sky130A

.subckt sky130_fd_sc_hd__or3_2 A B X C VGND VPWR VNB VPB
X0 VPWR.t1 a_30_53.t4 X.t3 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 VGND.t1 a_30_53.t5 X.t1 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 X.t2 a_30_53.t6 VPWR.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 a_112_297.t0 C.t0 a_30_53.t1 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 X.t0 a_30_53.t7 VGND.t0 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 VGND.t3 A.t0 a_30_53.t2 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 a_30_53.t0 B.t0 VGND.t2 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7 VGND.t4 C.t1 a_30_53.t3 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 a_184_297.t0 B.t1 a_112_297.t1 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9 VPWR.t2 A.t1 a_184_297.t1 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
R0 a_30_53.n2 a_30_53.t1 486.628
R1 a_30_53.n0 a_30_53.t4 212.079
R2 a_30_53.n1 a_30_53.t6 212.079
R3 a_30_53.n3 a_30_53.t3 201.47
R4 a_30_53.n0 a_30_53.t5 139.779
R5 a_30_53.n1 a_30_53.t7 139.779
R6 a_30_53.n4 a_30_53.n3 106.429
R7 a_30_53.n2 a_30_53.n1 79.651
R8 a_30_53.n3 a_30_53.n2 63.397
R9 a_30_53.n1 a_30_53.n0 61.345
R10 a_30_53.n4 a_30_53.t2 38.571
R11 a_30_53.t0 a_30_53.n4 38.571
R12 X X.n1 169.251
R13 X X.n0 152.895
R14 X.n0 X.t3 26.595
R15 X.n0 X.t2 26.595
R16 X.n1 X.t1 24.923
R17 X.n1 X.t0 24.923
R18 VPWR.n1 VPWR.n0 172.493
R19 VPWR.n1 VPWR.t1 159.625
R20 VPWR.n0 VPWR.t2 96.154
R21 VPWR.n0 VPWR.t0 26.595
R22 VPWR VPWR.n1 0.456
R23 VPB.t4 VPB.t0 290.031
R24 VPB.t2 VPB.t4 284.112
R25 VPB.t0 VPB.t1 248.598
R26 VPB.t3 VPB.t2 213.084
R27 VPB VPB.t3 201.246
R28 VGND.n6 VGND.n5 108.015
R29 VGND.n1 VGND.n0 105.973
R30 VGND.n2 VGND.t1 100.988
R31 VGND.n0 VGND.t3 52.857
R32 VGND.n5 VGND.t2 38.571
R33 VGND.n5 VGND.t4 38.571
R34 VGND.n0 VGND.t0 27.568
R35 VGND.n4 VGND.n3 4.65
R36 VGND.n7 VGND.n6 3.958
R37 VGND.n2 VGND.n1 3.881
R38 VGND.n4 VGND.n2 0.231
R39 VGND.n7 VGND.n4 0.137
R40 VGND VGND.n7 0.124
R41 VNB VNB.t4 7344.12
R42 VNB.t2 VNB.t3 2717.65
R43 VNB.t4 VNB.t2 2717.65
R44 VNB.t3 VNB.t0 2327.87
R45 VNB.t0 VNB.t1 2030.77
R46 C.n0 C.t1 185.168
R47 C.n0 C.t0 136.968
R48 C C.n0 80.266
R49 a_112_297.t0 a_112_297.t1 98.5
R50 A.n0 A.t0 196.548
R51 A.n0 A.t1 148.348
R52 A A.n0 85.503
R53 A.n1 A 13.575
R54 A.n1 A 6.826
R55 A A.n1 4.266
R56 B.t1 B.t0 378.254
R57 B B.t1 253.559
R58 a_184_297.t0 a_184_297.t1 154.785
C0 VPWR X 0.26fF
C1 VPWR B 0.20fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__or3_4.ext - technology: sky130A

.subckt sky130_fd_sc_hd__or3_4 A X B C VPWR VGND VNB VPB
X0 X.t7 a_27_47.t4 VGND.t3 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 X.t3 a_27_47.t5 VPWR.t3 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 X.t6 a_27_47.t6 VGND.t2 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 VGND.t1 a_27_47.t7 X.t5 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 VPWR.t4 A.t0 a_193_297.t0 VPB.t6 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 a_193_297.t1 B.t0 a_109_297.t1 VPB.t5 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 a_27_47.t2 B.t1 VGND.t5 VNB.t5 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 VPWR.t2 a_27_47.t8 X.t2 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 VGND.t6 A.t1 a_27_47.t3 VNB.t6 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 VGND.t0 a_27_47.t9 X.t4 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 X.t1 a_27_47.t10 VPWR.t1 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 VPWR.t0 a_27_47.t11 X.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 a_109_297.t0 C.t0 a_27_47.t0 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13 VGND.t4 C.t1 a_27_47.t1 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
R0 a_27_47.t0 a_27_47.n13 284.358
R1 a_27_47.n0 a_27_47.t8 212.079
R2 a_27_47.n2 a_27_47.t10 212.079
R3 a_27_47.n5 a_27_47.t11 212.079
R4 a_27_47.n10 a_27_47.t5 212.079
R5 a_27_47.n0 a_27_47.t7 139.779
R6 a_27_47.n2 a_27_47.t6 139.779
R7 a_27_47.n5 a_27_47.t9 139.779
R8 a_27_47.n10 a_27_47.t4 139.779
R9 a_27_47.n12 a_27_47.t1 127.762
R10 a_27_47.n13 a_27_47.n10 104.481
R11 a_27_47.n4 a_27_47.n1 101.6
R12 a_27_47.n4 a_27_47.n3 76
R13 a_27_47.n7 a_27_47.n6 76
R14 a_27_47.n9 a_27_47.n8 76
R15 a_27_47.n13 a_27_47.n12 63.094
R16 a_27_47.n12 a_27_47.n11 52.237
R17 a_27_47.n7 a_27_47.n4 25.6
R18 a_27_47.n9 a_27_47.n7 25.6
R19 a_27_47.n11 a_27_47.t3 24.923
R20 a_27_47.n11 a_27_47.t2 24.923
R21 a_27_47.n13 a_27_47.n9 23.717
R22 a_27_47.n1 a_27_47.n0 13.875
R23 a_27_47.n6 a_27_47.n5 9.493
R24 a_27_47.n3 a_27_47.n2 2.19
R25 VGND.n2 VGND.t1 190.732
R26 VGND.n1 VGND.n0 115.464
R27 VGND.n16 VGND.n15 115.464
R28 VGND.n6 VGND.n5 92.5
R29 VGND.n10 VGND.n9 92.5
R30 VGND.n5 VGND.t3 24.923
R31 VGND.n9 VGND.t6 24.923
R32 VGND.n0 VGND.t2 24.923
R33 VGND.n0 VGND.t0 24.923
R34 VGND.n15 VGND.t5 24.923
R35 VGND.n15 VGND.t4 24.923
R36 VGND.n2 VGND.n1 11.464
R37 VGND.n4 VGND.n3 4.65
R38 VGND.n8 VGND.n7 4.65
R39 VGND.n12 VGND.n11 4.65
R40 VGND.n14 VGND.n13 4.65
R41 VGND.n18 VGND.n17 4.65
R42 VGND.n11 VGND.n10 1.8
R43 VGND.n17 VGND.n16 0.752
R44 VGND.n7 VGND.n6 0.4
R45 VGND.n4 VGND.n2 0.339
R46 VGND.n8 VGND.n4 0.119
R47 VGND.n12 VGND.n8 0.119
R48 VGND.n14 VGND.n12 0.119
R49 VGND.n18 VGND.n14 0.119
R50 VGND.n19 VGND.n18 0.119
R51 VGND VGND.n19 0.02
R52 X.n5 X.n3 155.184
R53 X.n5 X.n4 110.76
R54 X.n2 X.n0 91.218
R55 X.n6 X.n5 56.626
R56 X.n2 X.n1 52.818
R57 X.n3 X.t0 26.595
R58 X.n3 X.t3 26.595
R59 X.n4 X.t2 26.595
R60 X.n4 X.t1 26.595
R61 X.n0 X.t4 24.923
R62 X.n0 X.t7 24.923
R63 X.n1 X.t5 24.923
R64 X.n1 X.t6 24.923
R65 X.n6 X.n2 21.835
R66 X X.n6 2.427
R67 VNB VNB.t4 6053.91
R68 VNB.t6 VNB.t3 4593.41
R69 VNB.t2 VNB.t1 2030.77
R70 VNB.t0 VNB.t2 2030.77
R71 VNB.t3 VNB.t0 2030.77
R72 VNB.t5 VNB.t6 2030.77
R73 VNB.t4 VNB.t5 2030.77
R74 VPWR.n2 VPWR.t2 204.188
R75 VPWR.n8 VPWR.n7 193.629
R76 VPWR.n9 VPWR.n6 176.568
R77 VPWR.n1 VPWR.n0 171.981
R78 VPWR.n5 VPWR.t4 39.4
R79 VPWR.n6 VPWR.n5 27.649
R80 VPWR.n0 VPWR.t1 26.595
R81 VPWR.n0 VPWR.t0 26.595
R82 VPWR.n7 VPWR.t3 26.595
R83 VPWR.n10 VPWR.n9 6.948
R84 VPWR.n4 VPWR.n3 4.65
R85 VPWR.n9 VPWR.n8 4.116
R86 VPWR.n2 VPWR.n1 3.929
R87 VPWR.n11 VPWR.n10 2.093
R88 VPWR VPWR.n11 0.421
R89 VPWR.n4 VPWR.n2 0.318
R90 VPWR.n11 VPWR.n4 0.195
R91 VPB.t6 VPB.t3 562.305
R92 VPB.t1 VPB.t2 248.598
R93 VPB.t0 VPB.t1 248.598
R94 VPB.t3 VPB.t0 248.598
R95 VPB.t5 VPB.t6 248.598
R96 VPB.t4 VPB.t5 248.598
R97 VPB VPB.t4 189.408
R98 A.n0 A.t0 239.503
R99 A.n0 A.t1 167.203
R100 A A.n0 83.168
R101 a_193_297.t0 a_193_297.t1 53.19
R102 B.n0 B.t0 241.534
R103 B.n0 B.t1 169.234
R104 B B.n0 91.752
R105 a_109_297.t0 a_109_297.t1 53.19
R106 C.n0 C.t0 231.014
R107 C.n0 C.t1 158.714
R108 C C.n0 81.632
C0 X VGND 0.42fF
C1 B A 0.10fF
C2 VPWR X 0.63fF
C3 C B 0.10fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__or3b_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__or3b_1 A C_N X B VGND VPWR VNB VPB
X0 a_109_93.t1 C_N.t0 VGND.t1 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1 a_215_53.t3 B.t0 VGND.t2 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 VGND.t4 a_109_93.t2 a_215_53.t2 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3 VGND.t0 A.t0 a_215_53.t0 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 VPWR.t1 A.t1 a_369_297.t1 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 a_369_297.t0 B.t1 a_297_297.t1 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 X.t1 a_215_53.t4 VPWR.t2 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 a_297_297.t0 a_109_93.t3 a_215_53.t1 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 a_109_93.t0 C_N.t1 VPWR.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9 X.t0 a_215_53.t5 VGND.t3 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
R0 C_N.n0 C_N.t1 137.175
R1 C_N.n0 C_N.t0 121.108
R2 C_N C_N.n0 81.632
R3 VGND.n8 VGND.t1 167.009
R4 VGND.n3 VGND.n0 109.578
R5 VGND.n2 VGND.n1 108.015
R6 VGND.n0 VGND.t0 51.428
R7 VGND.n1 VGND.t2 38.571
R8 VGND.n1 VGND.t4 38.571
R9 VGND.n0 VGND.t3 28.378
R10 VGND.n9 VGND.n8 4.65
R11 VGND.n5 VGND.n4 4.65
R12 VGND.n7 VGND.n6 4.65
R13 VGND.n3 VGND.n2 3.797
R14 VGND.n5 VGND.n3 0.253
R15 VGND.n7 VGND.n5 0.119
R16 VGND.n9 VGND.n7 0.119
R17 VGND VGND.n9 0.022
R18 a_109_93.t0 a_109_93.n1 380.336
R19 a_109_93.n0 a_109_93.t2 183.49
R20 a_109_93.n1 a_109_93.t1 142.079
R21 a_109_93.n0 a_109_93.t3 135.29
R22 a_109_93.n1 a_109_93.n0 92.096
R23 VNB VNB.t1 6894.12
R24 VNB.t1 VNB.t2 5398.53
R25 VNB.t3 VNB.t0 2717.65
R26 VNB.t2 VNB.t3 2717.65
R27 VNB.t0 VNB.t4 2303.7
R28 B.t1 B.t0 378.254
R29 B B.t1 242.054
R30 a_215_53.n1 a_215_53.t1 486.628
R31 a_215_53.n0 a_215_53.t4 241.534
R32 a_215_53.n2 a_215_53.t2 203.671
R33 a_215_53.n0 a_215_53.t5 169.234
R34 a_215_53.n3 a_215_53.n2 106.429
R35 a_215_53.n1 a_215_53.n0 76
R36 a_215_53.n2 a_215_53.n1 63.021
R37 a_215_53.t0 a_215_53.n3 38.571
R38 a_215_53.n3 a_215_53.t3 38.571
R39 A.n0 A.t0 267.063
R40 A.n0 A.t1 148.348
R41 A A.n0 85.503
R42 A A.n1 13.187
R43 A.n1 A 5.296
R44 A.n1 A 4.654
R45 a_369_297.t0 a_369_297.t1 152.44
R46 VPWR.n1 VPWR.t0 412.018
R47 VPWR.n1 VPWR.n0 173.157
R48 VPWR.n0 VPWR.t1 96.154
R49 VPWR.n0 VPWR.t2 26.595
R50 VPWR VPWR.n1 0.04
R51 VPB.t0 VPB.t1 556.386
R52 VPB.t3 VPB.t4 290.031
R53 VPB.t2 VPB.t3 281.152
R54 VPB.t1 VPB.t2 213.084
R55 VPB VPB.t0 192.367
R56 a_297_297.t0 a_297_297.t1 98.5
R57 X X.t1 212.866
R58 X X.t0 194.174
C0 VPWR X 0.13fF
C1 VPWR B 0.34fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__or3b_2.ext - technology: sky130A

.subckt sky130_fd_sc_hd__or3b_2 A B C_N X VPWR VGND VNB VPB
X0 a_388_297.t0 A.t0 VPWR.t2 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1 VPWR.t3 C_N.t0 a_27_47.t0 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 VGND.t5 a_176_21.t4 X.t1 VNB.t5 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 X.t0 a_176_21.t5 VGND.t4 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 VPWR.t0 a_176_21.t6 X.t3 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 VGND.t3 B.t0 a_176_21.t3 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 X.t2 a_176_21.t7 VPWR.t1 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 a_176_21.t0 a_27_47.t2 a_472_297.t1 VPB.t5 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 a_472_297.t0 B.t1 a_388_297.t1 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9 a_176_21.t2 A.t1 VGND.t2 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10 a_176_21.t1 a_27_47.t3 VGND.t1 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11 VGND.t0 C_N.t1 a_27_47.t1 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
R0 A.n0 A.t1 196.548
R1 A.n0 A.t0 148.348
R2 A.n1 A.n0 76
R3  A.n1 6.818
R4 A.n1 A 1.315
R5 VPWR.n2 VPWR.n1 367.697
R6 VPWR.n2 VPWR.n0 315.909
R7 VPWR.n0 VPWR.t2 98.5
R8 VPWR.n1 VPWR.t3 96.154
R9 VPWR.n1 VPWR.t1 34.305
R10 VPWR.n0 VPWR.t0 25.61
R11 VPWR VPWR.n2 0.243
R12 a_388_297.t0 a_388_297.t1 126.642
R13 VPB.t0 VPB.t2 290.031
R14 VPB.t4 VPB.t1 287.071
R15 VPB.t3 VPB.t5 248.598
R16 VPB.t2 VPB.t3 248.598
R17 VPB.t1 VPB.t0 248.598
R18 VPB VPB.t4 189.408
R19 C_N.n0 C_N.t0 238.395
R20 C_N.n0 C_N.t1 195.015
R21 C_N.n1 C_N.n0 76
R22  C_N.n1 10.729
R23 C_N.n1 C_N 2.07
R24 a_27_47.t0 a_27_47.n1 377.117
R25 a_27_47.n1 a_27_47.n0 254.419
R26 a_27_47.n1 a_27_47.t1 242.404
R27 a_27_47.n0 a_27_47.t3 196.548
R28 a_27_47.n0 a_27_47.t2 148.348
R29 a_176_21.t0 a_176_21.n5 419.768
R30 a_176_21.n0 a_176_21.t6 212.079
R31 a_176_21.n1 a_176_21.t7 212.079
R32 a_176_21.n4 a_176_21.n2 145.068
R33 a_176_21.n0 a_176_21.t4 139.779
R34 a_176_21.n1 a_176_21.t5 139.779
R35 a_176_21.n5 a_176_21.t1 137.847
R36 a_176_21.n4 a_176_21.n3 112.829
R37 a_176_21.n2 a_176_21.n1 59.154
R38 a_176_21.n5 a_176_21.n4 57.719
R39 a_176_21.n3 a_176_21.t3 38.571
R40 a_176_21.n3 a_176_21.t2 38.571
R41 a_176_21.n2 a_176_21.n0 2.19
R42 X.n2 X.n0 375.351
R43 X.n2 X.n1 92.5
R44 X.n0 X.t3 26.595
R45 X.n0 X.t2 26.595
R46 X.n1 X.t1 24.923
R47 X.n1 X.t0 24.923
R48 X X.n2 0.182
R49 VGND.n2 VGND.n1 116.217
R50 VGND.n7 VGND.n6 116.217
R51 VGND.n3 VGND.n0 111.57
R52 VGND.n1 VGND.t2 52.857
R53 VGND.n6 VGND.t4 44
R54 VGND.n0 VGND.t1 38.571
R55 VGND.n0 VGND.t3 38.571
R56 VGND.n6 VGND.t0 38.571
R57 VGND.n1 VGND.t5 28.315
R58 VGND.n5 VGND.n4 4.65
R59 VGND.n9 VGND.n8 4.65
R60 VGND.n3 VGND.n2 4.441
R61 VGND.n8 VGND.n7 0.752
R62 VGND.n5 VGND.n3 0.205
R63 VGND.n9 VGND.n5 0.119
R64 VGND.n10 VGND.n9 0.119
R65 VGND VGND.n10 0.022
R66 VNB VNB.t0 6470.59
R67 VNB.t3 VNB.t1 2717.65
R68 VNB.t2 VNB.t3 2717.65
R69 VNB.t5 VNB.t2 2327.87
R70 VNB.t0 VNB.t4 2303.7
R71 VNB.t4 VNB.t5 2030.77
R72 B.t1 B.t0 392.026
R73 B B.t1 249.118
R74  B 24.533
R75 a_472_297.t0 a_472_297.t1 126.642
C0 VPWR B 0.15fF
C1 X VGND 0.13fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__or3b_4.ext - technology: sky130A

.subckt sky130_fd_sc_hd__or3b_4 A B C_N X VGND VPWR VNB VPB
X0 a_176_21.t3 a_27_47.t2 a_626_297.t1 VPB.t7 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_626_297.t0 B.t0 a_542_297.t0 VPB.t5 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 VPWR.t4 C_N.t0 a_27_47.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3 VGND.t4 a_176_21.t4 X.t7 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 a_542_297.t1 A.t0 VPWR.t5 VPB.t6 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 VPWR.t3 a_176_21.t5 X.t3 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 X.t2 a_176_21.t6 VPWR.t2 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 X.t6 a_176_21.t7 VGND.t3 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 X.t5 a_176_21.t8 VGND.t2 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 a_176_21.t1 A.t1 VGND.t6 VNB.t6 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 VPWR.t1 a_176_21.t9 X.t1 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 X.t0 a_176_21.t10 VPWR.t0 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 a_176_21.t2 a_27_47.t3 VGND.t7 VNB.t7 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 VGND.t1 a_176_21.t11 X.t4 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14 VGND.t0 B.t1 a_176_21.t0 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X15 VGND.t5 C_N.t1 a_27_47.t1 VNB.t5 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
R0 a_27_47.t0 a_27_47.n1 377.117
R1 a_27_47.n1 a_27_47.n0 320.719
R2 a_27_47.n1 a_27_47.t1 242.404
R3 a_27_47.n0 a_27_47.t2 241.534
R4 a_27_47.n0 a_27_47.t3 169.234
R5 a_626_297.t0 a_626_297.t1 65.01
R6 a_176_21.t3 a_176_21.n9 635.666
R7 a_176_21.n5 a_176_21.t5 212.079
R8 a_176_21.n1 a_176_21.t6 212.079
R9 a_176_21.n3 a_176_21.t9 212.079
R10 a_176_21.n2 a_176_21.t10 212.079
R11 a_176_21.n5 a_176_21.t11 139.779
R12 a_176_21.n1 a_176_21.t8 139.779
R13 a_176_21.n3 a_176_21.t4 139.779
R14 a_176_21.n2 a_176_21.t7 139.779
R15 a_176_21.n9 a_176_21.t2 124.199
R16 a_176_21.n8 a_176_21.n0 106.429
R17 a_176_21.n7 a_176_21.n6 76
R18 a_176_21.n9 a_176_21.n8 68.636
R19 a_176_21.n8 a_176_21.n7 65.459
R20 a_176_21.n3 a_176_21.n2 61.345
R21 a_176_21.n7 a_176_21.n4 59.577
R22 a_176_21.n4 a_176_21.n3 31.695
R23 a_176_21.n0 a_176_21.t0 24.923
R24 a_176_21.n0 a_176_21.t1 24.923
R25 a_176_21.n4 a_176_21.n1 18.798
R26 a_176_21.n6 a_176_21.n5 13.875
R27 VPB.t0 VPB.t1 287.071
R28 VPB.t5 VPB.t7 284.112
R29 VPB.t6 VPB.t5 248.598
R30 VPB.t4 VPB.t6 248.598
R31 VPB.t3 VPB.t4 248.598
R32 VPB.t2 VPB.t3 248.598
R33 VPB.t1 VPB.t2 248.598
R34 VPB VPB.t0 189.408
R35 B.n0 B.t0 241.534
R36 B.n0 B.t1 169.234
R37 B.n1 B.n0 76
R38  B.n1 11.767
R39 B.n1 B 2.27
R40 a_542_297.t0 a_542_297.t1 53.19
R41 C_N.n0 C_N.t0 238.395
R42 C_N.n0 C_N.t1 195.015
R43 C_N.n1 C_N.n0 76
R44  C_N.n1 10.729
R45 C_N.n1 C_N 2.07
R46 VPWR.n7 VPWR.n6 364.437
R47 VPWR.n3 VPWR.n2 311.884
R48 VPWR.n1 VPWR.n0 308.984
R49 VPWR.n6 VPWR.t4 96.154
R50 VPWR.n6 VPWR.t0 34.305
R51 VPWR.n2 VPWR.t5 26.595
R52 VPWR.n2 VPWR.t3 26.595
R53 VPWR.n0 VPWR.t2 26.595
R54 VPWR.n0 VPWR.t1 26.595
R55 VPWR.n5 VPWR.n4 4.65
R56 VPWR.n8 VPWR.n7 3.989
R57 VPWR.n3 VPWR.n1 3.847
R58 VPWR.n5 VPWR.n3 0.259
R59 VPWR.n8 VPWR.n5 0.136
R60 VPWR VPWR.n8 0.123
R61 X X.n0 293.173
R62 X.n5 X.n1 292.5
R63 X.n4 X.n2 171.133
R64 X.n5 X.n4 55.829
R65 X.n4 X.n3 49.327
R66 X X.n5 37.052
R67 X.n1 X.t1 26.595
R68 X.n1 X.t0 26.595
R69 X.n0 X.t3 26.595
R70 X.n0 X.t2 26.595
R71 X.n3 X.t7 24.923
R72 X.n3 X.t6 24.923
R73 X.n2 X.t4 24.923
R74 X.n2 X.t5 24.923
R75 VGND.n7 VGND.n6 116.217
R76 VGND.n13 VGND.n12 116.217
R77 VGND.n3 VGND.n0 108.748
R78 VGND.n2 VGND.n1 108.015
R79 VGND.n12 VGND.t5 45.714
R80 VGND.n12 VGND.t3 36.857
R81 VGND.n0 VGND.t7 36
R82 VGND.n0 VGND.t0 24.923
R83 VGND.n1 VGND.t6 24.923
R84 VGND.n1 VGND.t1 24.923
R85 VGND.n6 VGND.t2 24.923
R86 VGND.n6 VGND.t4 24.923
R87 VGND.n14 VGND.n13 5.276
R88 VGND.n5 VGND.n4 4.65
R89 VGND.n9 VGND.n8 4.65
R90 VGND.n11 VGND.n10 4.65
R91 VGND.n3 VGND.n2 3.932
R92 VGND.n8 VGND.n7 1.882
R93 VGND.n5 VGND.n3 0.274
R94 VGND.n14 VGND.n11 0.132
R95 VGND VGND.n14 0.127
R96 VGND.n9 VGND.n5 0.119
R97 VGND.n11 VGND.n9 0.119
R98 VNB VNB.t5 6438.23
R99 VNB.t0 VNB.t7 2320.88
R100 VNB.t5 VNB.t3 2303.7
R101 VNB.t6 VNB.t0 2030.77
R102 VNB.t1 VNB.t6 2030.77
R103 VNB.t2 VNB.t1 2030.77
R104 VNB.t4 VNB.t2 2030.77
R105 VNB.t3 VNB.t4 2030.77
R106 A.n0 A.t0 241.534
R107 A.n0 A.t1 169.234
R108 A A.n0 101.502
C0 X VGND 0.29fF
C1 A B 0.15fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__or4_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__or4_1 C A X B D VPWR VGND VNB VPB
X0 a_27_297.t0 B.t0 VGND.t0 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1 a_27_297.t1 D.t0 VGND.t1 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 a_277_297.t0 B.t1 a_205_297.t0 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3 VPWR.t1 A.t0 a_277_297.t1 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 X.t1 a_27_297.t5 VGND.t4 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 a_205_297.t1 C.t0 a_109_297.t1 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 X.t0 a_27_297.t6 VPWR.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 VGND.t3 C.t1 a_27_297.t4 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 a_109_297.t0 D.t1 a_27_297.t2 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9 VGND.t2 A.t1 a_27_297.t3 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
R0 B.t1 B.t0 618.106
R1 B B.t1 253.559
R2 VGND.n6 VGND.t1 150.464
R3 VGND.n3 VGND.n0 109.393
R4 VGND.n2 VGND.n1 108.015
R5 VGND.n0 VGND.t2 52.857
R6 VGND.n1 VGND.t0 38.571
R7 VGND.n1 VGND.t3 38.571
R8 VGND.n0 VGND.t4 27.568
R9 VGND.n7 VGND.n6 4.65
R10 VGND.n5 VGND.n4 4.65
R11 VGND.n3 VGND.n2 3.797
R12 VGND.n5 VGND.n3 0.253
R13 VGND.n7 VGND.n5 0.119
R14 VGND VGND.n7 0.02
R15 a_27_297.n1 a_27_297.t2 523.889
R16 a_27_297.n0 a_27_297.t6 240.999
R17 a_27_297.n3 a_27_297.n2 171.934
R18 a_27_297.n0 a_27_297.t5 168.699
R19 a_27_297.n4 a_27_297.n3 106.429
R20 a_27_297.n1 a_27_297.n0 76
R21 a_27_297.n3 a_27_297.n1 63.539
R22 a_27_297.n2 a_27_297.t4 47.142
R23 a_27_297.n2 a_27_297.t1 47.142
R24 a_27_297.n4 a_27_297.t3 38.571
R25 a_27_297.t0 a_27_297.n4 38.571
R26 VNB VNB.t2 7214.71
R27 VNB.t2 VNB.t4 3105.88
R28 VNB.t1 VNB.t3 2717.65
R29 VNB.t4 VNB.t1 2717.65
R30 VNB.t3 VNB.t0 2327.87
R31 D.n0 D.t0 186.028
R32 D.n0 D.t1 137.828
R33 D D.n0 78.011
R34 a_205_297.t0 a_205_297.t1 98.5
R35 a_277_297.t0 a_277_297.t1 154.785
R36 VPB.t2 VPB.t0 290.031
R37 VPB.t1 VPB.t2 284.112
R38 VPB.t3 VPB.t4 284.112
R39 VPB.t4 VPB.t1 213.084
R40 VPB VPB.t3 189.408
R41 A.n0 A.t1 196.548
R42 A.n0 A.t0 148.348
R43 A A.n0 85.309
R44 VPWR VPWR.n0 173.077
R45 VPWR.n0 VPWR.t1 96.154
R46 VPWR.n0 VPWR.t0 26.595
R47 X X.t0 214.087
R48 X X.t1 194.571
R49 C.n0 C.t1 196.548
R50 C.n0 C.t0 148.348
R51 C.n1 C.n0 76
R52 C C.n1 5.78
R53 C.n1 C 3.716
R54 a_109_297.t0 a_109_297.t1 154.785
C0 VPWR B 0.26fF
C1 X VPWR 0.13fF
C2 D C 0.12fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__or4_2.ext - technology: sky130A

.subckt sky130_fd_sc_hd__or4_2 C A X B D VPWR VGND VNB VPB
X0 a_27_297.t4 B.t0 VGND.t5 VNB.t5 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1 a_27_297.t1 D.t0 VGND.t1 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 a_277_297.t1 B.t1 a_205_297.t1 VPB.t5 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3 VPWR.t2 A.t0 a_277_297.t0 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 X.t3 a_27_297.t5 VGND.t3 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 a_205_297.t0 C.t0 a_109_297.t1 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 VPWR.t1 a_27_297.t6 X.t1 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 VGND.t4 a_27_297.t7 X.t2 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 X.t0 a_27_297.t8 VPWR.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 VGND.t0 C.t1 a_27_297.t0 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10 a_109_297.t0 D.t1 a_27_297.t2 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11 VGND.t2 A.t1 a_27_297.t3 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
R0 B.t1 B.t0 378.254
R1 B B.t1 253.559
R2 VGND.n10 VGND.t1 150.175
R3 VGND.n2 VGND.t4 112.172
R4 VGND.n6 VGND.n5 108.015
R5 VGND.n1 VGND.n0 105.973
R6 VGND.n0 VGND.t2 52.857
R7 VGND.n5 VGND.t5 38.571
R8 VGND.n5 VGND.t0 38.571
R9 VGND.n0 VGND.t3 27.568
R10 VGND.n11 VGND.n10 4.65
R11 VGND.n4 VGND.n3 4.65
R12 VGND.n7 VGND.n6 4.65
R13 VGND.n9 VGND.n8 4.65
R14 VGND.n2 VGND.n1 3.837
R15 VGND.n4 VGND.n2 0.271
R16 VGND.n7 VGND.n4 0.119
R17 VGND.n9 VGND.n7 0.119
R18 VGND.n11 VGND.n9 0.119
R19 VGND VGND.n11 0.02
R20 a_27_297.n3 a_27_297.t2 523.633
R21 a_27_297.n1 a_27_297.t6 212.079
R22 a_27_297.n2 a_27_297.t8 212.079
R23 a_27_297.n5 a_27_297.n4 171.934
R24 a_27_297.n1 a_27_297.t7 139.779
R25 a_27_297.n2 a_27_297.t5 139.779
R26 a_27_297.n4 a_27_297.n0 106.429
R27 a_27_297.n3 a_27_297.n2 79.651
R28 a_27_297.n4 a_27_297.n3 63.397
R29 a_27_297.n2 a_27_297.n1 61.345
R30 a_27_297.t0 a_27_297.n5 47.142
R31 a_27_297.n5 a_27_297.t1 47.142
R32 a_27_297.n0 a_27_297.t3 38.571
R33 a_27_297.n0 a_27_297.t4 38.571
R34 VNB VNB.t3 7214.71
R35 VNB.t3 VNB.t2 3105.88
R36 VNB.t5 VNB.t4 2717.65
R37 VNB.t2 VNB.t5 2717.65
R38 VNB.t4 VNB.t1 2327.87
R39 VNB.t1 VNB.t0 2030.77
R40 D.n0 D.t0 186.028
R41 D.n0 D.t1 137.828
R42 D D.n0 77.983
R43 a_205_297.t0 a_205_297.t1 98.5
R44 a_277_297.t0 a_277_297.t1 154.785
R45 VPB.t4 VPB.t0 290.031
R46 VPB.t5 VPB.t4 284.112
R47 VPB.t2 VPB.t3 284.112
R48 VPB.t0 VPB.t1 248.598
R49 VPB.t3 VPB.t5 213.084
R50 VPB VPB.t2 189.408
R51 A.n0 A.t1 196.548
R52 A.n0 A.t0 148.348
R53 A A.n0 85.503
R54 VPWR.n1 VPWR.n0 172.464
R55 VPWR.n1 VPWR.t1 171.472
R56 VPWR.n0 VPWR.t2 96.154
R57 VPWR.n0 VPWR.t0 26.595
R58 VPWR VPWR.n1 0.606
R59 X X.n1 169.251
R60 X X.n0 152.895
R61 X.n0 X.t1 26.595
R62 X.n0 X.t0 26.595
R63 X.n1 X.t2 24.923
R64 X.n1 X.t3 24.923
R65 C.n0 C.t1 196.548
R66 C.n0 C.t0 148.348
R67 C.n1 C.n0 76
R68 C C.n1 5.78
R69 C.n1 C 3.716
R70 a_109_297.t0 a_109_297.t1 154.785
C0 VPWR X 0.24fF
C1 D C 0.12fF
C2 VPWR B 0.26fF
C3 X VGND 0.11fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__or4_4.ext - technology: sky130A

.subckt sky130_fd_sc_hd__or4_4 B C A D X VPWR VGND VNB VPB
X0 VPWR.t0 A.t0 a_304_297.t0 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_304_297.t1 B.t0 a_220_297.t1 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 VGND.t7 C.t0 a_32_297.t4 VNB.t7 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 a_220_297.t0 C.t1 a_114_297.t1 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 a_32_297.t0 D.t0 VGND.t0 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 a_32_297.t3 B.t1 VGND.t6 VNB.t6 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 VPWR.t1 a_32_297.t5 X.t3 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 X.t2 a_32_297.t6 VPWR.t2 VPB.t5 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 VGND.t5 A.t1 a_32_297.t2 VNB.t5 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 VPWR.t3 a_32_297.t7 X.t1 VPB.t6 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 X.t7 a_32_297.t8 VGND.t4 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 X.t6 a_32_297.t9 VGND.t3 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 X.t0 a_32_297.t10 VPWR.t4 VPB.t7 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13 a_114_297.t0 D.t1 a_32_297.t1 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14 VGND.t2 a_32_297.t11 X.t5 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X15 VGND.t1 a_32_297.t12 X.t4 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
R0 A.n0 A.t0 241.534
R1 A.n0 A.t1 169.234
R2 A A.n0 101.599
R3 a_304_297.t0 a_304_297.t1 53.19
R4 VPWR.n4 VPWR.t1 202.594
R5 VPWR.n1 VPWR.n0 171.981
R6 VPWR.n3 VPWR.n2 171.981
R7 VPWR.n0 VPWR.t4 37.43
R8 VPWR.n0 VPWR.t0 37.43
R9 VPWR.n2 VPWR.t2 26.595
R10 VPWR.n2 VPWR.t3 26.595
R11 VPWR.n6 VPWR.n5 4.65
R12 VPWR.n7 VPWR.n1 4.075
R13 VPWR.n4 VPWR.n3 3.837
R14 VPWR VPWR.n7 0.485
R15 VPWR.n6 VPWR.n4 0.243
R16 VPWR.n7 VPWR.n6 0.136
R17 VPB.t2 VPB.t7 313.707
R18 VPB.t1 VPB.t0 313.707
R19 VPB.t5 VPB.t4 248.598
R20 VPB.t6 VPB.t5 248.598
R21 VPB.t7 VPB.t6 248.598
R22 VPB.t3 VPB.t2 248.598
R23 VPB.t0 VPB.t3 248.598
R24 VPB VPB.t1 210.124
R25 B.n0 B.t0 241.534
R26 B.n0 B.t1 169.234
R27 B B.n0 107.667
R28 a_220_297.t0 a_220_297.t1 53.19
R29 C.n0 C.t1 241.534
R30 C.n0 C.t0 169.234
R31 C C.n0 116.669
R32 a_32_297.n2 a_32_297.t5 212.079
R33 a_32_297.n4 a_32_297.t6 212.079
R34 a_32_297.n7 a_32_297.t7 212.079
R35 a_32_297.n10 a_32_297.t10 212.079
R36 a_32_297.t1 a_32_297.n14 209.754
R37 a_32_297.n2 a_32_297.t12 139.779
R38 a_32_297.n4 a_32_297.t9 139.779
R39 a_32_297.n7 a_32_297.t11 139.779
R40 a_32_297.n10 a_32_297.t8 139.779
R41 a_32_297.n14 a_32_297.n0 104.923
R42 a_32_297.n13 a_32_297.n1 104.923
R43 a_32_297.n6 a_32_297.n3 101.6
R44 a_32_297.n13 a_32_297.n12 79.057
R45 a_32_297.n6 a_32_297.n5 76
R46 a_32_297.n9 a_32_297.n8 76
R47 a_32_297.n12 a_32_297.n11 76
R48 a_32_297.n14 a_32_297.n13 65.505
R49 a_32_297.n0 a_32_297.t0 39.692
R50 a_32_297.n0 a_32_297.t4 30.461
R51 a_32_297.n3 a_32_297.n2 26.29
R52 a_32_297.n9 a_32_297.n6 25.6
R53 a_32_297.n12 a_32_297.n9 25.6
R54 a_32_297.n1 a_32_297.t2 24.923
R55 a_32_297.n1 a_32_297.t3 24.923
R56 a_32_297.n5 a_32_297.n4 14.606
R57 a_32_297.n11 a_32_297.n10 8.763
R58 a_32_297.n8 a_32_297.n7 2.921
R59 VGND.n0 VGND.t1 195.432
R60 VGND.n17 VGND.t0 178.619
R61 VGND.n2 VGND.n1 115.464
R62 VGND.n13 VGND.n12 108.015
R63 VGND.n8 VGND.n7 105.973
R64 VGND.n7 VGND.t5 43.384
R65 VGND.n7 VGND.t4 26.769
R66 VGND.n1 VGND.t3 24.923
R67 VGND.n1 VGND.t2 24.923
R68 VGND.n12 VGND.t6 24.923
R69 VGND.n12 VGND.t7 24.923
R70 VGND.n18 VGND.n17 4.65
R71 VGND.n4 VGND.n3 4.65
R72 VGND.n6 VGND.n5 4.65
R73 VGND.n9 VGND.n8 4.65
R74 VGND.n11 VGND.n10 4.65
R75 VGND.n14 VGND.n13 4.65
R76 VGND.n16 VGND.n15 4.65
R77 VGND.n3 VGND.n2 2.635
R78 VGND.n4 VGND.n0 0.981
R79 VGND.n6 VGND.n4 0.119
R80 VGND.n9 VGND.n6 0.119
R81 VGND.n11 VGND.n9 0.119
R82 VGND.n14 VGND.n11 0.119
R83 VGND.n16 VGND.n14 0.119
R84 VGND.n18 VGND.n16 0.119
R85 VGND VGND.n18 0.023
R86 VNB VNB.t0 6223.14
R87 VNB.t5 VNB.t4 2562.64
R88 VNB.t0 VNB.t7 2562.64
R89 VNB.t3 VNB.t1 2030.77
R90 VNB.t2 VNB.t3 2030.77
R91 VNB.t4 VNB.t2 2030.77
R92 VNB.t6 VNB.t5 2030.77
R93 VNB.t7 VNB.t6 2030.77
R94 a_114_297.t0 a_114_297.t1 74.86
R95 D.n0 D.t1 231.014
R96 D.n0 D.t0 158.714
R97 D D.n0 78.47
R98  D 15.27
R99 X.n5 X.n3 155.184
R100 X.n2 X.n0 145.662
R101 X.n5 X.n4 110.76
R102 X.n6 X.n5 55.947
R103 X.n2 X.n1 52.624
R104 X.n3 X.t1 26.595
R105 X.n3 X.t0 26.595
R106 X.n4 X.t3 26.595
R107 X.n4 X.t2 26.595
R108 X.n0 X.t5 24.923
R109 X.n0 X.t7 24.923
R110 X.n1 X.t4 24.923
R111 X.n1 X.t6 24.923
R112 X.n6 X.n2 14.222
R113 X X.n6 2.612
C0 X VGND 0.40fF
C1 B A 0.13fF
C2 VPWR X 0.66fF
C3 B VPWR 0.10fF
C4 C B 0.25fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__or4b_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__or4b_1 B D_N A X C VPWR VGND VNB VPB
X0 X.t0 a_215_297.t5 VPWR.t2 VPB.t5 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_109_53.t1 D_N.t0 VGND.t1 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 a_215_297.t3 a_109_53.t2 VGND.t4 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3 X.t1 a_215_297.t6 VGND.t5 VNB.t5 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 a_392_297.t0 C.t0 a_297_297.t0 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 a_465_297.t1 B.t0 a_392_297.t1 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 a_215_297.t2 B.t1 VGND.t3 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7 VPWR.t0 A.t0 a_465_297.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 a_297_297.t1 a_109_53.t3 a_215_297.t4 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9 a_109_53.t0 D_N.t1 VPWR.t1 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10 VGND.t2 C.t1 a_215_297.t1 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11 VGND.t0 A.t1 a_215_297.t0 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
R0 a_215_297.n1 a_215_297.t4 521.865
R1 a_215_297.n0 a_215_297.t5 241.534
R2 a_215_297.n3 a_215_297.n2 170.052
R3 a_215_297.n0 a_215_297.t6 169.234
R4 a_215_297.n4 a_215_297.n3 106.429
R5 a_215_297.n1 a_215_297.n0 76
R6 a_215_297.n3 a_215_297.n1 63.397
R7 a_215_297.n2 a_215_297.t3 47.142
R8 a_215_297.n2 a_215_297.t1 40
R9 a_215_297.t0 a_215_297.n4 38.571
R10 a_215_297.n4 a_215_297.t2 38.571
R11 VPWR.n1 VPWR.t1 397.348
R12 VPWR.n1 VPWR.n0 173.272
R13 VPWR.n0 VPWR.t0 96.154
R14 VPWR.n0 VPWR.t2 26.595
R15 VPWR VPWR.n1 0.042
R16 X X.t0 212.866
R17 X X.t1 194.174
R18 VPB.t3 VPB.t4 556.386
R19 VPB.t0 VPB.t5 290.031
R20 VPB.t4 VPB.t1 281.152
R21 VPB.t2 VPB.t0 269.314
R22 VPB.t1 VPB.t2 216.043
R23 VPB VPB.t3 189.408
R24 D_N.n0 D_N.t0 185.168
R25 D_N.n0 D_N.t1 136.968
R26 D_N D_N.n0 78.07
R27 VGND.n6 VGND.t4 150.464
R28 VGND.n10 VGND.t1 149.894
R29 VGND.n3 VGND.n0 109.388
R30 VGND.n2 VGND.n1 108.015
R31 VGND.n0 VGND.t0 52.857
R32 VGND.n1 VGND.t3 38.571
R33 VGND.n1 VGND.t2 38.571
R34 VGND.n0 VGND.t5 27.568
R35 VGND.n11 VGND.n10 4.65
R36 VGND.n5 VGND.n4 4.65
R37 VGND.n7 VGND.n6 4.65
R38 VGND.n9 VGND.n8 4.65
R39 VGND.n3 VGND.n2 3.805
R40 VGND.n5 VGND.n3 0.254
R41 VGND.n7 VGND.n5 0.119
R42 VGND.n9 VGND.n7 0.119
R43 VGND.n11 VGND.n9 0.119
R44 VGND VGND.n11 0.02
R45 a_109_53.t0 a_109_53.n1 376.887
R46 a_109_53.n0 a_109_53.t2 184.572
R47 a_109_53.n1 a_109_53.t1 156.932
R48 a_109_53.n0 a_109_53.t3 136.372
R49 a_109_53.n1 a_109_53.n0 93.454
R50 VNB VNB.t2 7214.71
R51 VNB.t2 VNB.t1 6082.35
R52 VNB.t1 VNB.t3 2944.12
R53 VNB.t4 VNB.t0 2717.65
R54 VNB.t3 VNB.t4 2717.65
R55 VNB.t0 VNB.t5 2327.87
R56 C.n0 C.t1 196.548
R57 C.n0 C.t0 148.348
R58 C.n1 C.n0 76
R59 C.n1 C 6.296
R60 C C.n1 3.2
R61 a_297_297.t0 a_297_297.t1 152.44
R62 a_392_297.t0 a_392_297.t1 100.845
R63 B.t0 B.t1 382.907
R64 B B.t0 242.315
R65 a_465_297.t0 a_465_297.t1 143.059
R66 A.n0 A.t1 196.548
R67 A.n0 A.t0 148.348
R68 A A.n0 85.503
C0 VPWR B 0.35fF
C1 VPWR X 0.13fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__or4b_2.ext - technology: sky130A

.subckt sky130_fd_sc_hd__or4b_2 C A X B D_N VPWR VGND VNB VPB
X0 a_176_21.t0 C.t0 VGND.t0 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1 VGND.t4 D_N.t0 a_27_53.t0 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 VGND.t1 a_176_21.t5 X.t1 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 X.t0 a_176_21.t6 VGND.t2 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 VPWR.t3 a_176_21.t7 X.t3 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 a_555_297.t0 C.t1 a_483_297.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 a_176_21.t2 a_27_53.t2 a_555_297.t1 VPB.t6 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7 X.t2 a_176_21.t8 VPWR.t2 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 a_387_297.t0 A.t0 VPWR.t1 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9 a_483_297.t1 B.t0 a_387_297.t1 VPB.t5 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10 VGND.t6 B.t1 a_176_21.t4 VNB.t6 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11 VGND.t5 a_27_53.t3 a_176_21.t3 VNB.t5 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12 VPWR.t0 D_N.t1 a_27_53.t1 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13 a_176_21.t1 A.t1 VGND.t3 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
R0 C.n0 C.t0 196.548
R1 C.n0 C.t1 148.348
R2 C C.n0 85.28
R3 VGND.n2 VGND.t5 154.337
R4 VGND.n11 VGND.n10 116.217
R5 VGND.n1 VGND.n0 108.015
R6 VGND.n6 VGND.n5 105.973
R7 VGND.n5 VGND.t3 52.857
R8 VGND.n10 VGND.t4 48.571
R9 VGND.n0 VGND.t0 38.571
R10 VGND.n0 VGND.t6 38.571
R11 VGND.n10 VGND.t2 31.236
R12 VGND.n5 VGND.t1 26.95
R13 VGND.n12 VGND.n11 6.029
R14 VGND.n4 VGND.n3 4.65
R15 VGND.n7 VGND.n6 4.65
R16 VGND.n9 VGND.n8 4.65
R17 VGND.n2 VGND.n1 3.765
R18 VGND.n4 VGND.n2 0.268
R19 VGND.n12 VGND.n9 0.132
R20 VGND VGND.n12 0.127
R21 VGND.n7 VGND.n4 0.119
R22 VGND.n9 VGND.n7 0.119
R23 a_176_21.n3 a_176_21.t2 518.819
R24 a_176_21.n2 a_176_21.t7 212.079
R25 a_176_21.n1 a_176_21.t8 212.079
R26 a_176_21.n5 a_176_21.n4 180.216
R27 a_176_21.n2 a_176_21.t5 139.779
R28 a_176_21.n1 a_176_21.t6 139.779
R29 a_176_21.n4 a_176_21.n0 112.452
R30 a_176_21.n3 a_176_21.n2 76
R31 a_176_21.n2 a_176_21.n1 61.345
R32 a_176_21.n4 a_176_21.n3 60.866
R33 a_176_21.n0 a_176_21.t4 55.714
R34 a_176_21.n0 a_176_21.t1 38.571
R35 a_176_21.n5 a_176_21.t3 38.571
R36 a_176_21.t0 a_176_21.n5 38.571
R37 VNB VNB.t4 6373.98
R38 VNB.t1 VNB.t6 3105.88
R39 VNB.t0 VNB.t5 2717.65
R40 VNB.t6 VNB.t0 2717.65
R41 VNB.t3 VNB.t1 2303.7
R42 VNB.t4 VNB.t2 2302.67
R43 VNB.t2 VNB.t3 2030.77
R44 D_N.n0 D_N.t0 186.028
R45 D_N.n0 D_N.t1 137.828
R46 D_N D_N.n0 79.911
R47 a_27_53.n0 a_27_53.t2 440.601
R48 a_27_53.t2 a_27_53.t3 392.026
R49 a_27_53.n0 a_27_53.t1 372.663
R50 a_27_53.t0 a_27_53.n0 226.1
R51 X.n2 X.n0 415.341
R52 X.n2 X.n1 92.5
R53 X.n0 X.t3 26.595
R54 X.n0 X.t2 26.595
R55 X.n1 X.t1 24.923
R56 X.n1 X.t0 24.923
R57 X X.n2 4.114
R58 VPWR.n2 VPWR.n0 433.174
R59 VPWR.n2 VPWR.n1 430.393
R60 VPWR.n1 VPWR.t0 96.154
R61 VPWR.n0 VPWR.t1 96.154
R62 VPWR.n0 VPWR.t3 27.807
R63 VPWR.n1 VPWR.t2 27.709
R64 VPWR VPWR.n2 0.194
R65 VPB.t4 VPB.t2 287.071
R66 VPB.t1 VPB.t3 287.071
R67 VPB.t0 VPB.t6 284.112
R68 VPB.t2 VPB.t5 284.112
R69 VPB.t3 VPB.t4 248.598
R70 VPB.t5 VPB.t0 213.084
R71 VPB VPB.t1 189.408
R72 a_483_297.t0 a_483_297.t1 98.5
R73 a_555_297.t0 a_555_297.t1 154.785
R74 A.n0 A.t1 196.548
R75 A.n0 A.t0 148.348
R76 A A.n0 80.16
R77 a_387_297.t0 a_387_297.t1 154.785
R78 B.t0 B.t1 392.026
R79 B B.t0 250.014
C0 X VGND 0.12fF
C1 VPWR B 0.11fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__or4b_4.ext - technology: sky130A

.subckt sky130_fd_sc_hd__or4b_4 D_N B C A X VGND VPWR VNB VPB
X0 X.t3 a_215_297.t5 VPWR.t3 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 VGND.t3 a_215_297.t6 X.t7 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 VPWR.t2 a_215_297.t7 X.t2 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 a_109_93.t0 D_N.t0 VGND.t5 VNB.t5 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 a_215_297.t0 a_109_93.t2 VGND.t4 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 VGND.t8 C.t0 a_215_297.t4 VNB.t8 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 VGND.t6 A.t0 a_215_297.t2 VNB.t6 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 X.t1 a_215_297.t8 VPWR.t1 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 a_215_297.t3 B.t0 VGND.t7 VNB.t7 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 a_109_93.t1 D_N.t1 VPWR.t4 VPB.t5 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10 VPWR.t5 A.t1 a_487_297.t0 VPB.t6 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 VGND.t2 a_215_297.t9 X.t6 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 a_487_297.t1 B.t1 a_403_297.t1 VPB.t7 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13 a_403_297.t0 C.t1 a_297_297.t0 VPB.t8 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14 VPWR.t0 a_215_297.t10 X.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 X.t5 a_215_297.t11 VGND.t1 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X16 X.t4 a_215_297.t12 VGND.t0 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X17 a_297_297.t1 a_109_93.t3 a_215_297.t1 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
R0 a_215_297.t1 a_215_297.n14 212.821
R1 a_215_297.n2 a_215_297.t10 212.079
R2 a_215_297.n4 a_215_297.t5 212.079
R3 a_215_297.n7 a_215_297.t7 212.079
R4 a_215_297.n10 a_215_297.t8 212.079
R5 a_215_297.n2 a_215_297.t6 139.779
R6 a_215_297.n4 a_215_297.t12 139.779
R7 a_215_297.n7 a_215_297.t9 139.779
R8 a_215_297.n10 a_215_297.t11 139.779
R9 a_215_297.n14 a_215_297.n0 104.923
R10 a_215_297.n13 a_215_297.n1 104.923
R11 a_215_297.n6 a_215_297.n3 101.6
R12 a_215_297.n13 a_215_297.n12 79.057
R13 a_215_297.n6 a_215_297.n5 76
R14 a_215_297.n9 a_215_297.n8 76
R15 a_215_297.n12 a_215_297.n11 76
R16 a_215_297.n14 a_215_297.n13 65.505
R17 a_215_297.n0 a_215_297.t0 39.692
R18 a_215_297.n0 a_215_297.t4 30.461
R19 a_215_297.n3 a_215_297.n2 26.29
R20 a_215_297.n9 a_215_297.n6 25.6
R21 a_215_297.n12 a_215_297.n9 25.6
R22 a_215_297.n1 a_215_297.t2 24.923
R23 a_215_297.n1 a_215_297.t3 24.923
R24 a_215_297.n5 a_215_297.n4 14.606
R25 a_215_297.n11 a_215_297.n10 8.763
R26 a_215_297.n8 a_215_297.n7 2.921
R27 VPWR.n18 VPWR.t4 375.021
R28 VPWR.n2 VPWR.t0 202.585
R29 VPWR.n6 VPWR.n5 171.981
R30 VPWR.n1 VPWR.n0 171.981
R31 VPWR.n5 VPWR.t1 37.43
R32 VPWR.n5 VPWR.t5 37.43
R33 VPWR.n0 VPWR.t3 26.595
R34 VPWR.n0 VPWR.t2 26.595
R35 VPWR.n4 VPWR.n3 4.65
R36 VPWR.n7 VPWR.n6 4.65
R37 VPWR.n9 VPWR.n8 4.65
R38 VPWR.n11 VPWR.n10 4.65
R39 VPWR.n13 VPWR.n12 4.65
R40 VPWR.n15 VPWR.n14 4.65
R41 VPWR.n17 VPWR.n16 4.65
R42 VPWR.n19 VPWR.n18 4.65
R43 VPWR.n2 VPWR.n1 3.845
R44 VPWR.n4 VPWR.n2 0.242
R45 VPWR.n7 VPWR.n4 0.119
R46 VPWR.n9 VPWR.n7 0.119
R47 VPWR.n11 VPWR.n9 0.119
R48 VPWR.n13 VPWR.n11 0.119
R49 VPWR.n15 VPWR.n13 0.119
R50 VPWR.n17 VPWR.n15 0.119
R51 VPWR.n19 VPWR.n17 0.119
R52 VPWR VPWR.n19 0.022
R53 X.n5 X.n3 155.184
R54 X.n2 X.n0 145.662
R55 X.n5 X.n4 110.76
R56 X.n6 X.n5 56.736
R57 X.n2 X.n1 52.624
R58 X.n3 X.t2 26.595
R59 X.n3 X.t1 26.595
R60 X.n4 X.t0 26.595
R61 X.n4 X.t3 26.595
R62 X.n0 X.t6 24.923
R63 X.n0 X.t5 24.923
R64 X.n1 X.t7 24.923
R65 X.n1 X.t4 24.923
R66 X.n6 X.n2 14.222
R67 X X.n6 2.666
R68 VPB.t5 VPB.t4 556.386
R69 VPB.t6 VPB.t1 313.707
R70 VPB.t4 VPB.t8 313.707
R71 VPB.t3 VPB.t0 248.598
R72 VPB.t2 VPB.t3 248.598
R73 VPB.t1 VPB.t2 248.598
R74 VPB.t7 VPB.t6 248.598
R75 VPB.t8 VPB.t7 248.598
R76 VPB VPB.t5 192.367
R77 VGND.n0 VGND.t3 195.626
R78 VGND.n21 VGND.t5 163.563
R79 VGND.n17 VGND.t4 139.243
R80 VGND.n2 VGND.n1 115.464
R81 VGND.n13 VGND.n12 108.015
R82 VGND.n8 VGND.n7 105.973
R83 VGND.n7 VGND.t6 43.384
R84 VGND.n7 VGND.t1 26.769
R85 VGND.n1 VGND.t0 24.923
R86 VGND.n1 VGND.t2 24.923
R87 VGND.n12 VGND.t7 24.923
R88 VGND.n12 VGND.t8 24.923
R89 VGND.n22 VGND.n21 4.65
R90 VGND.n4 VGND.n3 4.65
R91 VGND.n6 VGND.n5 4.65
R92 VGND.n9 VGND.n8 4.65
R93 VGND.n11 VGND.n10 4.65
R94 VGND.n14 VGND.n13 4.65
R95 VGND.n16 VGND.n15 4.65
R96 VGND.n18 VGND.n17 4.65
R97 VGND.n20 VGND.n19 4.65
R98 VGND.n3 VGND.n2 2.258
R99 VGND.n4 VGND.n0 1.02
R100 VGND.n6 VGND.n4 0.119
R101 VGND.n9 VGND.n6 0.119
R102 VGND.n11 VGND.n9 0.119
R103 VGND.n14 VGND.n11 0.119
R104 VGND.n16 VGND.n14 0.119
R105 VGND.n18 VGND.n16 0.119
R106 VGND.n20 VGND.n18 0.119
R107 VGND.n22 VGND.n20 0.119
R108 VGND VGND.n22 0.022
R109 VNB VNB.t5 6078.09
R110 VNB.t5 VNB.t4 4545.05
R111 VNB.t6 VNB.t1 2562.64
R112 VNB.t4 VNB.t8 2562.64
R113 VNB.t0 VNB.t3 2030.77
R114 VNB.t2 VNB.t0 2030.77
R115 VNB.t1 VNB.t2 2030.77
R116 VNB.t7 VNB.t6 2030.77
R117 VNB.t8 VNB.t7 2030.77
R118 D_N.n0 D_N.t1 328.657
R119 D_N.n0 D_N.t0 126.217
R120 D_N.n1 D_N.n0 76
R121  D_N.n1 10.729
R122 D_N.n1 D_N 2.07
R123 a_109_93.n1 a_109_93.t1 425.685
R124 a_109_93.n0 a_109_93.t3 228.309
R125 a_109_93.n0 a_109_93.t2 156.009
R126 a_109_93.n2 a_109_93.n1 110.391
R127 a_109_93.n1 a_109_93.n0 92.678
R128 a_109_93.n2 a_109_93.t0 30
R129 C.n0 C.t1 241.534
R130 C.n0 C.t0 169.234
R131 C C.n0 116.501
R132 A.n0 A.t1 241.534
R133 A.n0 A.t0 169.234
R134 A A.n0 102.352
R135 B.n0 B.t1 241.534
R136 B.n0 B.t0 169.234
R137 B B.n0 109.816
R138 a_487_297.t0 a_487_297.t1 53.19
R139 a_403_297.t0 a_403_297.t1 53.19
R140 a_297_297.t0 a_297_297.t1 74.86
C0 VPWR VGND 0.12fF
C1 X VGND 0.40fF
C2 B A 0.13fF
C3 VPWR X 0.66fF
C4 B VPWR 0.10fF
C5 VPB VPWR 0.11fF
C6 C B 0.25fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__or4bb_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__or4bb_1 A X B D_N C_N VPWR VGND VNB VPB
X0 VGND.t0 A.t0 a_311_413.t0 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1 VPWR.t0 A.t1 a_561_297.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 a_393_413.t1 a_205_93.t2 a_311_413.t1 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3 VGND.t2 C_N.t0 a_27_410.t1 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 VPWR.t1 C_N.t1 a_27_410.t0 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 X.t0 a_311_413.t5 VPWR.t2 VPB.t5 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 VGND.t3 a_27_410.t2 a_311_413.t3 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7 a_561_297.t1 B.t0 a_489_297.t1 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 a_205_93.t0 D_N.t0 VGND.t6 VNB.t6 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9 a_205_93.t1 D_N.t1 VPWR.t3 VPB.t6 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10 a_489_297.t0 a_27_410.t3 a_393_413.t0 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11 a_311_413.t4 B.t1 VGND.t4 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12 a_311_413.t2 a_205_93.t3 VGND.t1 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13 X.t1 a_311_413.t6 VGND.t5 VNB.t5 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
R0 A.n0 A.t0 206.188
R1 A.n0 A.t1 148.348
R2 A A.n0 85.503
R3 a_311_413.n1 a_311_413.t1 543.076
R4 a_311_413.n0 a_311_413.t5 241.534
R5 a_311_413.n3 a_311_413.n2 170.805
R6 a_311_413.n0 a_311_413.t6 169.234
R7 a_311_413.n4 a_311_413.n3 106.429
R8 a_311_413.n1 a_311_413.n0 76
R9 a_311_413.n3 a_311_413.n1 63.397
R10 a_311_413.n2 a_311_413.t3 42.857
R11 a_311_413.n2 a_311_413.t2 38.571
R12 a_311_413.t0 a_311_413.n4 38.571
R13 a_311_413.n4 a_311_413.t4 38.571
R14 VGND.n6 VGND.t1 144.724
R15 VGND.n11 VGND.n10 135.794
R16 VGND.n3 VGND.n0 109.388
R17 VGND.n2 VGND.n1 108.015
R18 VGND.n0 VGND.t0 52.857
R19 VGND.n10 VGND.t2 45.714
R20 VGND.n1 VGND.t4 38.571
R21 VGND.n1 VGND.t3 38.571
R22 VGND.n10 VGND.t6 38.571
R23 VGND.n0 VGND.t5 30.637
R24 VGND.n12 VGND.n11 7.911
R25 VGND.n5 VGND.n4 4.65
R26 VGND.n7 VGND.n6 4.65
R27 VGND.n9 VGND.n8 4.65
R28 VGND.n3 VGND.n2 3.805
R29 VGND.n5 VGND.n3 0.254
R30 VGND.n12 VGND.n9 0.132
R31 VGND VGND.n12 0.129
R32 VGND.n7 VGND.n5 0.119
R33 VGND.n9 VGND.n7 0.119
R34 VNB VNB.t2 12650
R35 VNB.t6 VNB.t1 6115.42
R36 VNB.t2 VNB.t6 2879.41
R37 VNB.t1 VNB.t3 2814.71
R38 VNB.t4 VNB.t0 2717.65
R39 VNB.t3 VNB.t4 2717.65
R40 VNB.t0 VNB.t5 2327.87
R41 a_561_297.t0 a_561_297.t1 133.678
R42 VPWR.n1 VPWR.t3 327.591
R43 VPWR.n2 VPWR.n1 312.596
R44 VPWR.n2 VPWR.n0 173.297
R45 VPWR.n0 VPWR.t0 96.154
R46 VPWR.n1 VPWR.t1 63.321
R47 VPWR.n0 VPWR.t2 26.595
R48 VPWR VPWR.n2 0.143
R49 VPB.t6 VPB.t1 553.426
R50 VPB.t0 VPB.t5 290.031
R51 VPB.t2 VPB.t6 287.071
R52 VPB.t1 VPB.t3 284.112
R53 VPB.t4 VPB.t0 257.476
R54 VPB.t3 VPB.t4 213.084
R55 VPB VPB.t2 192.367
R56 a_205_93.n1 a_205_93.t1 403.933
R57 a_205_93.n0 a_205_93.t2 322.745
R58 a_205_93.n0 a_205_93.t3 194.212
R59 a_205_93.t0 a_205_93.n1 177.301
R60 a_205_93.n1 a_205_93.n0 76
R61 a_393_413.t0 a_393_413.t1 499.581
R62 C_N.n0 C_N.t1 329.901
R63 C_N.n0 C_N.t0 132.281
R64 C_N.n1 C_N.n0 76
R65  C_N.n1 10.422
R66 C_N.n1 C_N 2.011
R67 a_27_410.t0 a_27_410.n1 372.559
R68 a_27_410.n1 a_27_410.n0 264.234
R69 a_27_410.n1 a_27_410.t1 220.264
R70 a_27_410.n0 a_27_410.t2 206.188
R71 a_27_410.n0 a_27_410.t3 148.348
R72 X X.t0 212.866
R73 X X.t1 194.174
R74 B.t0 B.t1 397.284
R75 B B.t0 262.191
R76 a_489_297.t0 a_489_297.t1 98.5
R77 D_N.n0 D_N.t1 142.993
R78 D_N.n0 D_N.t0 126.926
R79 D_N D_N.n0 78.427
C0 VPWR X 0.13fF
C1 VPWR B 0.16fF
C2 C_N D_N 0.11fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__or4bb_2.ext - technology: sky130A

.subckt sky130_fd_sc_hd__or4bb_2 A X B D_N C_N VPWR VGND VNB VPB
X0 a_398_413.t1 a_206_93.t2 a_316_413.t4 VPB.t7 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1 VPWR.t2 a_316_413.t5 X.t3 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 X.t1 a_316_413.t6 VGND.t3 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 X.t2 a_316_413.t7 VPWR.t1 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 VGND.t5 C_N.t0 a_27_410.t1 VNB.t5 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 VPWR.t4 C_N.t1 a_27_410.t0 VPB.t5 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 VGND.t0 a_27_410.t2 a_316_413.t0 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7 VGND.t4 A.t0 a_316_413.t1 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 VGND.t2 a_316_413.t8 X.t0 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 a_566_297.t1 B.t0 a_494_297.t0 VPB.t6 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10 a_206_93.t1 D_N.t0 VGND.t1 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11 a_316_413.t2 B.t1 VGND.t6 VNB.t6 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12 a_206_93.t0 D_N.t1 VPWR.t0 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13 a_494_297.t1 a_27_410.t3 a_398_413.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14 a_316_413.t3 a_206_93.t3 VGND.t7 VNB.t7 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15 VPWR.t3 A.t1 a_566_297.t0 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
R0 a_206_93.t0 a_206_93.n1 404.583
R1 a_206_93.n0 a_206_93.t2 322.745
R2 a_206_93.n0 a_206_93.t3 194.212
R3 a_206_93.n1 a_206_93.t1 177.812
R4 a_206_93.n1 a_206_93.n0 81.27
R5 a_316_413.n3 a_316_413.t4 543.076
R6 a_316_413.n1 a_316_413.t5 212.079
R7 a_316_413.n2 a_316_413.t7 212.079
R8 a_316_413.n5 a_316_413.n4 171.934
R9 a_316_413.n1 a_316_413.t8 139.779
R10 a_316_413.n2 a_316_413.t6 139.779
R11 a_316_413.n4 a_316_413.n0 106.429
R12 a_316_413.n3 a_316_413.n2 79.651
R13 a_316_413.n4 a_316_413.n3 63.397
R14 a_316_413.n2 a_316_413.n1 61.345
R15 a_316_413.t0 a_316_413.n5 47.142
R16 a_316_413.n5 a_316_413.t3 40
R17 a_316_413.n0 a_316_413.t1 38.571
R18 a_316_413.n0 a_316_413.t2 38.571
R19 a_398_413.t0 a_398_413.t1 499.581
R20 VPB.t1 VPB.t7 568.224
R21 VPB.t4 VPB.t2 290.031
R22 VPB.t5 VPB.t1 287.071
R23 VPB.t7 VPB.t0 284.112
R24 VPB.t6 VPB.t4 257.476
R25 VPB.t2 VPB.t3 248.598
R26 VPB.t0 VPB.t6 213.084
R27 VPB VPB.t5 189.408
R28 X X.n1 169.251
R29 X X.n0 152.895
R30 X.n0 X.t3 26.595
R31 X.n0 X.t2 26.595
R32 X.n1 X.t0 24.923
R33 X.n1 X.t1 24.923
R34 VPWR.n13 VPWR.t0 327.591
R35 VPWR.n14 VPWR.n13 309.178
R36 VPWR.n2 VPWR.t2 170.512
R37 VPWR.n1 VPWR.n0 169.105
R38 VPWR.n0 VPWR.t3 96.154
R39 VPWR.n13 VPWR.t4 63.321
R40 VPWR.n0 VPWR.t1 26.595
R41 VPWR.n4 VPWR.n3 4.65
R42 VPWR.n6 VPWR.n5 4.65
R43 VPWR.n8 VPWR.n7 4.65
R44 VPWR.n10 VPWR.n9 4.65
R45 VPWR.n12 VPWR.n11 4.65
R46 VPWR.n15 VPWR.n14 3.932
R47 VPWR.n2 VPWR.n1 3.86
R48 VPWR.n4 VPWR.n2 0.248
R49 VPWR.n15 VPWR.n12 0.137
R50 VPWR VPWR.n15 0.121
R51 VPWR.n6 VPWR.n4 0.119
R52 VPWR.n8 VPWR.n6 0.119
R53 VPWR.n10 VPWR.n8 0.119
R54 VPWR.n12 VPWR.n10 0.119
R55 VGND.n10 VGND.t7 145.493
R56 VGND.n15 VGND.n14 135.794
R57 VGND.n2 VGND.t2 117.062
R58 VGND.n6 VGND.n5 108.015
R59 VGND.n1 VGND.n0 105.973
R60 VGND.n0 VGND.t4 52.857
R61 VGND.n14 VGND.t5 45.714
R62 VGND.n5 VGND.t6 38.571
R63 VGND.n5 VGND.t0 38.571
R64 VGND.n14 VGND.t1 38.571
R65 VGND.n0 VGND.t3 30.637
R66 VGND.n16 VGND.n15 8.288
R67 VGND.n4 VGND.n3 4.65
R68 VGND.n7 VGND.n6 4.65
R69 VGND.n9 VGND.n8 4.65
R70 VGND.n11 VGND.n10 4.65
R71 VGND.n13 VGND.n12 4.65
R72 VGND.n2 VGND.n1 3.822
R73 VGND.n4 VGND.n2 0.254
R74 VGND.n16 VGND.n13 0.132
R75 VGND VGND.n16 0.127
R76 VGND.n7 VGND.n4 0.119
R77 VGND.n9 VGND.n7 0.119
R78 VGND.n11 VGND.n9 0.119
R79 VGND.n13 VGND.n11 0.119
R80 VNB VNB.t5 12650
R81 VNB.t1 VNB.t7 6115.42
R82 VNB.t7 VNB.t0 2944.12
R83 VNB.t5 VNB.t1 2879.41
R84 VNB.t6 VNB.t4 2717.65
R85 VNB.t0 VNB.t6 2717.65
R86 VNB.t4 VNB.t3 2327.87
R87 VNB.t3 VNB.t2 2030.77
R88 C_N.n0 C_N.t1 329.901
R89 C_N.n0 C_N.t0 132.281
R90 C_N.n1 C_N.n0 76
R91  C_N.n1 10.422
R92 C_N.n1 C_N 2.011
R93 a_27_410.t0 a_27_410.n1 372.559
R94 a_27_410.n1 a_27_410.n0 266.117
R95 a_27_410.n1 a_27_410.t1 217.923
R96 a_27_410.n0 a_27_410.t2 206.188
R97 a_27_410.n0 a_27_410.t3 148.348
R98 A.n0 A.t0 206.188
R99 A.n0 A.t1 148.348
R100 A A.n0 85.503
R101 B.t0 B.t1 397.284
R102 B B.t0 262.191
R103 a_494_297.t0 a_494_297.t1 98.5
R104 a_566_297.t0 a_566_297.t1 133.678
R105 D_N.n0 D_N.t1 142.993
R106 D_N.n0 D_N.t0 126.926
R107 D_N D_N.n0 78.427
C0 VPWR X 0.24fF
C1 C_N D_N 0.11fF
C2 VPWR B 0.16fF
C3 VPB VPWR 0.10fF
C4 VPWR VGND 0.12fF
C5 X VGND 0.12fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__or4bb_4.ext - technology: sky130A

.subckt sky130_fd_sc_hd__or4bb_4 D_N B A C_N X VGND VPWR VNB VPB
X0 VPWR.t6 a_315_380.t5 X.t7 VPB.t9 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 X.t6 a_315_380.t6 VPWR.t5 VPB.t8 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 a_315_380.t1 B.t0 VGND.t9 VNB.t9 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 VGND.t0 C_N.t0 a_27_410.t0 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 VPWR.t0 C_N.t1 a_27_410.t1 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 VPWR.t1 A.t0 a_583_297.t0 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 VGND.t1 a_27_410.t2 a_315_380.t0 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 a_583_297.t1 B.t1 a_499_297.t1 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 VGND.t2 A.t1 a_315_380.t2 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 a_397_297.t1 a_205_93.t2 a_315_380.t3 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 X.t3 a_315_380.t7 VGND.t8 VNB.t8 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 X.t2 a_315_380.t8 VGND.t7 VNB.t7 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 a_499_297.t0 a_27_410.t3 a_397_297.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13 VPWR.t4 a_315_380.t9 X.t5 VPB.t7 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14 a_205_93.t0 D_N.t0 VGND.t4 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15 a_205_93.t1 D_N.t1 VPWR.t2 VPB.t5 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16 VGND.t6 a_315_380.t10 X.t1 VNB.t6 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X17 VGND.t5 a_315_380.t11 X.t0 VNB.t5 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X18 a_315_380.t4 a_205_93.t3 VGND.t3 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X19 X.t4 a_315_380.t12 VPWR.t3 VPB.t6 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
R0 a_315_380.n15 a_315_380.n14 415.406
R1 a_315_380.n2 a_315_380.t9 212.079
R2 a_315_380.n4 a_315_380.t12 212.079
R3 a_315_380.n7 a_315_380.t5 212.079
R4 a_315_380.n10 a_315_380.t6 212.079
R5 a_315_380.n16 a_315_380.n15 162.235
R6 a_315_380.n2 a_315_380.t11 139.779
R7 a_315_380.n4 a_315_380.t8 139.779
R8 a_315_380.n7 a_315_380.t10 139.779
R9 a_315_380.n10 a_315_380.t7 139.779
R10 a_315_380.n14 a_315_380.n0 104.923
R11 a_315_380.n13 a_315_380.n1 104.923
R12 a_315_380.n6 a_315_380.n3 101.6
R13 a_315_380.n13 a_315_380.n12 79.057
R14 a_315_380.n6 a_315_380.n5 76
R15 a_315_380.n9 a_315_380.n8 76
R16 a_315_380.n12 a_315_380.n11 76
R17 a_315_380.n14 a_315_380.n13 65.505
R18 a_315_380.n0 a_315_380.t4 39.692
R19 a_315_380.n0 a_315_380.t0 30.461
R20 a_315_380.n3 a_315_380.n2 26.29
R21 a_315_380.n15 a_315_380.t3 26.266
R22 a_315_380.n9 a_315_380.n6 25.6
R23 a_315_380.n12 a_315_380.n9 25.6
R24 a_315_380.n1 a_315_380.t2 24.923
R25 a_315_380.n1 a_315_380.t1 24.923
R26 a_315_380.n5 a_315_380.n4 14.606
R27 a_315_380.n11 a_315_380.n10 8.763
R28 a_315_380.n8 a_315_380.n7 2.921
R29 X.n5 X.n3 155.184
R30 X.n2 X.n0 145.662
R31 X.n5 X.n4 110.76
R32 X.n6 X.n5 58.417
R33 X.n2 X.n1 52.624
R34 X.n3 X.t7 26.595
R35 X.n3 X.t6 26.595
R36 X.n4 X.t5 26.595
R37 X.n4 X.t4 26.595
R38 X.n0 X.t1 24.923
R39 X.n0 X.t3 24.923
R40 X.n1 X.t0 24.923
R41 X.n1 X.t2 24.923
R42 X.n6 X.n2 14.222
R43 X X.n6 2.782
R44 VPWR.n18 VPWR.t2 327.591
R45 VPWR.n19 VPWR.n18 309.178
R46 VPWR.n2 VPWR.t4 202.619
R47 VPWR.n1 VPWR.n0 171.981
R48 VPWR.n6 VPWR.n5 171.981
R49 VPWR.n18 VPWR.t0 63.321
R50 VPWR.n5 VPWR.t5 37.43
R51 VPWR.n5 VPWR.t1 37.43
R52 VPWR.n0 VPWR.t3 26.595
R53 VPWR.n0 VPWR.t6 26.595
R54 VPWR.n4 VPWR.n3 4.65
R55 VPWR.n7 VPWR.n6 4.65
R56 VPWR.n9 VPWR.n8 4.65
R57 VPWR.n11 VPWR.n10 4.65
R58 VPWR.n13 VPWR.n12 4.65
R59 VPWR.n15 VPWR.n14 4.65
R60 VPWR.n17 VPWR.n16 4.65
R61 VPWR.n20 VPWR.n19 3.932
R62 VPWR.n2 VPWR.n1 3.811
R63 VPWR.n4 VPWR.n2 0.243
R64 VPWR.n20 VPWR.n17 0.137
R65 VPWR VPWR.n20 0.123
R66 VPWR.n7 VPWR.n4 0.119
R67 VPWR.n9 VPWR.n7 0.119
R68 VPWR.n11 VPWR.n9 0.119
R69 VPWR.n13 VPWR.n11 0.119
R70 VPWR.n15 VPWR.n13 0.119
R71 VPWR.n17 VPWR.n15 0.119
R72 VPB.t5 VPB.t4 565.264
R73 VPB.t3 VPB.t8 313.707
R74 VPB.t4 VPB.t0 301.869
R75 VPB.t1 VPB.t5 287.071
R76 VPB.t6 VPB.t7 248.598
R77 VPB.t9 VPB.t6 248.598
R78 VPB.t8 VPB.t9 248.598
R79 VPB.t2 VPB.t3 248.598
R80 VPB.t0 VPB.t2 248.598
R81 VPB VPB.t1 192.367
R82 B.n0 B.t1 241.534
R83 B.n0 B.t0 169.234
R84 B B.n0 107.667
R85 VGND.n0 VGND.t5 199.091
R86 VGND.n17 VGND.t3 183.974
R87 VGND.n22 VGND.n21 135.794
R88 VGND.n2 VGND.n1 115.464
R89 VGND.n13 VGND.n12 108.015
R90 VGND.n8 VGND.n7 105.973
R91 VGND.n21 VGND.t0 45.714
R92 VGND.n7 VGND.t2 43.384
R93 VGND.n21 VGND.t4 38.571
R94 VGND.n7 VGND.t8 26.769
R95 VGND.n1 VGND.t7 24.923
R96 VGND.n1 VGND.t6 24.923
R97 VGND.n12 VGND.t9 24.923
R98 VGND.n12 VGND.t1 24.923
R99 VGND.n23 VGND.n22 7.911
R100 VGND.n4 VGND.n3 4.65
R101 VGND.n6 VGND.n5 4.65
R102 VGND.n9 VGND.n8 4.65
R103 VGND.n11 VGND.n10 4.65
R104 VGND.n14 VGND.n13 4.65
R105 VGND.n16 VGND.n15 4.65
R106 VGND.n18 VGND.n17 4.65
R107 VGND.n20 VGND.n19 4.65
R108 VGND.n3 VGND.n2 3.764
R109 VGND.n4 VGND.n0 0.861
R110 VGND.n23 VGND.n20 0.132
R111 VGND VGND.n23 0.129
R112 VGND.n6 VGND.n4 0.119
R113 VGND.n9 VGND.n6 0.119
R114 VGND.n11 VGND.n9 0.119
R115 VGND.n14 VGND.n11 0.119
R116 VGND.n16 VGND.n14 0.119
R117 VGND.n18 VGND.n16 0.119
R118 VGND.n20 VGND.n18 0.119
R119 VNB VNB.t0 12650
R120 VNB.t4 VNB.t3 5321.88
R121 VNB.t0 VNB.t4 2879.41
R122 VNB.t2 VNB.t8 2562.64
R123 VNB.t3 VNB.t1 2562.64
R124 VNB.t7 VNB.t5 2030.77
R125 VNB.t6 VNB.t7 2030.77
R126 VNB.t8 VNB.t6 2030.77
R127 VNB.t9 VNB.t2 2030.77
R128 VNB.t1 VNB.t9 2030.77
R129 C_N.n0 C_N.t1 329.901
R130 C_N.n0 C_N.t0 132.281
R131 C_N.n1 C_N.n0 76
R132  C_N.n1 10.422
R133 C_N.n1 C_N 2.011
R134 a_27_410.n1 a_27_410.t1 372.559
R135 a_27_410.n1 a_27_410.n0 332.751
R136 a_27_410.n0 a_27_410.t3 241.534
R137 a_27_410.t0 a_27_410.n1 220.264
R138 a_27_410.n0 a_27_410.t2 169.234
R139 A.n0 A.t0 241.534
R140 A.n0 A.t1 169.234
R141 A A.n0 102.352
R142 a_583_297.t0 a_583_297.t1 53.19
R143 a_499_297.t0 a_499_297.t1 53.19
R144 a_205_93.n1 a_205_93.t1 403.116
R145 a_205_93.n0 a_205_93.t2 227.673
R146 a_205_93.t0 a_205_93.n1 173.978
R147 a_205_93.n0 a_205_93.t3 155.373
R148 a_205_93.n1 a_205_93.n0 76
R149 a_397_297.t0 a_397_297.t1 70.92
R150 D_N.n0 D_N.t1 142.993
R151 D_N.n0 D_N.t0 126.926
R152 D_N D_N.n0 78.427
C0 B A 0.13fF
C1 B VPWR 0.10fF
C2 C_N D_N 0.11fF
C3 X VGND 0.40fF
C4 VPWR X 0.65fF
C5 VPB VPWR 0.11fF
C6 VPWR VGND 0.12fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__probe_p_8.ext - technology: sky130A

.subckt sky130_fd_sc_hd__probe_p_8 X A VGND VPWR VNB VPB
X0 a_361_47.t7 a_27_47.t6 VGND.t10 VNB.t10 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 a_361_47.t6 a_27_47.t7 VGND.t9 VNB.t9 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 a_361_47.t5 a_27_47.t8 VGND.t8 VNB.t8 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 VPWR.t10 a_27_47.t9 a_361_47.t15 VPB.t10 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 a_361_47.t14 a_27_47.t10 VPWR.t9 VPB.t9 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 VGND.t7 a_27_47.t11 a_361_47.t4 VNB.t7 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 VPWR.t1 A.t0 a_27_47.t2 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 VPWR.t8 a_27_47.t12 a_361_47.t13 VPB.t8 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 a_27_47.t0 A.t1 VPWR.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 a_361_47.t12 a_27_47.t13 VPWR.t7 VPB.t7 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 a_27_47.t1 A.t2 VGND.t0 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 a_361_47.t3 a_27_47.t14 VGND.t6 VNB.t6 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 VPWR.t6 a_27_47.t15 a_361_47.t11 VPB.t6 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13 a_361_47.t10 a_27_47.t16 VPWR.t5 VPB.t5 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14 VGND.t1 A.t3 a_27_47.t3 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X15 VGND.t5 a_27_47.t17 a_361_47.t2 VNB.t5 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X16 VPWR.t4 a_27_47.t18 a_361_47.t9 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17 VGND.t4 a_27_47.t19 a_361_47.t1 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X18 VGND.t3 a_27_47.t20 a_361_47.t0 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X19 a_361_47.t8 a_27_47.t21 VPWR.t3 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X20 VPWR.t2 A.t4 a_27_47.t4 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X21 VGND.t2 A.t5 a_27_47.t5 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
R0 a_27_47.n0 a_27_47.t12 221.719
R1 a_27_47.n1 a_27_47.t13 221.719
R2 a_27_47.n2 a_27_47.t15 221.719
R3 a_27_47.n6 a_27_47.t16 221.719
R4 a_27_47.n9 a_27_47.t18 221.719
R5 a_27_47.n12 a_27_47.t21 221.719
R6 a_27_47.n15 a_27_47.t9 221.719
R7 a_27_47.n18 a_27_47.t10 221.719
R8 a_27_47.n22 a_27_47.t5 193.846
R9 a_27_47.n24 a_27_47.t4 173.405
R10 a_27_47.n0 a_27_47.t11 149.419
R11 a_27_47.n1 a_27_47.t8 149.419
R12 a_27_47.n2 a_27_47.t20 149.419
R13 a_27_47.n6 a_27_47.t7 149.419
R14 a_27_47.n9 a_27_47.t19 149.419
R15 a_27_47.n12 a_27_47.t6 149.419
R16 a_27_47.n15 a_27_47.t17 149.419
R17 a_27_47.n18 a_27_47.t14 149.419
R18 a_27_47.n25 a_27_47.n24 108.41
R19 a_27_47.n22 a_27_47.n21 105.676
R20 a_27_47.n5 a_27_47.n3 101.6
R21 a_27_47.n5 a_27_47.n4 76
R22 a_27_47.n8 a_27_47.n7 76
R23 a_27_47.n11 a_27_47.n10 76
R24 a_27_47.n14 a_27_47.n13 76
R25 a_27_47.n17 a_27_47.n16 76
R26 a_27_47.n20 a_27_47.n19 76
R27 a_27_47.n1 a_27_47.n0 74.977
R28 a_27_47.n3 a_27_47.n1 66.051
R29 a_27_47.n23 a_27_47.n22 48.962
R30 a_27_47.n24 a_27_47.n23 38.732
R31 a_27_47.n7 a_27_47.n6 37.488
R32 a_27_47.n25 a_27_47.t2 26.595
R33 a_27_47.t0 a_27_47.n25 26.595
R34 a_27_47.n8 a_27_47.n5 25.6
R35 a_27_47.n11 a_27_47.n8 25.6
R36 a_27_47.n14 a_27_47.n11 25.6
R37 a_27_47.n17 a_27_47.n14 25.6
R38 a_27_47.n20 a_27_47.n17 25.6
R39 a_27_47.n21 a_27_47.t3 24.923
R40 a_27_47.n21 a_27_47.t1 24.923
R41 a_27_47.n10 a_27_47.n9 23.207
R42 a_27_47.n19 a_27_47.n18 19.637
R43 a_27_47.n23 a_27_47.n20 18.447
R44 a_27_47.n3 a_27_47.n2 8.925
R45 a_27_47.n13 a_27_47.n12 8.925
R46 a_27_47.n16 a_27_47.n15 5.355
R47 VGND.n1 VGND.n0 108.015
R48 VGND.n6 VGND.n5 108.015
R49 VGND.n10 VGND.n9 108.015
R50 VGND.n16 VGND.n15 108.015
R51 VGND.n21 VGND.n20 108.015
R52 VGND.n2 VGND.t7 106.996
R53 VGND.n0 VGND.t8 24.923
R54 VGND.n0 VGND.t3 24.923
R55 VGND.n5 VGND.t9 24.923
R56 VGND.n5 VGND.t4 24.923
R57 VGND.n9 VGND.t10 24.923
R58 VGND.n9 VGND.t5 24.923
R59 VGND.n15 VGND.t6 24.923
R60 VGND.n15 VGND.t1 24.923
R61 VGND.n20 VGND.t0 24.923
R62 VGND.n20 VGND.t2 24.923
R63 VGND.n4 VGND.n3 4.65
R64 VGND.n8 VGND.n7 4.65
R65 VGND.n12 VGND.n11 4.65
R66 VGND.n14 VGND.n13 4.65
R67 VGND.n17 VGND.n16 4.65
R68 VGND.n19 VGND.n18 4.65
R69 VGND.n22 VGND.n21 3.932
R70 VGND.n2 VGND.n1 3.488
R71 VGND.n7 VGND.n6 3.388
R72 VGND.n11 VGND.n10 0.376
R73 VGND.n4 VGND.n2 0.263
R74 VGND.n22 VGND.n19 0.137
R75 VGND VGND.n22 0.121
R76 VGND.n8 VGND.n4 0.119
R77 VGND.n12 VGND.n8 0.119
R78 VGND.n14 VGND.n12 0.119
R79 VGND.n17 VGND.n14 0.119
R80 VGND.n19 VGND.n17 0.119
R81 a_361_47.n5 a_361_47.n4 228.465
R82 a_361_47.n8 a_361_47.n7 169.484
R83 a_361_47.n14 a_361_47.n13 168.923
R84 a_361_47.n6 a_361_47.n2 165.218
R85 a_361_47.n5 a_361_47.n3 165.218
R86 a_361_47.n11 a_361_47.n10 109.942
R87 a_361_47.n12 a_361_47.n1 105.676
R88 a_361_47.n15 a_361_47.n14 105.676
R89 a_361_47.n6 a_361_47.n5 63.247
R90 a_361_47.n14 a_361_47.n12 63.247
R91 a_361_47.n8 a_361_47.n6 50.447
R92 a_361_47.n12 a_361_47.n11 50.447
R93 a_361_47.n2 a_361_47.t11 26.595
R94 a_361_47.n2 a_361_47.t10 26.595
R95 a_361_47.n3 a_361_47.t9 26.595
R96 a_361_47.n3 a_361_47.t8 26.595
R97 a_361_47.n4 a_361_47.t15 26.595
R98 a_361_47.n4 a_361_47.t14 26.595
R99 a_361_47.n7 a_361_47.t13 26.595
R100 a_361_47.n7 a_361_47.t12 26.595
R101 a_361_47.n10 a_361_47.t4 24.923
R102 a_361_47.n10 a_361_47.t5 24.923
R103 a_361_47.n13 a_361_47.t2 24.923
R104 a_361_47.n13 a_361_47.t3 24.923
R105 a_361_47.n1 a_361_47.t0 24.923
R106 a_361_47.n1 a_361_47.t6 24.923
R107 a_361_47.n15 a_361_47.t1 24.923
R108 a_361_47.t7 a_361_47.n15 24.923
R109 a_361_47.n11 a_361_47.n9 11.796
R110 a_361_47.n9 a_361_47.n8 10.792
R111 a_361_47.n9 a_361_47.n0 6.376
R112 VNB VNB.t2 6053.91
R113 VNB.t8 VNB.t7 2030.77
R114 VNB.t3 VNB.t8 2030.77
R115 VNB.t9 VNB.t3 2030.77
R116 VNB.t4 VNB.t9 2030.77
R117 VNB.t10 VNB.t4 2030.77
R118 VNB.t5 VNB.t10 2030.77
R119 VNB.t6 VNB.t5 2030.77
R120 VNB.t1 VNB.t6 2030.77
R121 VNB.t0 VNB.t1 2030.77
R122 VNB.t2 VNB.t0 2030.77
R123 VPWR.n22 VPWR.n21 174.594
R124 VPWR.n16 VPWR.n15 174.594
R125 VPWR.n1 VPWR.n0 164.214
R126 VPWR.n6 VPWR.n5 164.214
R127 VPWR.n10 VPWR.n9 164.214
R128 VPWR.n2 VPWR.t8 149.356
R129 VPWR.n0 VPWR.t7 26.595
R130 VPWR.n0 VPWR.t6 26.595
R131 VPWR.n5 VPWR.t5 26.595
R132 VPWR.n5 VPWR.t4 26.595
R133 VPWR.n9 VPWR.t3 26.595
R134 VPWR.n9 VPWR.t10 26.595
R135 VPWR.n21 VPWR.t0 26.595
R136 VPWR.n21 VPWR.t2 26.595
R137 VPWR.n15 VPWR.t9 26.595
R138 VPWR.n15 VPWR.t1 26.595
R139 VPWR.n17 VPWR.n16 6.776
R140 VPWR.n24 VPWR.n23 4.65
R141 VPWR.n4 VPWR.n3 4.65
R142 VPWR.n8 VPWR.n7 4.65
R143 VPWR.n12 VPWR.n11 4.65
R144 VPWR.n14 VPWR.n13 4.65
R145 VPWR.n18 VPWR.n17 4.65
R146 VPWR.n20 VPWR.n19 4.65
R147 VPWR.n2 VPWR.n1 3.488
R148 VPWR.n7 VPWR.n6 3.388
R149 VPWR.n23 VPWR.n22 0.752
R150 VPWR.n11 VPWR.n10 0.376
R151 VPWR.n4 VPWR.n2 0.263
R152 VPWR.n8 VPWR.n4 0.119
R153 VPWR.n12 VPWR.n8 0.119
R154 VPWR.n14 VPWR.n12 0.119
R155 VPWR.n18 VPWR.n14 0.119
R156 VPWR.n20 VPWR.n18 0.119
R157 VPWR.n24 VPWR.n20 0.119
R158 VPWR.n25 VPWR.n24 0.119
R159 VPWR VPWR.n25 0.02
R160 VPB.t7 VPB.t8 248.598
R161 VPB.t6 VPB.t7 248.598
R162 VPB.t5 VPB.t6 248.598
R163 VPB.t4 VPB.t5 248.598
R164 VPB.t3 VPB.t4 248.598
R165 VPB.t10 VPB.t3 248.598
R166 VPB.t9 VPB.t10 248.598
R167 VPB.t1 VPB.t9 248.598
R168 VPB.t0 VPB.t1 248.598
R169 VPB.t2 VPB.t0 248.598
R170 VPB VPB.t2 189.408
R171 A.n6 A.t4 235.762
R172 A.n0 A.t0 221.719
R173 A.n2 A.t1 221.719
R174 A.n6 A.t5 163.462
R175 A.n0 A.t3 149.419
R176 A.n2 A.t2 149.419
R177 A.n5 A.n4 76
R178 A.n7 A.n6 76
R179 A.n1 A.n0 58.018
R180 A.n5 A.n2 43.737
R181 A.n4 A.n3 21.76
R182 A.n7 A 19.52
R183 A.n6 A.n5 17.851
R184 A.n2 A.n1 16.959
R185 A A.n7 9.92
R186 A.n3 A 5.44
R187 A.n4 A 2.24
C0 VPWR VGND 0.12fF
C1 VPB VPWR 0.12fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__probec_p_8.ext - technology: sky130A

.subckt sky130_fd_sc_hd__probec_p_8 X A VGND VPWR VNB VPB
X0 a_361_47.t7 a_27_47.t6 VGND.t7 VNB.t7 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
R0 VPWR m5_872_595# sky130_fd_pr__res_generic_m5 w=2.11616e+11u l=1.2e+06u
X1 a_361_47.t6 a_27_47.t7 VGND.t6 VNB.t6 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 a_361_47.t5 a_27_47.t8 VGND.t5 VNB.t5 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 VPWR.t7 a_27_47.t9 a_361_47.t15 VPB.t7 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
R1 VGND m5_872_n71# sky130_fd_pr__res_generic_m5 w=2.11616e+11u l=1.2e+06u
X4 a_361_47.t14 a_27_47.t10 VPWR.t6 VPB.t6 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 VGND.t4 a_27_47.t11 a_361_47.t4 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 VPWR.t8 A.t0 a_27_47.t0 VPB.t8 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 VPWR.t5 a_27_47.t12 a_361_47.t13 VPB.t5 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 a_27_47.t1 A.t1 VPWR.t9 VPB.t9 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 a_361_47.t12 a_27_47.t13 VPWR.t4 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 a_27_47.t2 A.t2 VGND.t8 VNB.t8 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 a_361_47.t3 a_27_47.t14 VGND.t3 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 VPWR.t3 a_27_47.t15 a_361_47.t11 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13 a_361_47.t10 a_27_47.t16 VPWR.t2 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14 VGND.t9 A.t3 a_27_47.t3 VNB.t9 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X15 VGND.t2 a_27_47.t17 a_361_47.t2 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X16 VPWR.t1 a_27_47.t18 a_361_47.t9 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17 VGND.t1 a_27_47.t19 a_361_47.t1 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X18 VGND.t0 a_27_47.t20 a_361_47.t0 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X19 a_361_47.t8 a_27_47.t21 VPWR.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X20 VPWR.t10 A.t4 a_27_47.t4 VPB.t10 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X21 VGND.t10 A.t5 a_27_47.t5 VNB.t10 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
R2 a_27_47.n0 a_27_47.t12 221.719
R3 a_27_47.n1 a_27_47.t13 221.719
R4 a_27_47.n2 a_27_47.t15 221.719
R5 a_27_47.n6 a_27_47.t16 221.719
R6 a_27_47.n9 a_27_47.t18 221.719
R7 a_27_47.n12 a_27_47.t21 221.719
R8 a_27_47.n15 a_27_47.t9 221.719
R9 a_27_47.n18 a_27_47.t10 221.719
R10 a_27_47.n22 a_27_47.t5 193.846
R11 a_27_47.n24 a_27_47.t4 173.405
R12 a_27_47.n0 a_27_47.t11 149.419
R13 a_27_47.n1 a_27_47.t8 149.419
R14 a_27_47.n2 a_27_47.t20 149.419
R15 a_27_47.n6 a_27_47.t7 149.419
R16 a_27_47.n9 a_27_47.t19 149.419
R17 a_27_47.n12 a_27_47.t6 149.419
R18 a_27_47.n15 a_27_47.t17 149.419
R19 a_27_47.n18 a_27_47.t14 149.419
R20 a_27_47.n25 a_27_47.n24 108.41
R21 a_27_47.n22 a_27_47.n21 105.676
R22 a_27_47.n5 a_27_47.n3 101.6
R23 a_27_47.n5 a_27_47.n4 76
R24 a_27_47.n8 a_27_47.n7 76
R25 a_27_47.n11 a_27_47.n10 76
R26 a_27_47.n14 a_27_47.n13 76
R27 a_27_47.n17 a_27_47.n16 76
R28 a_27_47.n20 a_27_47.n19 76
R29 a_27_47.n1 a_27_47.n0 74.977
R30 a_27_47.n3 a_27_47.n1 66.051
R31 a_27_47.n23 a_27_47.n22 48.962
R32 a_27_47.n24 a_27_47.n23 38.732
R33 a_27_47.n7 a_27_47.n6 37.488
R34 a_27_47.t0 a_27_47.n25 26.595
R35 a_27_47.n25 a_27_47.t1 26.595
R36 a_27_47.n8 a_27_47.n5 25.6
R37 a_27_47.n11 a_27_47.n8 25.6
R38 a_27_47.n14 a_27_47.n11 25.6
R39 a_27_47.n17 a_27_47.n14 25.6
R40 a_27_47.n20 a_27_47.n17 25.6
R41 a_27_47.n21 a_27_47.t3 24.923
R42 a_27_47.n21 a_27_47.t2 24.923
R43 a_27_47.n10 a_27_47.n9 23.207
R44 a_27_47.n19 a_27_47.n18 19.637
R45 a_27_47.n23 a_27_47.n20 18.447
R46 a_27_47.n3 a_27_47.n2 8.925
R47 a_27_47.n13 a_27_47.n12 8.925
R48 a_27_47.n16 a_27_47.n15 5.355
R49 VGND.n27 VGND.n26 108.015
R50 VGND.n32 VGND.n31 108.015
R51 VGND.n36 VGND.n35 108.015
R52 VGND.n42 VGND.n41 108.015
R53 VGND.n47 VGND.n46 108.015
R54 VGND.n22 VGND.t4 103.506
R55 VGND.n26 VGND.t5 24.923
R56 VGND.n26 VGND.t0 24.923
R57 VGND.n31 VGND.t6 24.923
R58 VGND.n31 VGND.t1 24.923
R59 VGND.n35 VGND.t7 24.923
R60 VGND.n35 VGND.t2 24.923
R61 VGND.n41 VGND.t3 24.923
R62 VGND.n41 VGND.t9 24.923
R63 VGND.n46 VGND.t8 24.923
R64 VGND.n46 VGND.t10 24.923
R65 VGND.n25 VGND.n24 4.65
R66 VGND.n28 VGND.n27 4.65
R67 VGND.n30 VGND.n29 4.65
R68 VGND.n34 VGND.n33 4.65
R69 VGND.n38 VGND.n37 4.65
R70 VGND.n40 VGND.n39 4.65
R71 VGND.n43 VGND.n42 4.65
R72 VGND.n45 VGND.n44 4.65
R73 VGND.n48 VGND.n47 3.932
R74 VGND.n23 VGND.n22 3.65
R75 VGND.n33 VGND.n32 3.388
R76 VGND.n16 VGND.n15 0.864
R77 VGND.n21 VGND.n20 0.521
R78 VGND.n37 VGND.n36 0.376
R79 VGND.n14 VGND.n13 0.285
R80 VGND.n25 VGND.n23 0.143
R81 VGND.n48 VGND.n45 0.137
R82 VGND VGND.n48 0.121
R83 VGND.n28 VGND.n25 0.119
R84 VGND.n30 VGND.n28 0.119
R85 VGND.n34 VGND.n30 0.119
R86 VGND.n38 VGND.n34 0.119
R87 VGND.n40 VGND.n38 0.119
R88 VGND.n43 VGND.n40 0.119
R89 VGND.n45 VGND.n43 0.119
R90 VGND.n23 VGND.n21 0.1
R91 VGND.n11 VGND.n7 0.095
R92 VGND.n20 VGND.n16 0.092
R93 VGND.n20 VGND.n19 0.061
R94 VGND.n5 VGND.n4 0.017
R95 VGND.n3 VGND.n2 0.017
R96 VGND.n1 VGND.n0 0.016
R97 VGND.n4 VGND.n3 0.014
R98 VGND.n19 VGND.n18 0.011
R99 VGND.n18 VGND.n17 0.008
R100 VGND.n13 VGND.n12 0.005
R101 VGND.n10 VGND.n9 0.005
R102 VGND.n15 VGND.n14 0.004
R103 VGND.n14 VGND.n5 0.003
R104 VGND.n2 VGND.n1 0.003
R105 VGND.n13 VGND.n6 0.003
R106 VGND.n9 VGND.n8 0.003
R107 VGND.n12 VGND.n11 0.001
R108 VGND.n11 VGND.n10 0.001
R109 a_361_47.n4 a_361_47.n3 228.465
R110 a_361_47.n7 a_361_47.n6 169.484
R111 a_361_47.n12 a_361_47.n11 168.923
R112 a_361_47.n5 a_361_47.n1 165.218
R113 a_361_47.n4 a_361_47.n2 165.218
R114 a_361_47.n9 a_361_47.n8 109.942
R115 a_361_47.n10 a_361_47.n0 105.676
R116 a_361_47.n13 a_361_47.n12 105.676
R117 a_361_47.n5 a_361_47.n4 63.247
R118 a_361_47.n12 a_361_47.n10 63.247
R119 a_361_47.n7 a_361_47.n5 50.447
R120 a_361_47.n10 a_361_47.n9 50.447
R121 a_361_47.n1 a_361_47.t11 26.595
R122 a_361_47.n1 a_361_47.t10 26.595
R123 a_361_47.n2 a_361_47.t9 26.595
R124 a_361_47.n2 a_361_47.t8 26.595
R125 a_361_47.n3 a_361_47.t15 26.595
R126 a_361_47.n3 a_361_47.t14 26.595
R127 a_361_47.n6 a_361_47.t13 26.595
R128 a_361_47.n6 a_361_47.t12 26.595
R129 a_361_47.n8 a_361_47.t4 24.923
R130 a_361_47.n8 a_361_47.t5 24.923
R131 a_361_47.n11 a_361_47.t2 24.923
R132 a_361_47.n11 a_361_47.t3 24.923
R133 a_361_47.n0 a_361_47.t0 24.923
R134 a_361_47.n0 a_361_47.t6 24.923
R135 a_361_47.n13 a_361_47.t1 24.923
R136 a_361_47.t7 a_361_47.n13 24.923
R137 a_361_47.n9 a_361_47.n7 22.588
R138 VNB VNB.t10 6053.91
R139 VNB.t5 VNB.t4 2030.77
R140 VNB.t0 VNB.t5 2030.77
R141 VNB.t6 VNB.t0 2030.77
R142 VNB.t1 VNB.t6 2030.77
R143 VNB.t7 VNB.t1 2030.77
R144 VNB.t2 VNB.t7 2030.77
R145 VNB.t3 VNB.t2 2030.77
R146 VNB.t9 VNB.t3 2030.77
R147 VNB.t8 VNB.t9 2030.77
R148 VNB.t10 VNB.t8 2030.77
R149 VPWR.n48 VPWR.n47 174.594
R150 VPWR.n42 VPWR.n41 174.594
R151 VPWR.n27 VPWR.n26 164.214
R152 VPWR.n32 VPWR.n31 164.214
R153 VPWR.n36 VPWR.n35 164.214
R154 VPWR.n22 VPWR.t5 145.866
R155 VPWR.n26 VPWR.t4 26.595
R156 VPWR.n26 VPWR.t3 26.595
R157 VPWR.n31 VPWR.t2 26.595
R158 VPWR.n31 VPWR.t1 26.595
R159 VPWR.n35 VPWR.t0 26.595
R160 VPWR.n35 VPWR.t7 26.595
R161 VPWR.n47 VPWR.t9 26.595
R162 VPWR.n47 VPWR.t10 26.595
R163 VPWR.n41 VPWR.t6 26.595
R164 VPWR.n41 VPWR.t8 26.595
R165 VPWR.n43 VPWR.n42 6.776
R166 VPWR.n50 VPWR.n49 4.65
R167 VPWR.n25 VPWR.n24 4.65
R168 VPWR.n28 VPWR.n27 4.65
R169 VPWR.n30 VPWR.n29 4.65
R170 VPWR.n34 VPWR.n33 4.65
R171 VPWR.n38 VPWR.n37 4.65
R172 VPWR.n40 VPWR.n39 4.65
R173 VPWR.n44 VPWR.n43 4.65
R174 VPWR.n46 VPWR.n45 4.65
R175 VPWR.n23 VPWR.n22 3.65
R176 VPWR.n33 VPWR.n32 3.388
R177 VPWR.n16 VPWR.n15 0.864
R178 VPWR.n49 VPWR.n48 0.752
R179 VPWR.n21 VPWR.n20 0.521
R180 VPWR.n37 VPWR.n36 0.376
R181 VPWR.n14 VPWR.n13 0.285
R182 VPWR.n25 VPWR.n23 0.143
R183 VPWR.n28 VPWR.n25 0.119
R184 VPWR.n30 VPWR.n28 0.119
R185 VPWR.n34 VPWR.n30 0.119
R186 VPWR.n38 VPWR.n34 0.119
R187 VPWR.n40 VPWR.n38 0.119
R188 VPWR.n44 VPWR.n40 0.119
R189 VPWR.n46 VPWR.n44 0.119
R190 VPWR.n50 VPWR.n46 0.119
R191 VPWR.n51 VPWR.n50 0.119
R192 VPWR.n23 VPWR.n21 0.1
R193 VPWR.n11 VPWR.n7 0.095
R194 VPWR.n20 VPWR.n16 0.092
R195 VPWR.n20 VPWR.n19 0.061
R196 VPWR VPWR.n51 0.02
R197 VPWR.n5 VPWR.n4 0.017
R198 VPWR.n3 VPWR.n2 0.017
R199 VPWR.n1 VPWR.n0 0.016
R200 VPWR.n4 VPWR.n3 0.014
R201 VPWR.n19 VPWR.n18 0.011
R202 VPWR.n18 VPWR.n17 0.008
R203 VPWR.n13 VPWR.n12 0.005
R204 VPWR.n10 VPWR.n9 0.005
R205 VPWR.n15 VPWR.n14 0.004
R206 VPWR.n14 VPWR.n5 0.003
R207 VPWR.n2 VPWR.n1 0.003
R208 VPWR.n13 VPWR.n6 0.003
R209 VPWR.n9 VPWR.n8 0.003
R210 VPWR.n12 VPWR.n11 0.001
R211 VPWR.n11 VPWR.n10 0.001
R212 VPB.t4 VPB.t5 248.598
R213 VPB.t3 VPB.t4 248.598
R214 VPB.t2 VPB.t3 248.598
R215 VPB.t1 VPB.t2 248.598
R216 VPB.t0 VPB.t1 248.598
R217 VPB.t7 VPB.t0 248.598
R218 VPB.t6 VPB.t7 248.598
R219 VPB.t8 VPB.t6 248.598
R220 VPB.t9 VPB.t8 248.598
R221 VPB.t10 VPB.t9 248.598
R222 VPB VPB.t10 189.408
R223 A.n6 A.t4 235.762
R224 A.n0 A.t0 221.719
R225 A.n2 A.t1 221.719
R226 A.n6 A.t5 163.462
R227 A.n0 A.t3 149.419
R228 A.n2 A.t2 149.419
R229 A.n5 A.n4 76
R230 A.n7 A.n6 76
R231 A.n1 A.n0 58.018
R232 A.n5 A.n2 43.737
R233 A.n4 A.n3 21.76
R234 A.n7 A 19.52
R235 A.n6 A.n5 17.851
R236 A.n2 A.n1 16.959
R237 A A.n7 9.92
R238 A.n3 A 5.44
R239 A.n4 A 2.24
C0 VPWR VGND 0.38fF
C1 VPB VPWR 0.15fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__sdfbbn_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__sdfbbn_1 SCD SCE RESET_B VGND CLK_N SET_B Q VPWR D Q_N VNB
+ VPB
X0 a_381_363.t1 SCD.t0 VPWR.t15 VPB.t23 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1 a_1102_21.t0 SET_B.t0 VPWR.t12 VPB.t17 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 VPWR.t1 a_1396_21.t2 a_2122_329.t1 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X3 Q.t0 a_2596_47.t2 VPWR.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 a_917_47.t2 a_27_47.t2 a_453_47.t3 VPB.t20 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 VPWR.t2 a_1396_21.t3 a_1351_329.t1 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X6 VPWR.t3 SCE.t0 a_423_315.t0 VPB.t5 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7 VGND.t13 SCE.t1 a_423_315.t1 VNB.t23 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 a_1030_47.t0 a_27_47.t3 a_917_47.t3 VNB.t7 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X9 a_1614_47.t1 a_1102_21.t4 VGND.t9 VNB.t16 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X10 a_1351_329.t0 a_917_47.t4 a_1102_21.t2 VPB.t7 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X11 VPWR.t9 RESET_B.t0 a_1396_21.t0 VPB.t14 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X12 VPWR.t8 CLK_N.t0 a_27_47.t0 VPB.t13 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X13 a_1572_329.t1 a_1102_21.t5 VPWR.t10 VPB.t15 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X14 a_2122_329.t0 a_1714_47.t4 a_1887_21.t1 VPB.t12 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X15 VGND.t4 a_1887_21.t4 a_1822_47.t0 VNB.t9 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16 VPWR.t11 a_1102_21.t6 a_1017_413.t1 VPB.t16 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17 VPWR.t5 a_1887_21.t5 a_1800_413.t0 VPB.t9 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18 a_1887_21.t2 a_1714_47.t5 a_2004_47.t1 VNB.t12 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X19 a_1887_21.t0 SET_B.t1 VPWR.t13 VPB.t18 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20 a_1800_413.t1 a_27_47.t4 a_1714_47.t3 VPB.t21 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21 a_1102_21.t3 a_917_47.t5 a_1241_47.t1 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X22 a_193_47.t1 a_27_47.t5 VGND.t2 VNB.t6 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23 a_453_47.t4 D.t0 a_735_47.t0 VNB.t17 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24 a_1714_47.t0 a_193_47.t2 a_1572_329.t0 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X25 a_2004_47.t2 a_1396_21.t4 a_1887_21.t3 VNB.t19 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X26 Q.t1 a_2596_47.t3 VGND.t3 VNB.t8 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X27 VGND.t5 a_1887_21.t6 a_2596_47.t0 VNB.t10 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X28 a_193_47.t0 a_27_47.t6 VPWR.t14 VPB.t22 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X29 a_1241_47.t0 SET_B.t2 VGND.t1 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X30 a_1241_47.t2 a_1396_21.t5 a_1102_21.t1 VNB.t18 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X31 a_1017_413.t0 a_193_47.t3 a_917_47.t0 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X32 VGND.t10 a_1102_21.t7 a_1030_47.t1 VNB.t15 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X33 a_735_47.t1 a_423_315.t2 VGND.t11 VNB.t20 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X34 VPWR.t6 a_1887_21.t7 a_2596_47.t1 VPB.t10 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X35 a_453_47.t2 a_423_315.t3 a_381_363.t0 VPB.t8 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X36 a_381_47.t0 SCD.t1 VGND.t12 VNB.t21 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X37 a_1714_47.t2 a_27_47.t7 a_1614_47.t0 VNB.t5 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X38 a_1822_47.t1 a_193_47.t4 a_1714_47.t1 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X39 Q_N.t1 a_1887_21.t8 VGND.t6 VNB.t11 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X40 a_917_47.t1 a_193_47.t5 a_453_47.t0 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X41 Q_N.t0 a_1887_21.t9 VPWR.t7 VPB.t11 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X42 a_453_47.t5 D.t1 a_752_413.t0 VPB.t19 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X43 a_2004_47.t0 SET_B.t3 VGND.t0 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X44 a_752_413.t1 SCE.t2 VPWR.t4 VPB.t6 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X45 VGND.t7 CLK_N.t1 a_27_47.t1 VNB.t13 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X46 a_453_47.t1 SCE.t3 a_381_47.t1 VNB.t22 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X47 VGND.t8 RESET_B.t1 a_1396_21.t1 VNB.t14 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
R0 SCD.n0 SCD.t1 301.529
R1 SCD.n0 SCD.t0 197.618
R2 SCD SCD.n0 78.057
R3 VPWR.n6 VPWR.t1 500.865
R4 VPWR.n1 VPWR.n0 440.25
R5 VPWR.n60 VPWR.n59 311.893
R6 VPWR.n47 VPWR.n46 308.79
R7 VPWR.n36 VPWR.n35 306.984
R8 VPWR.n14 VPWR.n13 292.5
R9 VPWR.n55 VPWR.t15 228.496
R10 VPWR.n3 VPWR.n2 173.154
R11 VPWR.n28 VPWR.n27 164.214
R12 VPWR.n13 VPWR.t13 91.464
R13 VPWR.n13 VPWR.t5 91.464
R14 VPWR.n35 VPWR.t12 91.464
R15 VPWR.n27 VPWR.t10 86.773
R16 VPWR.n35 VPWR.t11 86.773
R17 VPWR.n46 VPWR.t4 63.321
R18 VPWR.n46 VPWR.t3 63.321
R19 VPWR.n0 VPWR.t9 63.101
R20 VPWR.n2 VPWR.t6 57.733
R21 VPWR.n59 VPWR.t14 41.554
R22 VPWR.n59 VPWR.t8 41.554
R23 VPWR.n27 VPWR.t2 38.696
R24 VPWR.n2 VPWR.t0 32.579
R25 VPWR.n0 VPWR.t7 28.032
R26 VPWR.n5 VPWR.n4 4.65
R27 VPWR.n8 VPWR.n7 4.65
R28 VPWR.n10 VPWR.n9 4.65
R29 VPWR.n12 VPWR.n11 4.65
R30 VPWR.n16 VPWR.n15 4.65
R31 VPWR.n18 VPWR.n17 4.65
R32 VPWR.n20 VPWR.n19 4.65
R33 VPWR.n22 VPWR.n21 4.65
R34 VPWR.n24 VPWR.n23 4.65
R35 VPWR.n26 VPWR.n25 4.65
R36 VPWR.n30 VPWR.n29 4.65
R37 VPWR.n32 VPWR.n31 4.65
R38 VPWR.n34 VPWR.n33 4.65
R39 VPWR.n37 VPWR.n36 4.65
R40 VPWR.n39 VPWR.n38 4.65
R41 VPWR.n41 VPWR.n40 4.65
R42 VPWR.n43 VPWR.n42 4.65
R43 VPWR.n45 VPWR.n44 4.65
R44 VPWR.n48 VPWR.n47 4.65
R45 VPWR.n50 VPWR.n49 4.65
R46 VPWR.n52 VPWR.n51 4.65
R47 VPWR.n54 VPWR.n53 4.65
R48 VPWR.n56 VPWR.n55 4.65
R49 VPWR.n58 VPWR.n57 4.65
R50 VPWR.n3 VPWR.n1 4.611
R51 VPWR.n61 VPWR.n60 3.932
R52 VPWR.n7 VPWR.n6 3.84
R53 VPWR.n29 VPWR.n28 3.388
R54 VPWR.n15 VPWR.n14 2.443
R55 VPWR.n5 VPWR.n3 0.144
R56 VPWR.n61 VPWR.n58 0.137
R57 VPWR VPWR.n61 0.123
R58 VPWR.n8 VPWR.n5 0.119
R59 VPWR.n10 VPWR.n8 0.119
R60 VPWR.n12 VPWR.n10 0.119
R61 VPWR.n16 VPWR.n12 0.119
R62 VPWR.n18 VPWR.n16 0.119
R63 VPWR.n20 VPWR.n18 0.119
R64 VPWR.n22 VPWR.n20 0.119
R65 VPWR.n24 VPWR.n22 0.119
R66 VPWR.n26 VPWR.n24 0.119
R67 VPWR.n30 VPWR.n26 0.119
R68 VPWR.n32 VPWR.n30 0.119
R69 VPWR.n34 VPWR.n32 0.119
R70 VPWR.n37 VPWR.n34 0.119
R71 VPWR.n39 VPWR.n37 0.119
R72 VPWR.n41 VPWR.n39 0.119
R73 VPWR.n43 VPWR.n41 0.119
R74 VPWR.n45 VPWR.n43 0.119
R75 VPWR.n48 VPWR.n45 0.119
R76 VPWR.n50 VPWR.n48 0.119
R77 VPWR.n52 VPWR.n50 0.119
R78 VPWR.n54 VPWR.n52 0.119
R79 VPWR.n56 VPWR.n54 0.119
R80 VPWR.n58 VPWR.n56 0.119
R81 a_381_363.t0 a_381_363.t1 64.64
R82 VPB.t8 VPB.t5 636.292
R83 VPB.t1 VPB.t14 588.94
R84 VPB.t11 VPB.t10 556.386
R85 VPB.t22 VPB.t23 556.386
R86 VPB.t15 VPB.t3 426.168
R87 VPB.t2 VPB.t15 405.451
R88 VPB.t4 VPB.t16 355.14
R89 VPB.t21 VPB.t9 349.221
R90 VPB.t9 VPB.t18 319.626
R91 VPB.t17 VPB.t7 319.626
R92 VPB.t16 VPB.t17 313.707
R93 VPB.t14 VPB.t11 287.071
R94 VPB.t19 VPB.t20 287.071
R95 VPB.t18 VPB.t12 284.112
R96 VPB.t10 VPB.t0 281.152
R97 VPB.t3 VPB.t21 248.598
R98 VPB.t7 VPB.t2 248.598
R99 VPB.t20 VPB.t4 248.598
R100 VPB.t6 VPB.t19 248.598
R101 VPB.t5 VPB.t6 248.598
R102 VPB.t13 VPB.t22 248.598
R103 VPB.t12 VPB.t1 213.084
R104 VPB.t23 VPB.t8 213.084
R105 VPB VPB.t13 142.056
R106 SET_B.n0 SET_B.t0 438.597
R107 SET_B.n1 SET_B.t1 393.971
R108 SET_B.n0 SET_B.t2 142.633
R109 SET_B.n1 SET_B.t3 134.267
R110 SET_B.n2 SET_B.n0 80.823
R111 SET_B.n2 SET_B.n1 17.667
R112 SET_B SET_B.n2 5.008
R113 SET_B.n2 SET_B 3.153
R114 a_1102_21.n5 a_1102_21.t7 386.158
R115 a_1102_21.n2 a_1102_21.t5 299.91
R116 a_1102_21.n7 a_1102_21.n6 292.5
R117 a_1102_21.n2 a_1102_21.t4 167.627
R118 a_1102_21.n5 a_1102_21.t6 141.945
R119 a_1102_21.n4 a_1102_21.n2 141.698
R120 a_1102_21.n6 a_1102_21.n5 114.656
R121 a_1102_21.n4 a_1102_21.n3 111.206
R122 a_1102_21.n0 a_1102_21.t0 110.226
R123 a_1102_21.n6 a_1102_21.n4 81.806
R124 a_1102_21.t2 a_1102_21.n1 63.321
R125 a_1102_21.t2 a_1102_21.n7 63.321
R126 a_1102_21.n3 a_1102_21.t1 25.312
R127 a_1102_21.n3 a_1102_21.t3 25.312
R128 a_1102_21.n1 a_1102_21.n0 9.38
R129 a_1396_21.t0 a_1396_21.n3 448.039
R130 a_1396_21.n0 a_1396_21.t5 212.988
R131 a_1396_21.n1 a_1396_21.t4 211.511
R132 a_1396_21.n1 a_1396_21.t2 206.934
R133 a_1396_21.n0 a_1396_21.t3 204.868
R134 a_1396_21.n2 a_1396_21.t1 194.213
R135 a_1396_21.n3 a_1396_21.n0 126.544
R136 a_1396_21.n2 a_1396_21.n1 76
R137 a_1396_21.n3 a_1396_21.n2 9.774
R138 a_2122_329.t0 a_2122_329.t1 49.25
R139 a_2596_47.n0 a_2596_47.t2 239.503
R140 a_2596_47.t1 a_2596_47.n1 237.868
R141 a_2596_47.n0 a_2596_47.t3 167.203
R142 a_2596_47.n1 a_2596_47.t0 150.778
R143 a_2596_47.n1 a_2596_47.n0 99.078
R144 Q.n1 Q.t0 207.372
R145 Q.n0 Q.t1 117.423
R146 Q Q.n0 68.335
R147 Q.n1 Q 9.019
R148 Q Q.n1 7.458
R149 Q.n0 Q 6.646
R150 a_27_47.n2 a_27_47.t2 498.224
R151 a_27_47.t0 a_27_47.n5 274.546
R152 a_27_47.n1 a_27_47.t4 267.397
R153 a_27_47.n0 a_27_47.t6 262.942
R154 a_27_47.n0 a_27_47.t5 227.596
R155 a_27_47.n1 a_27_47.t7 207.657
R156 a_27_47.n4 a_27_47.t1 168.633
R157 a_27_47.n2 a_27_47.t3 133.466
R158 a_27_47.n5 a_27_47.n0 76
R159 a_27_47.n5 a_27_47.n4 21.426
R160 a_27_47.n3 a_27_47.n2 10.359
R161 a_27_47.n4 a_27_47.n3 8.606
R162 a_27_47.n3 a_27_47.n1 7.542
R163 a_453_47.n2 a_453_47.n0 370.577
R164 a_453_47.t2 a_453_47.n3 277.904
R165 a_453_47.n3 a_453_47.t1 198.545
R166 a_453_47.n2 a_453_47.n1 163.58
R167 a_453_47.n0 a_453_47.t3 93.809
R168 a_453_47.n1 a_453_47.t0 63.333
R169 a_453_47.n0 a_453_47.t5 63.321
R170 a_453_47.n1 a_453_47.t4 29.726
R171 a_453_47.n3 a_453_47.n2 25.313
R172 a_917_47.n3 a_917_47.n2 412.288
R173 a_917_47.n1 a_917_47.t5 220.704
R174 a_917_47.n1 a_917_47.t4 214.132
R175 a_917_47.n2 a_917_47.n0 201.436
R176 a_917_47.n2 a_917_47.n1 144.216
R177 a_917_47.n0 a_917_47.t3 93.333
R178 a_917_47.t0 a_917_47.n3 63.321
R179 a_917_47.n3 a_917_47.t2 63.321
R180 a_917_47.n0 a_917_47.t1 45
R181 a_1351_329.t0 a_1351_329.t1 63.321
R182 SCE.n2 SCE.n1 285.986
R183 SCE.n3 SCE.n2 266.589
R184 SCE.n1 SCE.t2 228.146
R185 SCE.n3 SCE.t3 97.831
R186 SCE.n2 SCE.t1 93.186
R187 SCE.n1 SCE.t0 93.186
R188 SCE.n4 SCE.n3 76
R189 SCE SCE.n4 28.416
R190 SCE.n0 SCE 17.163
R191 SCE.n4 SCE 4.042
R192 SCE.n0 SCE 2.618
R193 SCE SCE.n0 1.515
R194 a_423_315.n1 a_423_315.t3 402.702
R195 a_423_315.t0 a_423_315.n1 385.562
R196 a_423_315.n0 a_423_315.t2 208.281
R197 a_423_315.n0 a_423_315.t1 191.602
R198 a_423_315.n1 a_423_315.n0 76.279
R199 VGND.n24 VGND.t9 186.97
R200 VGND.n54 VGND.t12 152.947
R201 VGND.n34 VGND.n33 113.205
R202 VGND.n3 VGND.n0 113.067
R203 VGND.n13 VGND.n12 110.223
R204 VGND.n59 VGND.n58 107.239
R205 VGND.n46 VGND.n45 106.463
R206 VGND.n33 VGND.t10 74.285
R207 VGND.n2 VGND.n1 64.275
R208 VGND.n1 VGND.t8 57.796
R209 VGND.n0 VGND.t5 54.285
R210 VGND.n12 VGND.t4 42.857
R211 VGND.n45 VGND.t13 42.857
R212 VGND.n12 VGND.t0 38.571
R213 VGND.n33 VGND.t1 38.571
R214 VGND.n45 VGND.t11 38.571
R215 VGND.n58 VGND.t2 38.571
R216 VGND.n58 VGND.t7 38.571
R217 VGND.n0 VGND.t3 25.934
R218 VGND.n1 VGND.t6 24.765
R219 VGND.n35 VGND.n34 12.8
R220 VGND.n14 VGND.n13 5.27
R221 VGND.n5 VGND.n4 4.65
R222 VGND.n7 VGND.n6 4.65
R223 VGND.n9 VGND.n8 4.65
R224 VGND.n11 VGND.n10 4.65
R225 VGND.n15 VGND.n14 4.65
R226 VGND.n17 VGND.n16 4.65
R227 VGND.n19 VGND.n18 4.65
R228 VGND.n21 VGND.n20 4.65
R229 VGND.n23 VGND.n22 4.65
R230 VGND.n26 VGND.n25 4.65
R231 VGND.n28 VGND.n27 4.65
R232 VGND.n30 VGND.n29 4.65
R233 VGND.n32 VGND.n31 4.65
R234 VGND.n36 VGND.n35 4.65
R235 VGND.n38 VGND.n37 4.65
R236 VGND.n40 VGND.n39 4.65
R237 VGND.n42 VGND.n41 4.65
R238 VGND.n44 VGND.n43 4.65
R239 VGND.n47 VGND.n46 4.65
R240 VGND.n49 VGND.n48 4.65
R241 VGND.n51 VGND.n50 4.65
R242 VGND.n53 VGND.n52 4.65
R243 VGND.n55 VGND.n54 4.65
R244 VGND.n57 VGND.n56 4.65
R245 VGND.n3 VGND.n2 3.969
R246 VGND.n60 VGND.n59 3.932
R247 VGND.n25 VGND.n24 2.258
R248 VGND.n5 VGND.n3 0.146
R249 VGND.n60 VGND.n57 0.137
R250 VGND VGND.n60 0.123
R251 VGND.n7 VGND.n5 0.119
R252 VGND.n9 VGND.n7 0.119
R253 VGND.n11 VGND.n9 0.119
R254 VGND.n15 VGND.n11 0.119
R255 VGND.n17 VGND.n15 0.119
R256 VGND.n19 VGND.n17 0.119
R257 VGND.n21 VGND.n19 0.119
R258 VGND.n23 VGND.n21 0.119
R259 VGND.n26 VGND.n23 0.119
R260 VGND.n28 VGND.n26 0.119
R261 VGND.n30 VGND.n28 0.119
R262 VGND.n32 VGND.n30 0.119
R263 VGND.n36 VGND.n32 0.119
R264 VGND.n38 VGND.n36 0.119
R265 VGND.n40 VGND.n38 0.119
R266 VGND.n42 VGND.n40 0.119
R267 VGND.n44 VGND.n42 0.119
R268 VGND.n47 VGND.n44 0.119
R269 VGND.n49 VGND.n47 0.119
R270 VGND.n51 VGND.n49 0.119
R271 VGND.n53 VGND.n51 0.119
R272 VGND.n55 VGND.n53 0.119
R273 VGND.n57 VGND.n55 0.119
R274 VNB.t22 VNB.t23 6308.82
R275 VNB.t6 VNB.t21 6082.35
R276 VNB.t19 VNB.t14 4595.56
R277 VNB.t18 VNB.t16 4595.56
R278 VNB.t11 VNB.t10 4545.05
R279 VNB VNB.t13 4270.59
R280 VNB.t3 VNB.t7 3655.88
R281 VNB.t15 VNB.t1 3526.47
R282 VNB.t5 VNB.t2 3494.12
R283 VNB.t7 VNB.t15 3300
R284 VNB.t2 VNB.t9 3073.53
R285 VNB.t17 VNB.t3 3073.53
R286 VNB.t0 VNB.t12 3065.62
R287 VNB.t9 VNB.t0 2814.71
R288 VNB.t20 VNB.t17 2814.71
R289 VNB.t23 VNB.t20 2814.71
R290 VNB.t13 VNB.t6 2717.65
R291 VNB.t1 VNB.t4 2363.68
R292 VNB.t16 VNB.t5 2349.76
R293 VNB.t21 VNB.t22 2329.41
R294 VNB.t14 VNB.t11 2296.97
R295 VNB.t10 VNB.t8 2296.7
R296 VNB.t12 VNB.t19 2053.33
R297 VNB.t4 VNB.t18 2053.33
R298 a_1030_47.t1 a_1030_47.t0 99.046
R299 a_1614_47.n0 a_1614_47.t0 75
R300 a_1614_47.n1 a_1614_47.n0 67.2
R301 a_1614_47.n0 a_1614_47.t1 13.143
R302 RESET_B.n0 RESET_B.t1 203.042
R303 RESET_B.n0 RESET_B.t0 174.121
R304 RESET_B RESET_B.n0 78.109
R305 CLK_N.n0 CLK_N.t0 272.06
R306 CLK_N.n0 CLK_N.t1 236.714
R307 CLK_N.n1 CLK_N.n0 76
R308 CLK_N CLK_N.n1 7.68
R309 CLK_N.n1 CLK_N 4.754
R310 a_1572_329.t1 a_1572_329.t0 236.868
R311 a_1714_47.n3 a_1714_47.n2 399.793
R312 a_1714_47.n1 a_1714_47.t4 241.535
R313 a_1714_47.n1 a_1714_47.t5 196.547
R314 a_1714_47.n2 a_1714_47.n0 183.436
R315 a_1714_47.n2 a_1714_47.n1 159.918
R316 a_1714_47.n0 a_1714_47.t2 70
R317 a_1714_47.n3 a_1714_47.t3 63.321
R318 a_1714_47.t0 a_1714_47.n3 63.321
R319 a_1714_47.n0 a_1714_47.t1 60
R320 a_1887_21.n5 a_1887_21.t4 386.846
R321 a_1887_21.n7 a_1887_21.n6 301.911
R322 a_1887_21.n1 a_1887_21.t9 292.412
R323 a_1887_21.n0 a_1887_21.t7 231.942
R324 a_1887_21.n4 a_1887_21.n2 229.286
R325 a_1887_21.n1 a_1887_21.t8 220.112
R326 a_1887_21.n4 a_1887_21.n3 185.612
R327 a_1887_21.n0 a_1887_21.t6 164.463
R328 a_1887_21.n2 a_1887_21.n0 151.74
R329 a_1887_21.n5 a_1887_21.t5 142.633
R330 a_1887_21.n6 a_1887_21.n5 128.841
R331 a_1887_21.n7 a_1887_21.t0 91.464
R332 a_1887_21.t1 a_1887_21.n7 32.833
R333 a_1887_21.n6 a_1887_21.n4 30.494
R334 a_1887_21.n3 a_1887_21.t3 25.312
R335 a_1887_21.n3 a_1887_21.t2 25.312
R336 a_1887_21.n2 a_1887_21.n1 2.677
R337 a_1822_47.t0 a_1822_47.t1 93.059
R338 a_1017_413.t0 a_1017_413.t1 211.071
R339 a_1800_413.t0 a_1800_413.t1 206.38
R340 a_2004_47.n0 a_2004_47.t2 270.96
R341 a_2004_47.n0 a_2004_47.t0 64.285
R342 a_2004_47.t1 a_2004_47.n0 47.722
R343 a_1241_47.n0 a_1241_47.t2 280.603
R344 a_1241_47.n0 a_1241_47.t0 62.857
R345 a_1241_47.t1 a_1241_47.n0 26.294
R346 a_193_47.n0 a_193_47.t4 532.86
R347 a_193_47.n1 a_193_47.t5 245.063
R348 a_193_47.n1 a_193_47.t3 231.324
R349 a_193_47.n3 a_193_47.t1 210.124
R350 a_193_47.n0 a_193_47.t2 137.933
R351 a_193_47.t0 a_193_47.n3 121.825
R352 a_193_47.n2 a_193_47.n0 12.947
R353 a_193_47.n3 a_193_47.n2 4.716
R354 a_193_47.n2 a_193_47.n1 4.65
R355 D.n0 D.t0 308.479
R356 D.n0 D.t1 224.932
R357 D.n1 D.n0 76
R358 D D.n1 24.51
R359 D.n1 D 5.451
R360 a_735_47.t0 a_735_47.t1 81.428
R361 a_381_47.t0 a_381_47.t1 60
R362 Q_N.n1 Q_N.t0 207.566
R363 Q_N.n0 Q_N.t1 117.423
R364 Q_N Q_N.n0 79.437
R365 Q_N.n1 Q_N 8.185
R366 Q_N Q_N.n1 6.859
R367 Q_N.n0 Q_N 5.614
R368 a_752_413.t0 a_752_413.t1 126.642
C0 SCD SCE 0.11fF
C1 SET_B VGND 0.36fF
C2 VPB VPWR 0.30fF
C3 VPWR Q 0.14fF
C4 VGND Q_N 0.12fF
C5 VPWR VGND 0.14fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__sdfbbn_2.ext - technology: sky130A

.subckt sky130_fd_sc_hd__sdfbbn_2 SCD SCE RESET_B VGND CLK_N SET_B Q VPWR D Q_N VNB
+ VPB
X0 a_381_363.t1 SCD.t0 VPWR.t16 VPB.t20 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1 a_1107_21.t0 SET_B.t0 VPWR.t12 VPB.t15 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 VPWR.t8 a_1401_21.t2 a_2122_329.t0 VPB.t11 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X3 a_1251_47.t1 a_1401_21.t3 a_1107_21.t1 VNB.t15 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X4 a_931_47.t2 a_27_47.t2 a_453_47.t4 VPB.t23 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 VPWR.t9 a_1401_21.t4 a_1351_329.t0 VPB.t12 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X6 VPWR.t3 SCE.t0 a_423_315.t0 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7 a_1351_329.t1 a_931_47.t4 a_1107_21.t2 VPB.t21 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X8 VPWR.t5 CLK_N.t0 a_27_47.t1 VPB.t5 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X9 a_1572_329.t1 a_1107_21.t4 VPWR.t10 VPB.t13 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X10 a_2122_329.t1 a_1714_47.t4 a_1888_21.t1 VPB.t22 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X11 VGND.t9 a_1888_21.t4 a_1823_47.t1 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12 a_1041_47.t1 a_27_47.t3 a_931_47.t3 VNB.t21 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X13 a_1107_21.t3 a_931_47.t5 a_1251_47.t2 VNB.t15 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X14 VPWR.t11 a_1107_21.t5 a_1017_413.t1 VPB.t14 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15 VPWR.t1 a_1888_21.t5 a_1800_413.t0 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16 a_1888_21.t2 a_1714_47.t5 a_2004_47.t1 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X17 a_764_47.t1 a_423_315.t2 VGND.t15 VNB.t12 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18 Q.t3 a_2696_47.t2 VGND.t7 VNB.t17 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X19 a_1888_21.t0 SET_B.t1 VPWR.t13 VPB.t16 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20 a_931_47.t0 a_193_47.t2 a_453_47.t1 VNB.t6 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X21 a_1800_413.t1 a_27_47.t4 a_1714_47.t3 VPB.t24 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22 VGND.t10 a_1888_21.t6 a_2696_47.t1 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23 a_193_47.t1 a_27_47.t5 VGND.t13 VNB.t22 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24 VPWR.t0 a_1888_21.t7 a_2696_47.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X25 a_453_47.t5 D.t0 a_764_47.t0 VNB.t20 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X26 VGND.t0 SCE.t1 a_423_315.t1 VNB.t5 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X27 a_1714_47.t0 a_193_47.t3 a_1572_329.t0 VPB.t9 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X28 VPWR.t15 a_1888_21.t8 Q_N.t1 VPB.t18 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X29 a_2004_47.t2 a_1401_21.t5 a_1888_21.t3 VNB.t19 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X30 VGND.t5 a_1107_21.t6 a_1041_47.t0 VNB.t16 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X31 VGND.t12 a_1888_21.t9 Q_N.t3 VNB.t11 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X32 VGND.t8 a_2696_47.t3 Q.t2 VNB.t18 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X33 VPWR.t6 a_2696_47.t4 Q.t1 VPB.t7 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X34 Q_N.t0 a_1888_21.t10 VPWR.t2 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X35 a_193_47.t0 a_27_47.t6 VPWR.t17 VPB.t25 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X36 Q.t0 a_2696_47.t5 VPWR.t7 VPB.t8 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X37 a_1017_413.t0 a_193_47.t4 a_931_47.t1 VPB.t10 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X38 a_1823_47.t0 a_193_47.t5 a_1714_47.t1 VNB.t8 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X39 Q_N.t2 a_1888_21.t11 VGND.t11 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X40 a_453_47.t2 a_423_315.t3 a_381_363.t0 VPB.t19 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X41 a_381_47.t1 SCD.t1 VGND.t4 VNB.t14 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X42 a_1714_47.t2 a_27_47.t7 a_1619_47.t1 VNB.t23 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X43 a_453_47.t0 D.t1 a_752_413.t1 VPB.t6 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X44 a_1251_47.t0 SET_B.t2 VGND.t3 VNB.t10 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X45 a_1619_47.t0 a_1107_21.t7 VGND.t6 VNB.t15 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X46 a_2004_47.t0 SET_B.t3 VGND.t2 VNB.t9 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X47 VPWR.t14 RESET_B.t0 a_1401_21.t1 VPB.t17 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X48 VGND.t1 RESET_B.t1 a_1401_21.t0 VNB.t7 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X49 a_752_413.t0 SCE.t2 VPWR.t4 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X50 VGND.t14 CLK_N.t1 a_27_47.t0 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X51 a_453_47.t3 SCE.t3 a_381_47.t0 VNB.t13 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
R0 SCD.n0 SCD.t1 301.268
R1 SCD.n0 SCD.t0 172.734
R2 SCD SCD.n0 78.057
R3 VPWR.n15 VPWR.t8 500.865
R4 VPWR.n10 VPWR.n9 440.25
R5 VPWR.n69 VPWR.n68 311.893
R6 VPWR.n56 VPWR.n55 308.082
R7 VPWR.n45 VPWR.n44 306.984
R8 VPWR.n23 VPWR.n22 292.5
R9 VPWR.n64 VPWR.t16 228.496
R10 VPWR.n1 VPWR.n0 168.939
R11 VPWR.n37 VPWR.n36 164.214
R12 VPWR.n2 VPWR.t6 157.987
R13 VPWR.n5 VPWR.t15 154.509
R14 VPWR.n22 VPWR.t13 91.464
R15 VPWR.n22 VPWR.t1 91.464
R16 VPWR.n44 VPWR.t12 91.464
R17 VPWR.n36 VPWR.t10 86.773
R18 VPWR.n44 VPWR.t11 86.773
R19 VPWR.n55 VPWR.t4 63.321
R20 VPWR.n55 VPWR.t3 63.321
R21 VPWR.n9 VPWR.t14 63.101
R22 VPWR.n0 VPWR.t0 58.484
R23 VPWR.n68 VPWR.t17 41.554
R24 VPWR.n68 VPWR.t5 41.554
R25 VPWR.n36 VPWR.t9 38.696
R26 VPWR.n0 VPWR.t7 31.83
R27 VPWR.n9 VPWR.t2 27.786
R28 VPWR.n4 VPWR.n3 4.65
R29 VPWR.n6 VPWR.n5 4.65
R30 VPWR.n8 VPWR.n7 4.65
R31 VPWR.n12 VPWR.n11 4.65
R32 VPWR.n14 VPWR.n13 4.65
R33 VPWR.n17 VPWR.n16 4.65
R34 VPWR.n19 VPWR.n18 4.65
R35 VPWR.n21 VPWR.n20 4.65
R36 VPWR.n25 VPWR.n24 4.65
R37 VPWR.n27 VPWR.n26 4.65
R38 VPWR.n29 VPWR.n28 4.65
R39 VPWR.n31 VPWR.n30 4.65
R40 VPWR.n33 VPWR.n32 4.65
R41 VPWR.n35 VPWR.n34 4.65
R42 VPWR.n39 VPWR.n38 4.65
R43 VPWR.n41 VPWR.n40 4.65
R44 VPWR.n43 VPWR.n42 4.65
R45 VPWR.n46 VPWR.n45 4.65
R46 VPWR.n48 VPWR.n47 4.65
R47 VPWR.n50 VPWR.n49 4.65
R48 VPWR.n52 VPWR.n51 4.65
R49 VPWR.n54 VPWR.n53 4.65
R50 VPWR.n57 VPWR.n56 4.65
R51 VPWR.n59 VPWR.n58 4.65
R52 VPWR.n61 VPWR.n60 4.65
R53 VPWR.n63 VPWR.n62 4.65
R54 VPWR.n65 VPWR.n64 4.65
R55 VPWR.n67 VPWR.n66 4.65
R56 VPWR.n70 VPWR.n69 3.932
R57 VPWR.n16 VPWR.n15 3.84
R58 VPWR.n2 VPWR.n1 3.73
R59 VPWR.n38 VPWR.n37 3.388
R60 VPWR.n24 VPWR.n23 2.443
R61 VPWR.n11 VPWR.n10 1.28
R62 VPWR.n4 VPWR.n2 0.247
R63 VPWR.n70 VPWR.n67 0.137
R64 VPWR VPWR.n70 0.123
R65 VPWR.n6 VPWR.n4 0.119
R66 VPWR.n8 VPWR.n6 0.119
R67 VPWR.n12 VPWR.n8 0.119
R68 VPWR.n14 VPWR.n12 0.119
R69 VPWR.n17 VPWR.n14 0.119
R70 VPWR.n19 VPWR.n17 0.119
R71 VPWR.n21 VPWR.n19 0.119
R72 VPWR.n25 VPWR.n21 0.119
R73 VPWR.n27 VPWR.n25 0.119
R74 VPWR.n29 VPWR.n27 0.119
R75 VPWR.n31 VPWR.n29 0.119
R76 VPWR.n33 VPWR.n31 0.119
R77 VPWR.n35 VPWR.n33 0.119
R78 VPWR.n39 VPWR.n35 0.119
R79 VPWR.n41 VPWR.n39 0.119
R80 VPWR.n43 VPWR.n41 0.119
R81 VPWR.n46 VPWR.n43 0.119
R82 VPWR.n48 VPWR.n46 0.119
R83 VPWR.n50 VPWR.n48 0.119
R84 VPWR.n52 VPWR.n50 0.119
R85 VPWR.n54 VPWR.n52 0.119
R86 VPWR.n57 VPWR.n54 0.119
R87 VPWR.n59 VPWR.n57 0.119
R88 VPWR.n61 VPWR.n59 0.119
R89 VPWR.n63 VPWR.n61 0.119
R90 VPWR.n65 VPWR.n63 0.119
R91 VPWR.n67 VPWR.n65 0.119
R92 a_381_363.t0 a_381_363.t1 64.64
R93 VPB.t11 VPB.t17 636.292
R94 VPB.t19 VPB.t3 636.292
R95 VPB.t18 VPB.t0 556.386
R96 VPB.t25 VPB.t20 556.386
R97 VPB.t13 VPB.t9 426.168
R98 VPB.t12 VPB.t13 405.451
R99 VPB.t10 VPB.t14 355.14
R100 VPB.t24 VPB.t1 349.221
R101 VPB.t1 VPB.t16 319.626
R102 VPB.t15 VPB.t21 319.626
R103 VPB.t14 VPB.t15 313.707
R104 VPB.t17 VPB.t2 287.071
R105 VPB.t6 VPB.t23 287.071
R106 VPB.t16 VPB.t22 284.112
R107 VPB.t0 VPB.t8 281.152
R108 VPB.t8 VPB.t7 248.598
R109 VPB.t2 VPB.t18 248.598
R110 VPB.t9 VPB.t24 248.598
R111 VPB.t21 VPB.t12 248.598
R112 VPB.t23 VPB.t10 248.598
R113 VPB.t4 VPB.t6 248.598
R114 VPB.t3 VPB.t4 248.598
R115 VPB.t5 VPB.t25 248.598
R116 VPB.t22 VPB.t11 213.084
R117 VPB.t20 VPB.t19 213.084
R118 VPB VPB.t5 142.056
R119 SET_B.n0 SET_B.t0 396.831
R120 SET_B.n3 SET_B.t1 394.428
R121 SET_B.n3 SET_B.t3 134.495
R122 SET_B.n0 SET_B.t2 134.063
R123 SET_B SET_B.n6 13.6
R124 SET_B.n5 SET_B.n3 13.011
R125 SET_B.n1 SET_B.n0 6.985
R126 SET_B.n6 SET_B.n5 6.318
R127 SET_B.n6 SET_B.n1 2.521
R128 SET_B.n2 SET_B 2.521
R129 SET_B.n6 SET_B.n2 0.775
R130 SET_B.n5 SET_B.n4 0.001
R131 a_1107_21.n5 a_1107_21.t6 387.959
R132 a_1107_21.n2 a_1107_21.t4 299.91
R133 a_1107_21.n7 a_1107_21.n6 292.5
R134 a_1107_21.n2 a_1107_21.t7 167.627
R135 a_1107_21.n5 a_1107_21.t5 143.746
R136 a_1107_21.n4 a_1107_21.n2 139.816
R137 a_1107_21.n6 a_1107_21.n5 114.656
R138 a_1107_21.n0 a_1107_21.t0 110.226
R139 a_1107_21.n4 a_1107_21.n3 109.954
R140 a_1107_21.n6 a_1107_21.n4 81.172
R141 a_1107_21.t2 a_1107_21.n1 63.321
R142 a_1107_21.t2 a_1107_21.n7 63.321
R143 a_1107_21.n3 a_1107_21.t1 25.312
R144 a_1107_21.n3 a_1107_21.t3 25.312
R145 a_1107_21.n1 a_1107_21.n0 9.38
R146 a_1401_21.t1 a_1401_21.n3 454.063
R147 a_1401_21.n1 a_1401_21.t5 211.734
R148 a_1401_21.n1 a_1401_21.t2 207.402
R149 a_1401_21.n0 a_1401_21.t3 205.623
R150 a_1401_21.n0 a_1401_21.t4 204.868
R151 a_1401_21.n2 a_1401_21.t0 196.688
R152 a_1401_21.n3 a_1401_21.n0 126.544
R153 a_1401_21.n2 a_1401_21.n1 76
R154 a_1401_21.n3 a_1401_21.n2 9.774
R155 a_2122_329.t0 a_2122_329.t1 49.25
R156 a_1251_47.t1 a_1251_47.n0 283.512
R157 a_1251_47.n0 a_1251_47.t2 43.437
R158 a_1251_47.n0 a_1251_47.t0 38.571
R159 VNB.t13 VNB.t5 6858.82
R160 VNB.t22 VNB.t14 6082.35
R161 VNB.t19 VNB.t7 4962.22
R162 VNB.t11 VNB.t0 4545.05
R163 VNB VNB.t3 4270.59
R164 VNB.t16 VNB.t10 3688.24
R165 VNB.t6 VNB.t21 3558.82
R166 VNB.t23 VNB.t8 3526.47
R167 VNB.t5 VNB.t12 3202.94
R168 VNB.t21 VNB.t16 3105.88
R169 VNB.t9 VNB.t4 3097.97
R170 VNB.t8 VNB.t1 3073.53
R171 VNB.t20 VNB.t6 3073.53
R172 VNB.t1 VNB.t9 2782.35
R173 VNB.t3 VNB.t22 2717.65
R174 VNB.t12 VNB.t20 2329.41
R175 VNB.t14 VNB.t13 2329.41
R176 VNB.t7 VNB.t2 2296.97
R177 VNB.t0 VNB.t17 2296.7
R178 VNB.t4 VNB.t19 2053.33
R179 VNB.t17 VNB.t18 2030.77
R180 VNB.t2 VNB.t11 2030.77
R181 VNB.t10 VNB.t15 213.215
R182 VNB.t10 VNB.t23 40.121
R183 a_27_47.n2 a_27_47.t2 538.597
R184 a_27_47.t1 a_27_47.n5 278.108
R185 a_27_47.n1 a_27_47.t4 267.397
R186 a_27_47.n0 a_27_47.t6 262.942
R187 a_27_47.n0 a_27_47.t5 227.596
R188 a_27_47.n1 a_27_47.t7 207.297
R189 a_27_47.n4 a_27_47.t0 173.241
R190 a_27_47.n2 a_27_47.t3 135.786
R191 a_27_47.n5 a_27_47.n0 76
R192 a_27_47.n5 a_27_47.n4 21.426
R193 a_27_47.n3 a_27_47.n2 10.203
R194 a_27_47.n4 a_27_47.n3 8.649
R195 a_27_47.n3 a_27_47.n1 7.5
R196 a_453_47.n2 a_453_47.n0 355.646
R197 a_453_47.t2 a_453_47.n3 325.164
R198 a_453_47.n3 a_453_47.t3 190.315
R199 a_453_47.n2 a_453_47.n1 133.46
R200 a_453_47.n0 a_453_47.t4 93.809
R201 a_453_47.n1 a_453_47.t1 63.333
R202 a_453_47.n0 a_453_47.t0 63.321
R203 a_453_47.n1 a_453_47.t5 29.726
R204 a_453_47.n3 a_453_47.n2 24.429
R205 a_931_47.n3 a_931_47.n2 415.031
R206 a_931_47.n1 a_931_47.t5 216.899
R207 a_931_47.n1 a_931_47.t4 210.473
R208 a_931_47.n2 a_931_47.n0 196.424
R209 a_931_47.n2 a_931_47.n1 140.828
R210 a_931_47.n0 a_931_47.t0 70
R211 a_931_47.n0 a_931_47.t3 63.333
R212 a_931_47.t1 a_931_47.n3 63.321
R213 a_931_47.n3 a_931_47.t2 63.321
R214 a_1351_329.t0 a_1351_329.t1 63.321
R215 SCE.n1 SCE.n0 310.086
R216 SCE.n2 SCE.n1 290.404
R217 SCE.n0 SCE.t2 228.146
R218 SCE.n2 SCE.t3 101.219
R219 SCE.n0 SCE.t0 93.186
R220 SCE.n1 SCE.t1 93.186
R221 SCE.n3 SCE.n2 76
R222 SCE.n3 SCE 26.003
R223 SCE SCE.n3 5.861
R224 a_423_315.t0 a_423_315.n1 427.341
R225 a_423_315.n1 a_423_315.t3 391.928
R226 a_423_315.n0 a_423_315.t2 209.832
R227 a_423_315.n0 a_423_315.t1 192.057
R228 a_423_315.n1 a_423_315.n0 89.034
R229 CLK_N.n0 CLK_N.t0 272.06
R230 CLK_N.n0 CLK_N.t1 236.714
R231 CLK_N.n1 CLK_N.n0 76
R232 CLK_N CLK_N.n1 7.68
R233 CLK_N.n1 CLK_N 4.754
R234 a_1572_329.t1 a_1572_329.t0 236.868
R235 a_1714_47.n3 a_1714_47.n2 399.793
R236 a_1714_47.n1 a_1714_47.t4 241.535
R237 a_1714_47.n1 a_1714_47.t5 196.547
R238 a_1714_47.n2 a_1714_47.n0 183.436
R239 a_1714_47.n2 a_1714_47.n1 159.918
R240 a_1714_47.n0 a_1714_47.t2 70
R241 a_1714_47.n3 a_1714_47.t3 63.321
R242 a_1714_47.t0 a_1714_47.n3 63.321
R243 a_1714_47.n0 a_1714_47.t1 61.666
R244 a_1888_21.n5 a_1888_21.t4 387.206
R245 a_1888_21.n2 a_1888_21.t10 308.479
R246 a_1888_21.n7 a_1888_21.n6 301.911
R247 a_1888_21.n2 a_1888_21.t11 236.179
R248 a_1888_21.n4 a_1888_21.n2 235.764
R249 a_1888_21.n0 a_1888_21.t7 231.473
R250 a_1888_21.n1 a_1888_21.t8 221.719
R251 a_1888_21.n4 a_1888_21.n3 183.133
R252 a_1888_21.n0 a_1888_21.t6 163.994
R253 a_1888_21.n1 a_1888_21.t9 149.419
R254 a_1888_21.n1 a_1888_21.n0 144.6
R255 a_1888_21.n5 a_1888_21.t5 142.993
R256 a_1888_21.n6 a_1888_21.n5 128.841
R257 a_1888_21.n7 a_1888_21.t0 91.464
R258 a_1888_21.n2 a_1888_21.n1 85.688
R259 a_1888_21.t1 a_1888_21.n7 32.833
R260 a_1888_21.n6 a_1888_21.n4 30.494
R261 a_1888_21.n3 a_1888_21.t3 25.312
R262 a_1888_21.n3 a_1888_21.t2 25.312
R263 a_1823_47.t1 a_1823_47.t0 93.059
R264 VGND.n32 VGND.t6 188.008
R265 VGND.n62 VGND.t4 152.947
R266 VGND.n2 VGND.t8 114.327
R267 VGND.n42 VGND.n41 113.205
R268 VGND.n5 VGND.t12 110.749
R269 VGND.n21 VGND.n20 110.223
R270 VGND.n1 VGND.n0 108.988
R271 VGND.n67 VGND.n66 107.239
R272 VGND.n54 VGND.n53 106.463
R273 VGND.n41 VGND.t5 81.428
R274 VGND.n10 VGND.n9 64.275
R275 VGND.n53 VGND.t0 60
R276 VGND.n9 VGND.t1 57.796
R277 VGND.n0 VGND.t10 54.285
R278 VGND.n20 VGND.t9 41.428
R279 VGND.n20 VGND.t2 38.571
R280 VGND.n41 VGND.t3 38.571
R281 VGND.n53 VGND.t15 38.571
R282 VGND.n66 VGND.t13 38.571
R283 VGND.n66 VGND.t14 38.571
R284 VGND.n0 VGND.t7 25.934
R285 VGND.n9 VGND.t11 24.765
R286 VGND.n43 VGND.n42 16.564
R287 VGND.n22 VGND.n21 5.27
R288 VGND.n4 VGND.n3 4.65
R289 VGND.n6 VGND.n5 4.65
R290 VGND.n8 VGND.n7 4.65
R291 VGND.n11 VGND.n10 4.65
R292 VGND.n13 VGND.n12 4.65
R293 VGND.n15 VGND.n14 4.65
R294 VGND.n17 VGND.n16 4.65
R295 VGND.n19 VGND.n18 4.65
R296 VGND.n23 VGND.n22 4.65
R297 VGND.n25 VGND.n24 4.65
R298 VGND.n27 VGND.n26 4.65
R299 VGND.n29 VGND.n28 4.65
R300 VGND.n31 VGND.n30 4.65
R301 VGND.n34 VGND.n33 4.65
R302 VGND.n36 VGND.n35 4.65
R303 VGND.n38 VGND.n37 4.65
R304 VGND.n40 VGND.n39 4.65
R305 VGND.n44 VGND.n43 4.65
R306 VGND.n46 VGND.n45 4.65
R307 VGND.n48 VGND.n47 4.65
R308 VGND.n50 VGND.n49 4.65
R309 VGND.n52 VGND.n51 4.65
R310 VGND.n55 VGND.n54 4.65
R311 VGND.n57 VGND.n56 4.65
R312 VGND.n59 VGND.n58 4.65
R313 VGND.n61 VGND.n60 4.65
R314 VGND.n63 VGND.n62 4.65
R315 VGND.n65 VGND.n64 4.65
R316 VGND.n33 VGND.n32 4.141
R317 VGND.n68 VGND.n67 3.932
R318 VGND.n2 VGND.n1 3.73
R319 VGND.n4 VGND.n2 0.247
R320 VGND.n68 VGND.n65 0.137
R321 VGND VGND.n68 0.123
R322 VGND.n6 VGND.n4 0.119
R323 VGND.n8 VGND.n6 0.119
R324 VGND.n11 VGND.n8 0.119
R325 VGND.n13 VGND.n11 0.119
R326 VGND.n15 VGND.n13 0.119
R327 VGND.n17 VGND.n15 0.119
R328 VGND.n19 VGND.n17 0.119
R329 VGND.n23 VGND.n19 0.119
R330 VGND.n25 VGND.n23 0.119
R331 VGND.n27 VGND.n25 0.119
R332 VGND.n29 VGND.n27 0.119
R333 VGND.n31 VGND.n29 0.119
R334 VGND.n34 VGND.n31 0.119
R335 VGND.n36 VGND.n34 0.119
R336 VGND.n38 VGND.n36 0.119
R337 VGND.n40 VGND.n38 0.119
R338 VGND.n44 VGND.n40 0.119
R339 VGND.n46 VGND.n44 0.119
R340 VGND.n48 VGND.n46 0.119
R341 VGND.n50 VGND.n48 0.119
R342 VGND.n52 VGND.n50 0.119
R343 VGND.n55 VGND.n52 0.119
R344 VGND.n57 VGND.n55 0.119
R345 VGND.n59 VGND.n57 0.119
R346 VGND.n61 VGND.n59 0.119
R347 VGND.n63 VGND.n61 0.119
R348 VGND.n65 VGND.n63 0.119
R349 a_1041_47.t0 a_1041_47.t1 93.516
R350 a_1017_413.t0 a_1017_413.t1 211.071
R351 a_1800_413.t0 a_1800_413.t1 206.38
R352 a_2004_47.n0 a_2004_47.t2 274.441
R353 a_2004_47.n0 a_2004_47.t0 64.285
R354 a_2004_47.t1 a_2004_47.n0 49.151
R355 a_764_47.t0 a_764_47.t1 60
R356 a_2696_47.t0 a_2696_47.n2 237.868
R357 a_2696_47.n0 a_2696_47.t4 212.079
R358 a_2696_47.n1 a_2696_47.t5 212.079
R359 a_2696_47.n2 a_2696_47.t1 150.778
R360 a_2696_47.n0 a_2696_47.t3 139.779
R361 a_2696_47.n1 a_2696_47.t2 139.779
R362 a_2696_47.n2 a_2696_47.n1 111.493
R363 a_2696_47.n1 a_2696_47.n0 61.345
R364 Q.n3 Q.n2 142.894
R365 Q.n1 Q.n0 92.5
R366 Q Q.n1 69.688
R367 Q.n2 Q.t1 26.595
R368 Q.n2 Q.t0 26.595
R369 Q.n0 Q.t2 24.923
R370 Q.n0 Q.t3 24.923
R371 Q.n3 Q 9.375
R372 Q Q.n3 7.629
R373 Q.n1 Q 6.912
R374 a_193_47.n0 a_193_47.t5 534.467
R375 a_193_47.n1 a_193_47.t2 236.795
R376 a_193_47.n1 a_193_47.t4 231.324
R377 a_193_47.n3 a_193_47.t1 210.124
R378 a_193_47.n0 a_193_47.t3 137.933
R379 a_193_47.t0 a_193_47.n3 121.825
R380 a_193_47.n2 a_193_47.n0 12.947
R381 a_193_47.n3 a_193_47.n2 4.716
R382 a_193_47.n2 a_193_47.n1 4.65
R383 D.n0 D.t0 308.479
R384 D.n0 D.t1 224.932
R385 D.n1 D.n0 76
R386 D.n1 D 40.64
R387 D D.n1 2.88
R388 Q_N.n3 Q_N.n2 142.77
R389 Q_N.n1 Q_N.n0 92.5
R390 Q_N Q_N.n1 85.278
R391 Q_N.n2 Q_N.t1 26.595
R392 Q_N.n2 Q_N.t0 26.595
R393 Q_N.n0 Q_N.t3 24.923
R394 Q_N.n0 Q_N.t2 24.923
R395 Q_N.n3 Q_N 9.243
R396 Q_N Q_N.n3 7.748
R397 Q_N.n1 Q_N 6.4
R398 a_381_47.t0 a_381_47.t1 60
R399 a_1619_47.n1 a_1619_47.n0 67.2
R400 a_1619_47.n0 a_1619_47.t1 66.666
R401 a_1619_47.n0 a_1619_47.t0 13.143
R402 a_752_413.t0 a_752_413.t1 126.642
R403 RESET_B.n0 RESET_B.t1 201.872
R404 RESET_B.n0 RESET_B.t0 172.951
R405 RESET_B RESET_B.n0 78
C0 SET_B VGND 0.36fF
C1 VPB VPWR 0.32fF
C2 VPWR Q 0.30fF
C3 VGND Q_N 0.22fF
C4 VPWR VGND 0.19fF
C5 VGND Q 0.15fF
C6 SCD SCE 0.11fF
C7 VPWR Q_N 0.23fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__sdfbbp_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__sdfbbp_1 SCD SCE RESET_B VGND CLK SET_B Q VPWR D Q_N VNB
+ VPB
X0 a_381_363.t1 SCD.t0 VPWR.t11 VPB.t17 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1 a_1107_21.t3 SET_B.t0 VPWR.t2 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 VPWR.t12 a_1400_21.t2 a_2122_329.t0 VPB.t19 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X3 Q.t1 a_2596_47.t2 VPWR.t6 VPB.t8 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 a_931_47.t2 a_193_47.t2 a_453_363.t5 VPB.t9 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 VPWR.t13 a_1400_21.t3 a_1351_329.t0 VPB.t20 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X6 a_1251_47.t0 a_1400_21.t4 a_1107_21.t2 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X7 VPWR.t0 SCE.t0 a_423_315.t1 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 a_1351_329.t1 a_931_47.t4 a_1107_21.t0 VPB.t18 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X9 VPWR.t7 RESET_B.t0 a_1400_21.t1 VPB.t11 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X10 VPWR.t4 CLK.t0 a_27_47.t0 VPB.t6 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X11 a_1572_329.t0 a_1107_21.t4 VPWR.t14 VPB.t21 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X12 a_2122_329.t1 a_1714_47.t4 a_1887_21.t2 VPB.t5 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X13 a_2026_47.t2 SET_B.t1 VGND.t12 VNB.t21 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14 a_1041_47.t1 a_193_47.t3 a_931_47.t1 VNB.t17 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X15 VGND.t1 a_1887_21.t4 a_1822_47.t0 VNB.t9 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16 VPWR.t15 a_1107_21.t5 a_1017_413.t0 VPB.t22 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17 a_1107_21.t1 a_931_47.t5 a_1251_47.t1 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X18 VPWR.t9 a_1887_21.t5 a_1800_413.t0 VPB.t13 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19 a_764_47.t0 a_423_315.t2 VGND.t6 VNB.t12 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20 a_1887_21.t1 a_1714_47.t5 a_2026_47.t1 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X21 a_1887_21.t3 SET_B.t2 VPWR.t3 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22 a_931_47.t0 a_27_47.t2 a_453_363.t2 VNB.t10 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X23 a_1800_413.t1 a_193_47.t4 a_1714_47.t2 VPB.t10 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24 a_193_47.t1 a_27_47.t3 VGND.t9 VNB.t11 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X25 a_453_363.t4 D.t0 a_764_47.t1 VNB.t13 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X26 VGND.t8 SCE.t1 a_423_315.t0 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X27 a_1714_47.t0 a_27_47.t4 a_1572_329.t1 VPB.t14 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X28 VGND.t4 a_1107_21.t6 a_1041_47.t0 VNB.t5 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X29 a_2026_47.t0 a_1400_21.t5 a_1887_21.t0 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X30 Q.t0 a_2596_47.t3 VGND.t11 VNB.t18 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X31 VGND.t3 a_1887_21.t6 a_2596_47.t0 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X32 a_193_47.t0 a_27_47.t5 VPWR.t10 VPB.t15 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X33 a_1017_413.t1 a_27_47.t6 a_931_47.t3 VPB.t23 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X34 a_453_363.t1 SCE.t2 a_381_47.t1 VNB.t7 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X35 VPWR.t8 a_1887_21.t7 a_2596_47.t1 VPB.t12 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X36 a_453_363.t3 a_423_315.t3 a_381_363.t0 VPB.t16 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X37 a_381_47.t0 SCD.t1 VGND.t7 VNB.t14 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X38 a_1714_47.t3 a_193_47.t5 a_1618_47.t1 VNB.t16 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X39 a_1822_47.t1 a_27_47.t7 a_1714_47.t1 VNB.t19 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X40 Q_N.t0 a_1887_21.t8 VGND.t2 VNB.t8 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X41 Q_N.t1 a_1887_21.t9 VPWR.t1 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X42 a_453_363.t0 D.t1 a_752_413.t0 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X43 a_1251_47.t2 SET_B.t3 VGND.t13 VNB.t20 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X44 a_1618_47.t0 a_1107_21.t7 VGND.t5 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X45 a_752_413.t1 SCE.t3 VPWR.t5 VPB.t7 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X46 VGND.t0 CLK.t1 a_27_47.t1 VNB.t15 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X47 VGND.t10 RESET_B.t1 a_1400_21.t0 VNB.t6 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
R0 SCD.n0 SCD.t1 302.41
R1 SCD.n0 SCD.t0 173.876
R2 SCD SCD.n0 78.057
R3 VPWR.n6 VPWR.t12 500.865
R4 VPWR.n1 VPWR.n0 440.25
R5 VPWR.n60 VPWR.n59 311.893
R6 VPWR.n47 VPWR.n46 308.79
R7 VPWR.n36 VPWR.n35 306.984
R8 VPWR.n14 VPWR.n13 292.5
R9 VPWR.n55 VPWR.t11 229.845
R10 VPWR.n3 VPWR.n2 172.733
R11 VPWR.n28 VPWR.n27 164.214
R12 VPWR.n13 VPWR.t3 91.464
R13 VPWR.n13 VPWR.t9 91.464
R14 VPWR.n35 VPWR.t2 91.464
R15 VPWR.n27 VPWR.t14 86.773
R16 VPWR.n35 VPWR.t15 86.773
R17 VPWR.n46 VPWR.t5 63.321
R18 VPWR.n46 VPWR.t0 63.321
R19 VPWR.n0 VPWR.t7 63.101
R20 VPWR.n2 VPWR.t8 58.484
R21 VPWR.n59 VPWR.t10 41.554
R22 VPWR.n59 VPWR.t4 41.554
R23 VPWR.n27 VPWR.t13 38.696
R24 VPWR.n2 VPWR.t6 31.83
R25 VPWR.n0 VPWR.t1 28.032
R26 VPWR.n5 VPWR.n4 4.65
R27 VPWR.n8 VPWR.n7 4.65
R28 VPWR.n10 VPWR.n9 4.65
R29 VPWR.n12 VPWR.n11 4.65
R30 VPWR.n16 VPWR.n15 4.65
R31 VPWR.n18 VPWR.n17 4.65
R32 VPWR.n20 VPWR.n19 4.65
R33 VPWR.n22 VPWR.n21 4.65
R34 VPWR.n24 VPWR.n23 4.65
R35 VPWR.n26 VPWR.n25 4.65
R36 VPWR.n30 VPWR.n29 4.65
R37 VPWR.n32 VPWR.n31 4.65
R38 VPWR.n34 VPWR.n33 4.65
R39 VPWR.n37 VPWR.n36 4.65
R40 VPWR.n39 VPWR.n38 4.65
R41 VPWR.n41 VPWR.n40 4.65
R42 VPWR.n43 VPWR.n42 4.65
R43 VPWR.n45 VPWR.n44 4.65
R44 VPWR.n48 VPWR.n47 4.65
R45 VPWR.n50 VPWR.n49 4.65
R46 VPWR.n52 VPWR.n51 4.65
R47 VPWR.n54 VPWR.n53 4.65
R48 VPWR.n56 VPWR.n55 4.65
R49 VPWR.n58 VPWR.n57 4.65
R50 VPWR.n3 VPWR.n1 4.611
R51 VPWR.n61 VPWR.n60 3.932
R52 VPWR.n7 VPWR.n6 3.84
R53 VPWR.n29 VPWR.n28 3.388
R54 VPWR.n15 VPWR.n14 2.443
R55 VPWR.n5 VPWR.n3 0.144
R56 VPWR.n61 VPWR.n58 0.137
R57 VPWR VPWR.n61 0.123
R58 VPWR.n8 VPWR.n5 0.119
R59 VPWR.n10 VPWR.n8 0.119
R60 VPWR.n12 VPWR.n10 0.119
R61 VPWR.n16 VPWR.n12 0.119
R62 VPWR.n18 VPWR.n16 0.119
R63 VPWR.n20 VPWR.n18 0.119
R64 VPWR.n22 VPWR.n20 0.119
R65 VPWR.n24 VPWR.n22 0.119
R66 VPWR.n26 VPWR.n24 0.119
R67 VPWR.n30 VPWR.n26 0.119
R68 VPWR.n32 VPWR.n30 0.119
R69 VPWR.n34 VPWR.n32 0.119
R70 VPWR.n37 VPWR.n34 0.119
R71 VPWR.n39 VPWR.n37 0.119
R72 VPWR.n41 VPWR.n39 0.119
R73 VPWR.n43 VPWR.n41 0.119
R74 VPWR.n45 VPWR.n43 0.119
R75 VPWR.n48 VPWR.n45 0.119
R76 VPWR.n50 VPWR.n48 0.119
R77 VPWR.n52 VPWR.n50 0.119
R78 VPWR.n54 VPWR.n52 0.119
R79 VPWR.n56 VPWR.n54 0.119
R80 VPWR.n58 VPWR.n56 0.119
R81 a_381_363.t0 a_381_363.t1 64.64
R82 VPB.t16 VPB.t0 636.292
R83 VPB.t19 VPB.t11 588.94
R84 VPB.t2 VPB.t12 556.386
R85 VPB.t15 VPB.t17 556.386
R86 VPB.t21 VPB.t14 426.168
R87 VPB.t20 VPB.t21 405.451
R88 VPB.t23 VPB.t22 355.14
R89 VPB.t10 VPB.t13 349.221
R90 VPB.t13 VPB.t4 319.626
R91 VPB.t3 VPB.t18 319.626
R92 VPB.t22 VPB.t3 313.707
R93 VPB.t11 VPB.t2 287.071
R94 VPB.t1 VPB.t9 287.071
R95 VPB.t4 VPB.t5 284.112
R96 VPB.t12 VPB.t8 281.152
R97 VPB.t14 VPB.t10 248.598
R98 VPB.t18 VPB.t20 248.598
R99 VPB.t9 VPB.t23 248.598
R100 VPB.t7 VPB.t1 248.598
R101 VPB.t0 VPB.t7 248.598
R102 VPB.t6 VPB.t15 248.598
R103 VPB.t5 VPB.t19 213.084
R104 VPB.t17 VPB.t16 213.084
R105 VPB VPB.t6 142.056
R106 SET_B.n0 SET_B.t0 396.831
R107 SET_B.n3 SET_B.t2 393.971
R108 SET_B.n3 SET_B.t1 134.267
R109 SET_B.n0 SET_B.t3 134.063
R110 SET_B SET_B.n6 13.6
R111 SET_B.n5 SET_B.n3 13.016
R112 SET_B.n1 SET_B.n0 6.985
R113 SET_B.n6 SET_B.n5 6.318
R114 SET_B.n6 SET_B.n1 2.521
R115 SET_B.n2 SET_B 2.521
R116 SET_B.n6 SET_B.n2 0.775
R117 SET_B.n5 SET_B.n4 0.001
R118 a_1107_21.n5 a_1107_21.t6 387.959
R119 a_1107_21.n2 a_1107_21.t4 299.91
R120 a_1107_21.n7 a_1107_21.n6 292.5
R121 a_1107_21.n2 a_1107_21.t7 167.627
R122 a_1107_21.n5 a_1107_21.t5 143.746
R123 a_1107_21.n4 a_1107_21.n2 140.193
R124 a_1107_21.n6 a_1107_21.n5 114.656
R125 a_1107_21.n4 a_1107_21.n3 110.36
R126 a_1107_21.n0 a_1107_21.t3 110.226
R127 a_1107_21.n6 a_1107_21.n4 81.287
R128 a_1107_21.t0 a_1107_21.n1 63.321
R129 a_1107_21.t0 a_1107_21.n7 63.321
R130 a_1107_21.n3 a_1107_21.t2 25.312
R131 a_1107_21.n3 a_1107_21.t1 25.312
R132 a_1107_21.n1 a_1107_21.n0 9.38
R133 a_1400_21.t1 a_1400_21.n3 448.039
R134 a_1400_21.n1 a_1400_21.t5 211.511
R135 a_1400_21.n1 a_1400_21.t2 206.934
R136 a_1400_21.n0 a_1400_21.t3 204.868
R137 a_1400_21.n0 a_1400_21.t4 204.408
R138 a_1400_21.n2 a_1400_21.t0 195.463
R139 a_1400_21.n3 a_1400_21.n0 126.544
R140 a_1400_21.n2 a_1400_21.n1 76
R141 a_1400_21.n3 a_1400_21.n2 9.774
R142 a_2122_329.t0 a_2122_329.t1 49.25
R143 a_2596_47.n0 a_2596_47.t2 238.589
R144 a_2596_47.t1 a_2596_47.n1 237.868
R145 a_2596_47.n0 a_2596_47.t3 166.289
R146 a_2596_47.n1 a_2596_47.t0 150.778
R147 a_2596_47.n1 a_2596_47.n0 99.078
R148 Q.n1 Q.t1 207.372
R149 Q.n0 Q.t0 117.423
R150 Q Q.n0 69.449
R151 Q.n1 Q 9.019
R152 Q Q.n1 7.458
R153 Q.n0 Q 6.646
R154 a_193_47.n1 a_193_47.t2 538.597
R155 a_193_47.t0 a_193_47.n3 278.596
R156 a_193_47.n0 a_193_47.t4 267.397
R157 a_193_47.n0 a_193_47.t5 207.657
R158 a_193_47.n3 a_193_47.t1 150.413
R159 a_193_47.n1 a_193_47.t3 135.786
R160 a_193_47.n2 a_193_47.n1 10.203
R161 a_193_47.n3 a_193_47.n2 8.238
R162 a_193_47.n2 a_193_47.n0 7.5
R163 a_453_363.n2 a_453_363.n0 355.646
R164 a_453_363.t3 a_453_363.n3 258.131
R165 a_453_363.n3 a_453_363.t1 177.756
R166 a_453_363.n2 a_453_363.n1 133.46
R167 a_453_363.n0 a_453_363.t5 93.809
R168 a_453_363.n1 a_453_363.t2 63.333
R169 a_453_363.n0 a_453_363.t0 63.321
R170 a_453_363.n1 a_453_363.t4 29.726
R171 a_453_363.n3 a_453_363.n2 24.553
R172 a_931_47.n3 a_931_47.n2 415.031
R173 a_931_47.n1 a_931_47.t5 216.899
R174 a_931_47.n1 a_931_47.t4 210.473
R175 a_931_47.n2 a_931_47.n0 196.424
R176 a_931_47.n2 a_931_47.n1 140.828
R177 a_931_47.n0 a_931_47.t0 70
R178 a_931_47.n0 a_931_47.t1 63.333
R179 a_931_47.n3 a_931_47.t3 63.321
R180 a_931_47.t2 a_931_47.n3 63.321
R181 a_1351_329.t0 a_1351_329.t1 63.321
R182 a_1251_47.t0 a_1251_47.n0 282.717
R183 a_1251_47.n0 a_1251_47.t1 42.008
R184 a_1251_47.n0 a_1251_47.t2 38.571
R185 VNB.t7 VNB.t0 6664.71
R186 VNB.t11 VNB.t14 6082.35
R187 VNB.t2 VNB.t6 4595.56
R188 VNB.t8 VNB.t4 4545.05
R189 VNB VNB.t15 4270.59
R190 VNB.t5 VNB.t20 3688.24
R191 VNB.t10 VNB.t17 3558.82
R192 VNB.t9 VNB.t21 3526.47
R193 VNB.t16 VNB.t19 3494.12
R194 VNB.t0 VNB.t12 3202.94
R195 VNB.t17 VNB.t5 3105.88
R196 VNB.t19 VNB.t9 3073.53
R197 VNB.t13 VNB.t10 3073.53
R198 VNB.t15 VNB.t11 2717.65
R199 VNB.t14 VNB.t7 2523.53
R200 VNB.t12 VNB.t13 2329.41
R201 VNB.t6 VNB.t8 2296.97
R202 VNB.t4 VNB.t18 2296.7
R203 VNB.t21 VNB.t1 2280.14
R204 VNB.t1 VNB.t2 2053.33
R205 VNB.t20 VNB.t3 213.215
R206 VNB.t20 VNB.t16 42.773
R207 SCE.n1 SCE.n0 310.086
R208 SCE.n2 SCE.n1 296.028
R209 SCE.n0 SCE.t3 228.146
R210 SCE.n2 SCE.t2 97.202
R211 SCE.n0 SCE.t0 93.186
R212 SCE.n1 SCE.t1 93.186
R213 SCE.n3 SCE.n2 81.27
R214 SCE SCE.n3 29.381
R215 SCE.n3 SCE 10.181
R216 a_423_315.n0 a_423_315.t1 427.341
R217 a_423_315.n0 a_423_315.t3 391.928
R218 a_423_315.n1 a_423_315.t2 209.832
R219 a_423_315.t0 a_423_315.n1 189.347
R220 a_423_315.n1 a_423_315.n0 89.034
R221 RESET_B.n0 RESET_B.t1 203.042
R222 RESET_B.n0 RESET_B.t0 174.121
R223 RESET_B RESET_B.n0 78.109
R224 CLK.n0 CLK.t0 272.06
R225 CLK.n0 CLK.t1 236.714
R226 CLK.n1 CLK.n0 76
R227 CLK CLK.n1 7.68
R228 CLK.n1 CLK 4.754
R229 a_27_47.n0 a_27_47.t7 532.86
R230 a_27_47.n3 a_27_47.t5 262.942
R231 a_27_47.t0 a_27_47.n5 242.769
R232 a_27_47.n1 a_27_47.t2 236.795
R233 a_27_47.n1 a_27_47.t6 231.324
R234 a_27_47.n3 a_27_47.t3 227.596
R235 a_27_47.n4 a_27_47.t1 194.667
R236 a_27_47.n0 a_27_47.t4 137.933
R237 a_27_47.n4 a_27_47.n3 76
R238 a_27_47.n5 a_27_47.n4 35.339
R239 a_27_47.n2 a_27_47.n0 12.947
R240 a_27_47.n5 a_27_47.n2 8.243
R241 a_27_47.n2 a_27_47.n1 4.65
R242 a_1572_329.t0 a_1572_329.t1 236.868
R243 a_1714_47.n3 a_1714_47.n2 399.793
R244 a_1714_47.n1 a_1714_47.t4 241.535
R245 a_1714_47.n1 a_1714_47.t5 196.547
R246 a_1714_47.n2 a_1714_47.n0 183.436
R247 a_1714_47.n2 a_1714_47.n1 159.918
R248 a_1714_47.n0 a_1714_47.t3 70
R249 a_1714_47.n3 a_1714_47.t2 63.321
R250 a_1714_47.t0 a_1714_47.n3 63.321
R251 a_1714_47.n0 a_1714_47.t1 60
R252 a_1887_21.n4 a_1887_21.t4 386.846
R253 a_1887_21.n6 a_1887_21.n5 301.911
R254 a_1887_21.n1 a_1887_21.t9 268.312
R255 a_1887_21.n0 a_1887_21.t7 231.942
R256 a_1887_21.n3 a_1887_21.n1 229.286
R257 a_1887_21.n1 a_1887_21.t8 196.012
R258 a_1887_21.n3 a_1887_21.n2 185.391
R259 a_1887_21.n0 a_1887_21.t6 164.463
R260 a_1887_21.n1 a_1887_21.n0 151.74
R261 a_1887_21.n4 a_1887_21.t5 142.633
R262 a_1887_21.n5 a_1887_21.n4 128.841
R263 a_1887_21.n6 a_1887_21.t3 91.464
R264 a_1887_21.t2 a_1887_21.n6 32.833
R265 a_1887_21.n5 a_1887_21.n3 30.494
R266 a_1887_21.n2 a_1887_21.t0 25.312
R267 a_1887_21.n2 a_1887_21.t1 25.312
R268 VGND.n24 VGND.t5 187.788
R269 VGND.n54 VGND.t7 155.135
R270 VGND.n34 VGND.n33 113.205
R271 VGND.n3 VGND.n0 113.067
R272 VGND.n13 VGND.n12 110.223
R273 VGND.n59 VGND.n58 107.239
R274 VGND.n46 VGND.n45 106.463
R275 VGND.n33 VGND.t4 81.428
R276 VGND.n12 VGND.t12 70
R277 VGND.n2 VGND.n1 64.275
R278 VGND.n45 VGND.t8 60
R279 VGND.n1 VGND.t10 57.796
R280 VGND.n0 VGND.t3 54.285
R281 VGND.n12 VGND.t1 42.857
R282 VGND.n33 VGND.t13 38.571
R283 VGND.n45 VGND.t6 38.571
R284 VGND.n58 VGND.t9 38.571
R285 VGND.n58 VGND.t0 38.571
R286 VGND.n0 VGND.t11 25.934
R287 VGND.n1 VGND.t2 24.765
R288 VGND.n35 VGND.n34 16.564
R289 VGND.n14 VGND.n13 5.27
R290 VGND.n5 VGND.n4 4.65
R291 VGND.n7 VGND.n6 4.65
R292 VGND.n9 VGND.n8 4.65
R293 VGND.n11 VGND.n10 4.65
R294 VGND.n15 VGND.n14 4.65
R295 VGND.n17 VGND.n16 4.65
R296 VGND.n19 VGND.n18 4.65
R297 VGND.n21 VGND.n20 4.65
R298 VGND.n23 VGND.n22 4.65
R299 VGND.n26 VGND.n25 4.65
R300 VGND.n28 VGND.n27 4.65
R301 VGND.n30 VGND.n29 4.65
R302 VGND.n32 VGND.n31 4.65
R303 VGND.n36 VGND.n35 4.65
R304 VGND.n38 VGND.n37 4.65
R305 VGND.n40 VGND.n39 4.65
R306 VGND.n42 VGND.n41 4.65
R307 VGND.n44 VGND.n43 4.65
R308 VGND.n47 VGND.n46 4.65
R309 VGND.n49 VGND.n48 4.65
R310 VGND.n51 VGND.n50 4.65
R311 VGND.n53 VGND.n52 4.65
R312 VGND.n55 VGND.n54 4.65
R313 VGND.n57 VGND.n56 4.65
R314 VGND.n3 VGND.n2 3.969
R315 VGND.n60 VGND.n59 3.932
R316 VGND.n25 VGND.n24 3.764
R317 VGND.n5 VGND.n3 0.146
R318 VGND.n60 VGND.n57 0.137
R319 VGND VGND.n60 0.123
R320 VGND.n7 VGND.n5 0.119
R321 VGND.n9 VGND.n7 0.119
R322 VGND.n11 VGND.n9 0.119
R323 VGND.n15 VGND.n11 0.119
R324 VGND.n17 VGND.n15 0.119
R325 VGND.n19 VGND.n17 0.119
R326 VGND.n21 VGND.n19 0.119
R327 VGND.n23 VGND.n21 0.119
R328 VGND.n26 VGND.n23 0.119
R329 VGND.n28 VGND.n26 0.119
R330 VGND.n30 VGND.n28 0.119
R331 VGND.n32 VGND.n30 0.119
R332 VGND.n36 VGND.n32 0.119
R333 VGND.n38 VGND.n36 0.119
R334 VGND.n40 VGND.n38 0.119
R335 VGND.n42 VGND.n40 0.119
R336 VGND.n44 VGND.n42 0.119
R337 VGND.n47 VGND.n44 0.119
R338 VGND.n49 VGND.n47 0.119
R339 VGND.n51 VGND.n49 0.119
R340 VGND.n53 VGND.n51 0.119
R341 VGND.n55 VGND.n53 0.119
R342 VGND.n57 VGND.n55 0.119
R343 a_2026_47.t0 a_2026_47.n0 272.229
R344 a_2026_47.n0 a_2026_47.t1 42.008
R345 a_2026_47.n0 a_2026_47.t2 38.571
R346 a_1041_47.t0 a_1041_47.t1 93.516
R347 a_1822_47.t0 a_1822_47.t1 93.059
R348 a_1017_413.t0 a_1017_413.t1 211.071
R349 a_1800_413.t0 a_1800_413.t1 206.38
R350 a_764_47.t0 a_764_47.t1 60
R351 D.n0 D.t0 308.479
R352 D.n0 D.t1 224.932
R353 D.n1 D.n0 76
R354 D.n1 D 40.64
R355 D D.n1 2.88
R356 a_381_47.t0 a_381_47.t1 68.571
R357 a_1618_47.n0 a_1618_47.t1 68.333
R358 a_1618_47.n1 a_1618_47.n0 67.2
R359 a_1618_47.n0 a_1618_47.t0 13.143
R360 Q_N.n1 Q_N.t1 207.566
R361 Q_N.n0 Q_N.t0 117.423
R362 Q_N Q_N.n0 79.437
R363 Q_N.n1 Q_N 8.185
R364 Q_N Q_N.n1 6.859
R365 Q_N.n0 Q_N 5.614
R366 a_752_413.t0 a_752_413.t1 126.642
C0 SCD SCE 0.11fF
C1 SET_B VGND 0.36fF
C2 VPB VPWR 0.30fF
C3 VGND Q_N 0.12fF
C4 VPWR Q 0.14fF
C5 VPWR VGND 0.14fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__sdfrbp_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__sdfrbp_1 VPWR VGND Q_N SCE SCD D RESET_B CLK Q VNB VPB
X0 a_193_47.t0 a_27_47.t2 VPWR.t12 VPB.t16 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_780_389.t1 a_299_66.t2 a_620_389.t1 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=540000u l=150000u
X2 VGND.t4 a_1767_21.t3 a_2324_47.t1 VNB sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X3 a_1245_303.t1 a_1079_413.t4 VPWR.t11 VPB.t13 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X4 VPWR.t7 a_1592_47.t4 a_1767_21.t1 VPB.t8 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 VGND.t5 a_1767_21.t4 a_1701_47.t0 VNB sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 a_1758_413.t1 a_193_47.t2 a_1592_47.t2 VPB.t18 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7 VPWR.t13 a_1767_21.t5 a_2324_47.t0 VPB.t19 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X8 a_1767_21.t2 a_1592_47.t5 a_1946_47.t1 VNB sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9 VGND.t11 SCD.t0 a_817_66.t1 VNB sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=180000u
X10 a_538_389.t1 SCE.t0 VPWR.t9 VPB.t11 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=540000u l=150000u
X11 VPWR.t4 SCD.t1 a_780_389.t0 VPB.t5 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=540000u l=150000u
X12 VPWR.t8 SCE.t1 a_299_66.t0 VPB.t9 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=540000u l=150000u
X13 a_1767_21.t0 RESET_B.t0 VPWR.t5 VPB.t6 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14 a_193_47.t1 a_27_47.t3 VGND.t8 VNB sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X15 a_620_389.t2 D.t0 a_569_119.t0 VNB sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16 a_1187_47.t0 a_193_47.t3 a_1079_413.t2 VNB sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X17 a_1293_47.t0 a_1245_303.t4 a_1187_47.t1 VNB sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18 VPWR.t10 a_1245_303.t5 a_1191_413.t1 VPB.t12 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19 a_620_389.t3 D.t1 a_538_389.t0 VPB.t10 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=540000u l=150000u
X20 a_1191_413.t0 a_27_47.t4 a_1079_413.t0 VPB.t15 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21 a_569_119.t1 a_299_66.t3 VGND.t6 VNB sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22 VPWR.t2 a_1767_21.t6 a_1758_413.t0 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23 VGND.t0 RESET_B.t1 a_1293_47.t1 VNB sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24 Q.t1 a_1767_21.t7 VPWR.t3 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X25 Q.t0 a_1767_21.t8 VGND.t3 VNB sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X26 Q_N.t0 a_2324_47.t2 VGND.t2 VNB sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X27 a_1079_413.t1 a_27_47.t5 a_620_389.t4 VNB sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X28 a_1191_413.t2 RESET_B.t2 VPWR.t6 VPB.t7 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X29 a_1701_47.t1 a_27_47.t6 a_1592_47.t0 VNB sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X30 a_1946_47.t0 RESET_B.t3 VGND.t1 VNB sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X31 Q_N.t1 a_2324_47.t3 VPWR.t1 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X32 a_1592_47.t3 a_193_47.t4 a_1245_303.t3 VNB sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X33 VGND.t10 SCE.t2 a_299_66.t1 VNB sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X34 a_1592_47.t1 a_27_47.t7 a_1245_303.t2 VPB.t14 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X35 a_1245_303.t0 a_1079_413.t5 VGND.t7 VNB sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X36 a_1079_413.t3 a_193_47.t5 a_620_389.t5 VPB.t17 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X37 VPWR.t0 CLK.t0 a_27_47.t0 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X38 a_817_66.t0 SCE.t3 a_620_389.t0 VNB sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=500000u
X39 VGND.t9 CLK.t1 a_27_47.t1 VNB sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
R0 a_27_47.n1 a_27_47.t4 534.047
R1 a_27_47.n0 a_27_47.t7 489.903
R2 a_27_47.n1 a_27_47.t5 276.816
R3 a_27_47.t0 a_27_47.n9 243.743
R4 a_27_47.n7 a_27_47.t2 238.856
R5 a_27_47.n0 a_27_47.t6 204.42
R6 a_27_47.n3 a_27_47.t1 175.866
R7 a_27_47.n5 a_27_47.t3 156.738
R8 a_27_47.n2 a_27_47.n0 14.808
R9 a_27_47.n6 a_27_47.n5 12.496
R10 a_27_47.n2 a_27_47.n1 11.633
R11 a_27_47.n8 a_27_47.n7 9.3
R12 a_27_47.n9 a_27_47.n2 6.029
R13 a_27_47.n4 a_27_47.n3 2.844
R14 a_27_47.n7 a_27_47.n6 2.677
R15 a_27_47.n9 a_27_47.n8 1.13
R16 a_27_47.n8 a_27_47.n4 0.609
R17 VPWR.n4 VPWR.t11 514.01
R18 VPWR.n5 VPWR.t4 408.48
R19 VPWR.n1 VPWR.t7 370.56
R20 VPWR.n16 VPWR.n15 323.37
R21 VPWR.n7 VPWR.n6 311.893
R22 VPWR.n3 VPWR.n2 310.932
R23 VPWR.n35 VPWR.n34 292.5
R24 VPWR.n55 VPWR.n54 168.669
R25 VPWR.n0 VPWR.t3 152.716
R26 VPWR.n2 VPWR.t2 114.916
R27 VPWR.n34 VPWR.t6 103.19
R28 VPWR.n34 VPWR.t10 93.809
R29 VPWR.n2 VPWR.t5 63.321
R30 VPWR.n15 VPWR.t9 49.25
R31 VPWR.n15 VPWR.t8 49.25
R32 VPWR.n54 VPWR.t1 36.158
R33 VPWR.n54 VPWR.t13 36.158
R34 VPWR.n6 VPWR.t0 29.55
R35 VPWR.n6 VPWR.t12 26.595
R36  VPWR.n55 10.815
R37 VPWR.n17 VPWR.n16 9.411
R38 VPWR.n53 VPWR.n52 4.65
R39 VPWR.n51 VPWR.n0 4.65
R40 VPWR.n50 VPWR.n1 4.65
R41 VPWR.n49 VPWR.n48 4.65
R42 VPWR.n47 VPWR.n3 4.65
R43 VPWR.n46 VPWR.n45 4.65
R44 VPWR.n44 VPWR.n43 4.65
R45 VPWR.n42 VPWR.n41 4.65
R46 VPWR.n40 VPWR.n4 4.65
R47 VPWR.n39 VPWR.n38 4.65
R48 VPWR.n37 VPWR.n36 4.65
R49 VPWR.n33 VPWR.n32 4.65
R50 VPWR.n31 VPWR.n30 4.65
R51 VPWR.n29 VPWR.n28 4.65
R52 VPWR.n27 VPWR.n26 4.65
R53 VPWR.n25 VPWR.n5 4.65
R54 VPWR.n24 VPWR.n23 4.65
R55 VPWR.n22 VPWR.n21 4.65
R56 VPWR.n20 VPWR.n19 4.65
R57 VPWR.n18 VPWR.n17 4.65
R58 VPWR.n14 VPWR.n13 4.65
R59 VPWR.n12 VPWR.n11 4.65
R60 VPWR.n10 VPWR.n9 4.65
R61 VPWR.n8 VPWR.n7 3.958
R62 VPWR.n36 VPWR.n35 2.702
R63 VPWR.n55 VPWR.n53 0.76
R64 VPWR.n10 VPWR.n8 0.137
R65 VPWR.n8 VPWR 0.121
R66 VPWR.n53 VPWR.n51 0.119
R67 VPWR.n51 VPWR.n50 0.119
R68 VPWR.n50 VPWR.n49 0.119
R69 VPWR.n49 VPWR.n47 0.119
R70 VPWR.n47 VPWR.n46 0.119
R71 VPWR.n46 VPWR.n44 0.119
R72 VPWR.n44 VPWR.n42 0.119
R73 VPWR.n42 VPWR.n40 0.119
R74 VPWR.n40 VPWR.n39 0.119
R75 VPWR.n39 VPWR.n37 0.119
R76 VPWR.n37 VPWR.n33 0.119
R77 VPWR.n33 VPWR.n31 0.119
R78 VPWR.n31 VPWR.n29 0.119
R79 VPWR.n29 VPWR.n27 0.119
R80 VPWR.n27 VPWR.n25 0.119
R81 VPWR.n25 VPWR.n24 0.119
R82 VPWR.n24 VPWR.n22 0.119
R83 VPWR.n22 VPWR.n20 0.119
R84 VPWR.n20 VPWR.n18 0.119
R85 VPWR.n18 VPWR.n14 0.119
R86 VPWR.n14 VPWR.n12 0.119
R87 VPWR.n12 VPWR.n10 0.119
R88 a_193_47.n1 a_193_47.t4 266.53
R89 a_193_47.n0 a_193_47.t3 265.71
R90 a_193_47.n1 a_193_47.t2 231.814
R91 a_193_47.n3 a_193_47.t1 210.139
R92 a_193_47.n0 a_193_47.t5 146.401
R93 a_193_47.t0 a_193_47.n3 38.199
R94 a_193_47.n2 a_193_47.n1 7.332
R95 a_193_47.n3 a_193_47.n2 6.062
R96 a_193_47.n2 a_193_47.n0 3.302
R97 VPB.t16 VPB.t9 774.312
R98 VPB.t5 VPB.t17 637.547
R99 VPB.t8 VPB.t4 556.386
R100 VPB.t7 VPB.t13 556.386
R101 VPB.t10 VPB.t0 511.784
R102 VPB.t4 VPB 414.33
R103 VPB.t12 VPB.t7 337.383
R104 VPB.t17 VPB.t15 331.464
R105 VPB.t3 VPB.t6 313.707
R106 VPB.t13 VPB.t14 281.152
R107 VPB.t0 VPB.t5 275.084
R108 VPB.t9 VPB.t11 268.686
R109 VPB.t11 VPB.t10 262.289
R110 VPB.t19 VPB.t2 260.436
R111 VPB.t1 VPB.t16 257.476
R112 VPB.t14 VPB.t18 254.517
R113 VPB.t6 VPB.t8 248.598
R114 VPB.t15 VPB.t12 248.598
R115 VPB.t18 VPB.t3 242.679
R116 VPB VPB.t1 177.57
R117 VPB VPB.t19 142.056
R118 a_299_66.n0 a_299_66.t2 1032.99
R119 a_299_66.t0 a_299_66.n0 408.174
R120 a_299_66.n0 a_299_66.t3 270.218
R121 a_299_66.n0 a_299_66.t1 195.971
R122 a_620_389.n0 a_620_389.t5 393.588
R123 a_620_389.n3 a_620_389.n2 307.182
R124 a_620_389.n0 a_620_389.t4 267.547
R125 a_620_389.n2 a_620_389.n1 184.051
R126 a_620_389.n3 a_620_389.t3 162.342
R127 a_620_389.n1 a_620_389.t0 106.635
R128 a_620_389.n2 a_620_389.n0 83.2
R129 a_620_389.t1 a_620_389.n3 74.787
R130 a_620_389.n1 a_620_389.t2 38.572
R131 a_780_389.t0 a_780_389.t1 102.148
R132 a_1767_21.n2 a_1767_21.t6 1015.03
R133 a_1767_21.n5 a_1767_21.n4 491.4
R134 a_1767_21.n0 a_1767_21.t5 239.392
R135 a_1767_21.n1 a_1767_21.t7 212.079
R136 a_1767_21.n3 a_1767_21.n2 181.032
R137 a_1767_21.n2 a_1767_21.t4 178.584
R138 a_1767_21.n0 a_1767_21.t3 154.239
R139 a_1767_21.n1 a_1767_21.t8 139.779
R140 a_1767_21.n1 a_1767_21.n0 132.915
R141 a_1767_21.n3 a_1767_21.t2 131.071
R142 a_1767_21.n4 a_1767_21.n1 97.924
R143 a_1767_21.n4 a_1767_21.n3 64.011
R144 a_1767_21.n5 a_1767_21.t1 63.321
R145 a_1767_21.t0 a_1767_21.n5 63.321
R146 a_2324_47.t0 a_2324_47.n1 259.364
R147 a_2324_47.n0 a_2324_47.t3 254.387
R148 a_2324_47.n0 a_2324_47.t2 211.007
R149 a_2324_47.n1 a_2324_47.t1 202.108
R150 a_2324_47.n1 a_2324_47.n0 76
R151 VGND.n1 VGND.t3 197.787
R152 VGND.n41 VGND.t6 159.774
R153 VGND.n43 VGND.t10 149.495
R154 VGND.n30 VGND.t11 148.719
R155 VGND.n9 VGND.t1 117.142
R156 VGND.n10 VGND.n9 113.205
R157 VGND.n2 VGND.n0 110.988
R158 VGND.n20 VGND.n19 107.239
R159 VGND.n50 VGND.n49 107.239
R160 VGND.n19 VGND.t0 72.857
R161 VGND.n19 VGND.t7 60.579
R162 VGND.n9 VGND.t5 52.857
R163 VGND.n0 VGND.t2 33.461
R164 VGND.n0 VGND.t4 33.461
R165 VGND.n49 VGND.t8 24.923
R166 VGND.n49 VGND.t9 24.923
R167 VGND.n11 VGND.n10 15.058
R168 VGND.n4 VGND.n3 4.65
R169 VGND.n6 VGND.n5 4.65
R170 VGND.n8 VGND.n7 4.65
R171 VGND.n12 VGND.n11 4.65
R172 VGND.n14 VGND.n13 4.65
R173 VGND.n16 VGND.n15 4.65
R174 VGND.n18 VGND.n17 4.65
R175 VGND.n21 VGND.n20 4.65
R176 VGND.n23 VGND.n22 4.65
R177 VGND.n25 VGND.n24 4.65
R178 VGND.n27 VGND.n26 4.65
R179 VGND.n29 VGND.n28 4.65
R180 VGND.n32 VGND.n31 4.65
R181 VGND.n34 VGND.n33 4.65
R182 VGND.n36 VGND.n35 4.65
R183 VGND.n38 VGND.n37 4.65
R184 VGND.n40 VGND.n39 4.65
R185 VGND.n42 VGND.n41 4.65
R186 VGND.n44 VGND.n43 4.65
R187 VGND.n46 VGND.n45 4.65
R188 VGND.n48 VGND.n47 4.65
R189 VGND.n2 VGND.n1 4.509
R190 VGND.n31 VGND.n30 4.141
R191 VGND.n51 VGND.n50 3.932
R192 VGND.n4 VGND.n2 0.141
R193 VGND.n51 VGND.n48 0.137
R194 VGND.n6 VGND.n4 0.119
R195 VGND.n8 VGND.n6 0.119
R196 VGND.n12 VGND.n8 0.119
R197 VGND.n14 VGND.n12 0.119
R198 VGND.n16 VGND.n14 0.119
R199 VGND.n18 VGND.n16 0.119
R200 VGND.n21 VGND.n18 0.119
R201 VGND.n23 VGND.n21 0.119
R202 VGND.n25 VGND.n23 0.119
R203 VGND.n27 VGND.n25 0.119
R204 VGND.n29 VGND.n27 0.119
R205 VGND.n32 VGND.n29 0.119
R206 VGND.n34 VGND.n32 0.119
R207 VGND.n36 VGND.n34 0.119
R208 VGND.n38 VGND.n36 0.119
R209 VGND.n40 VGND.n38 0.119
R210 VGND.n42 VGND.n40 0.119
R211 VGND.n44 VGND.n42 0.119
R212 VGND.n46 VGND.n44 0.119
R213 VGND.n48 VGND.n46 0.119
R214 VGND VGND.n51 0.11
R215 a_1079_413.n3 a_1079_413.n2 393.455
R216 a_1079_413.n1 a_1079_413.t4 339.006
R217 a_1079_413.n2 a_1079_413.n0 193.393
R218 a_1079_413.n1 a_1079_413.t5 168.699
R219 a_1079_413.n2 a_1079_413.n1 157.693
R220 a_1079_413.n3 a_1079_413.t3 128.988
R221 a_1079_413.n0 a_1079_413.t1 71.666
R222 a_1079_413.t0 a_1079_413.n3 63.321
R223 a_1079_413.n0 a_1079_413.t2 45
R224 a_1245_303.n0 a_1245_303.t4 365.917
R225 a_1245_303.n3 a_1245_303.n2 352.126
R226 a_1245_303.n2 a_1245_303.n1 177.291
R227 a_1245_303.n0 a_1245_303.t5 158.39
R228 a_1245_303.n2 a_1245_303.n0 151.67
R229 a_1245_303.n3 a_1245_303.t2 72.702
R230 a_1245_303.n1 a_1245_303.t3 63.333
R231 a_1245_303.t1 a_1245_303.n3 50.422
R232 a_1245_303.n1 a_1245_303.t0 26.77
R233 a_1592_47.n1 a_1592_47.t5 1025.84
R234 a_1592_47.n1 a_1592_47.t4 412.282
R235 a_1592_47.n3 a_1592_47.n2 342.717
R236 a_1592_47.n2 a_1592_47.n0 210.387
R237 a_1592_47.n2 a_1592_47.n1 144.894
R238 a_1592_47.n0 a_1592_47.t3 70
R239 a_1592_47.t1 a_1592_47.n3 68.011
R240 a_1592_47.n3 a_1592_47.t2 63.321
R241 a_1592_47.n0 a_1592_47.t0 61.666
R242 a_1701_47.t0 a_1701_47.t1 93.516
R243 a_1758_413.t0 a_1758_413.t1 121.952
R244 a_1946_47.t0 a_1946_47.t1 70
R245 SCD.n0 SCD.t0 248.765
R246 SCD.n0 SCD.t1 191.996
R247 SCD SCD.n0 79.072
R248 a_817_66.t1 a_817_66.t0 60
R249 SCE.t2 SCE.t3 729.319
R250 SCE.n0 SCE.t0 273.133
R251 SCE.n1 SCE.t2 215.9
R252 SCE.n1 SCE.n0 145.294
R253 SCE.n0 SCE.t1 138.173
R254 SCE SCE.n1 83.053
R255  SCE 34.974
R256 a_538_389.t0 a_538_389.t1 94.851
R257 RESET_B.n6 RESET_B.t0 2023.69
R258 RESET_B.n2 RESET_B.t2 396.265
R259 RESET_B.n6 RESET_B.t3 205.8
R260 RESET_B.n3 RESET_B.t1 126.39
R261 RESET_B.n3 RESET_B.n2 12.45
R262 RESET_B.n9 RESET_B 11.255
R263 RESET_B.n7 RESET_B.n6 9.81
R264 RESET_B.n4 RESET_B.n3 9.3
R265 RESET_B.n7 RESET_B 5.451
R266 RESET_B.n9 RESET_B.n8 4.659
R267 RESET_B.n5 RESET_B.n4 3.772
R268 RESET_B RESET_B.n9 3.751
R269 RESET_B.n4 RESET_B.n1 3.2
R270 RESET_B.n8 RESET_B.n5 2.364
R271 RESET_B.n8 RESET_B.n7 1.73
R272 RESET_B.n1 RESET_B.n0 0.685
R273 D.n0 D.t0 234.941
R274 D.n0 D.t1 164.248
R275 D.n1 D.n0 76
R276  D.n1 22.551
R277 D.n1 D 5.818
R278 a_569_119.t0 a_569_119.t1 60
R279 a_1187_47.t1 a_1187_47.t0 111.393
R280 a_1293_47.t0 a_1293_47.t1 60
R281 a_1191_413.n0 a_1191_413.t2 738.672
R282 a_1191_413.n0 a_1191_413.t1 63.321
R283 a_1191_413.t0 a_1191_413.n0 63.321
R284 Q.n2 Q.t1 207.372
R285 Q.n0 Q.t0 117.423
R286 Q.n1 Q 89.6
R287 Q.n1 Q.n0 64.808
R288 Q Q.n1 16
R289 Q.n0 Q 10.092
R290 Q.n2 Q 9.019
R291 Q Q.n2 7.458
R292 Q.n1 Q 0.738
R293 Q_N Q_N.t1 236.044
R294 Q_N Q_N.t0 199.212
R295 CLK.n0 CLK.t0 428.577
R296 CLK.n0 CLK.t1 426.167
R297 CLK.n1 CLK.n0 76
R298 CLK.n1 CLK 10.422
R299 CLK CLK.n1 2.011
C0 VPB VPWR 0.26fF
C1 VPWR VGND 0.12fF
C2 VPWR Q 0.11fF
C3 RESET_B VGND 0.35fF
C4 VPWR Q_N 0.13fF
C5 SCD VGND 0.11fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__sdfrbp_2.ext - technology: sky130A

.subckt sky130_fd_sc_hd__sdfrbp_2 VPWR VGND Q_N Q SCE SCD D RESET_B CLK VNB VPB
X0 a_193_47.t0 a_27_47.t2 VPWR.t15 VPB.t20 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_780_389.t1 a_299_66.t2 a_620_389.t5 VPB.t21 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=540000u l=150000u
X2 a_1245_303.t1 a_1079_413.t4 VPWR.t3 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X3 VPWR.t12 a_1592_47.t4 a_1767_21.t1 VPB.t12 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 VGND.t8 a_1767_21.t3 Q.t3 VNB.t11 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 VGND.t5 a_1767_21.t4 a_1701_47.t0 VNB.t10 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 a_1758_413.t1 a_193_47.t2 a_1592_47.t0 VPB.t14 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7 a_1767_21.t2 a_1592_47.t5 a_1946_47.t1 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 VPWR.t9 a_1767_21.t5 a_2135_47.t0 VPB.t9 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X9 VGND.t11 SCD.t0 a_817_66.t1 VNB.t16 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=180000u
X10 a_538_389.t0 SCE.t0 VPWR.t2 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=540000u l=150000u
X11 VPWR.t14 SCD.t1 a_780_389.t0 VPB.t17 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=540000u l=150000u
X12 VPWR.t6 SCE.t1 a_299_66.t0 VPB.t6 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=540000u l=150000u
X13 a_1767_21.t0 RESET_B.t0 VPWR.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14 a_193_47.t1 a_27_47.t3 VGND.t12 VNB.t20 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X15 a_620_389.t1 D.t0 a_569_119.t0 VNB.t7 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16 a_1187_47.t0 a_193_47.t3 a_1079_413.t1 VNB.t13 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X17 Q.t1 a_1767_21.t6 VPWR.t10 VPB.t10 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X18 a_1293_47.t1 a_1245_303.t4 a_1187_47.t1 VNB.t17 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19 VPWR.t8 a_1245_303.t5 a_1191_413.t1 VPB.t8 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20 Q.t2 a_1767_21.t7 VGND.t7 VNB.t9 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X21 a_620_389.t3 D.t1 a_538_389.t1 VPB.t15 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=540000u l=150000u
X22 a_1191_413.t2 a_27_47.t4 a_1079_413.t3 VPB.t19 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23 Q_N.t3 a_2135_47.t2 VGND.t2 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X24 a_569_119.t1 a_299_66.t3 VGND.t13 VNB.t21 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X25 VPWR.t11 a_1767_21.t8 a_1758_413.t0 VPB.t11 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X26 VGND.t0 RESET_B.t1 a_1293_47.t0 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X27 VPWR.t4 a_2135_47.t3 Q_N.t1 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X28 a_1079_413.t2 a_27_47.t5 a_620_389.t4 VNB.t19 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X29 VGND.t6 a_1767_21.t9 a_2135_47.t1 VNB.t8 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X30 a_1191_413.t0 RESET_B.t2 VPWR.t1 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X31 Q_N.t0 a_2135_47.t4 VPWR.t5 VPB.t5 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X32 a_1701_47.t1 a_27_47.t6 a_1592_47.t3 VNB.t18 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X33 a_1946_47.t0 RESET_B.t3 VGND.t1 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X34 VPWR.t7 a_1767_21.t10 Q.t0 VPB.t7 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X35 a_1592_47.t1 a_193_47.t4 a_1245_303.t0 VNB.t12 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X36 VGND.t4 SCE.t2 a_299_66.t1 VNB.t5 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X37 a_1592_47.t2 a_27_47.t7 a_1245_303.t3 VPB.t18 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X38 a_1245_303.t2 a_1079_413.t5 VGND.t9 VNB.t14 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X39 a_1079_413.t0 a_193_47.t5 a_620_389.t2 VPB.t13 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X40 VGND.t3 a_2135_47.t5 Q_N.t2 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X41 VPWR.t13 CLK.t0 a_27_47.t0 VPB.t16 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X42 a_817_66.t0 SCE.t3 a_620_389.t0 VNB.t6 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=500000u
X43 VGND.t10 CLK.t1 a_27_47.t1 VNB.t15 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
R0 a_27_47.n1 a_27_47.t4 534.047
R1 a_27_47.n0 a_27_47.t7 489.903
R2 a_27_47.n1 a_27_47.t5 276.816
R3 a_27_47.t0 a_27_47.n9 243.743
R4 a_27_47.n7 a_27_47.t2 238.856
R5 a_27_47.n0 a_27_47.t6 204.42
R6 a_27_47.n3 a_27_47.t1 175.866
R7 a_27_47.n5 a_27_47.t3 156.738
R8 a_27_47.n2 a_27_47.n0 14.808
R9 a_27_47.n6 a_27_47.n5 12.496
R10 a_27_47.n2 a_27_47.n1 11.633
R11 a_27_47.n8 a_27_47.n7 9.3
R12 a_27_47.n9 a_27_47.n2 6.029
R13 a_27_47.n4 a_27_47.n3 2.844
R14 a_27_47.n7 a_27_47.n6 2.677
R15 a_27_47.n9 a_27_47.n8 1.13
R16 a_27_47.n8 a_27_47.n4 0.609
R17 VPWR.n23 VPWR.t3 514.01
R18 VPWR.n39 VPWR.t14 408.48
R19 VPWR.n10 VPWR.t12 370.56
R20 VPWR.n48 VPWR.n47 323.37
R21 VPWR.n58 VPWR.n57 311.893
R22 VPWR.n15 VPWR.n14 310.932
R23 VPWR.n6 VPWR.n5 309.178
R24 VPWR.n1 VPWR.n0 307.239
R25 VPWR.n28 VPWR.n27 292.5
R26 VPWR.n2 VPWR.t4 166.684
R27 VPWR.n14 VPWR.t11 114.916
R28 VPWR.n27 VPWR.t1 103.19
R29 VPWR.n27 VPWR.t8 93.809
R30 VPWR.n14 VPWR.t0 63.321
R31 VPWR.n5 VPWR.t9 50.789
R32 VPWR.n47 VPWR.t2 49.25
R33 VPWR.n47 VPWR.t6 49.25
R34 VPWR.n5 VPWR.t10 38.707
R35 VPWR.n0 VPWR.t7 32.505
R36 VPWR.n57 VPWR.t13 29.55
R37 VPWR.n0 VPWR.t5 26.595
R38 VPWR.n57 VPWR.t15 26.595
R39 VPWR.n49 VPWR.n48 9.411
R40 VPWR.n4 VPWR.n3 4.65
R41 VPWR.n7 VPWR.n6 4.65
R42 VPWR.n9 VPWR.n8 4.65
R43 VPWR.n11 VPWR.n10 4.65
R44 VPWR.n13 VPWR.n12 4.65
R45 VPWR.n16 VPWR.n15 4.65
R46 VPWR.n18 VPWR.n17 4.65
R47 VPWR.n20 VPWR.n19 4.65
R48 VPWR.n22 VPWR.n21 4.65
R49 VPWR.n24 VPWR.n23 4.65
R50 VPWR.n26 VPWR.n25 4.65
R51 VPWR.n30 VPWR.n29 4.65
R52 VPWR.n32 VPWR.n31 4.65
R53 VPWR.n34 VPWR.n33 4.65
R54 VPWR.n36 VPWR.n35 4.65
R55 VPWR.n38 VPWR.n37 4.65
R56 VPWR.n40 VPWR.n39 4.65
R57 VPWR.n42 VPWR.n41 4.65
R58 VPWR.n44 VPWR.n43 4.65
R59 VPWR.n46 VPWR.n45 4.65
R60 VPWR.n50 VPWR.n49 4.65
R61 VPWR.n52 VPWR.n51 4.65
R62 VPWR.n54 VPWR.n53 4.65
R63 VPWR.n56 VPWR.n55 4.65
R64 VPWR.n59 VPWR.n58 3.958
R65 VPWR.n2 VPWR.n1 3.842
R66 VPWR.n29 VPWR.n28 2.702
R67 VPWR.n4 VPWR.n2 0.231
R68 VPWR.n59 VPWR.n56 0.137
R69 VPWR VPWR.n59 0.121
R70 VPWR.n7 VPWR.n4 0.119
R71 VPWR.n9 VPWR.n7 0.119
R72 VPWR.n11 VPWR.n9 0.119
R73 VPWR.n13 VPWR.n11 0.119
R74 VPWR.n16 VPWR.n13 0.119
R75 VPWR.n18 VPWR.n16 0.119
R76 VPWR.n20 VPWR.n18 0.119
R77 VPWR.n22 VPWR.n20 0.119
R78 VPWR.n24 VPWR.n22 0.119
R79 VPWR.n26 VPWR.n24 0.119
R80 VPWR.n30 VPWR.n26 0.119
R81 VPWR.n32 VPWR.n30 0.119
R82 VPWR.n34 VPWR.n32 0.119
R83 VPWR.n36 VPWR.n34 0.119
R84 VPWR.n38 VPWR.n36 0.119
R85 VPWR.n40 VPWR.n38 0.119
R86 VPWR.n42 VPWR.n40 0.119
R87 VPWR.n44 VPWR.n42 0.119
R88 VPWR.n46 VPWR.n44 0.119
R89 VPWR.n50 VPWR.n46 0.119
R90 VPWR.n52 VPWR.n50 0.119
R91 VPWR.n54 VPWR.n52 0.119
R92 VPWR.n56 VPWR.n54 0.119
R93 a_193_47.n1 a_193_47.t4 266.53
R94 a_193_47.n0 a_193_47.t3 265.71
R95 a_193_47.n1 a_193_47.t2 231.814
R96 a_193_47.n3 a_193_47.t1 210.139
R97 a_193_47.n0 a_193_47.t5 146.401
R98 a_193_47.t0 a_193_47.n3 38.199
R99 a_193_47.n2 a_193_47.n1 7.332
R100 a_193_47.n3 a_193_47.n2 6.062
R101 a_193_47.n2 a_193_47.n0 3.302
R102 VPB.t20 VPB.t6 774.312
R103 VPB.t17 VPB.t13 637.547
R104 VPB.t12 VPB.t9 556.386
R105 VPB.t1 VPB.t3 556.386
R106 VPB.t15 VPB.t21 511.784
R107 VPB.t8 VPB.t1 337.383
R108 VPB.t13 VPB.t19 331.464
R109 VPB.t11 VPB.t0 313.707
R110 VPB.t9 VPB.t10 281.152
R111 VPB.t3 VPB.t18 281.152
R112 VPB.t21 VPB.t17 275.084
R113 VPB.t10 VPB.t7 272.274
R114 VPB.t6 VPB.t2 268.686
R115 VPB.t7 VPB.t5 266.355
R116 VPB.t2 VPB.t15 262.289
R117 VPB.t16 VPB.t20 257.476
R118 VPB.t18 VPB.t14 254.517
R119 VPB.t5 VPB.t4 248.598
R120 VPB.t0 VPB.t12 248.598
R121 VPB.t19 VPB.t8 248.598
R122 VPB.t14 VPB.t11 242.679
R123 VPB VPB.t16 177.57
R124 a_299_66.n0 a_299_66.t2 1032.99
R125 a_299_66.t0 a_299_66.n0 408.174
R126 a_299_66.n0 a_299_66.t3 270.218
R127 a_299_66.n0 a_299_66.t1 195.971
R128 a_620_389.n0 a_620_389.t2 393.588
R129 a_620_389.n3 a_620_389.n2 307.182
R130 a_620_389.n0 a_620_389.t4 267.547
R131 a_620_389.n2 a_620_389.n1 184.051
R132 a_620_389.t3 a_620_389.n3 162.342
R133 a_620_389.n1 a_620_389.t0 106.635
R134 a_620_389.n2 a_620_389.n0 83.2
R135 a_620_389.n3 a_620_389.t5 74.787
R136 a_620_389.n1 a_620_389.t1 38.572
R137 a_780_389.t0 a_780_389.t1 102.148
R138 a_1079_413.n3 a_1079_413.n2 393.455
R139 a_1079_413.n1 a_1079_413.t4 339.006
R140 a_1079_413.n2 a_1079_413.n0 193.393
R141 a_1079_413.n1 a_1079_413.t5 168.699
R142 a_1079_413.n2 a_1079_413.n1 157.693
R143 a_1079_413.t0 a_1079_413.n3 128.988
R144 a_1079_413.n0 a_1079_413.t2 71.666
R145 a_1079_413.n3 a_1079_413.t3 63.321
R146 a_1079_413.n0 a_1079_413.t1 45
R147 a_1245_303.n0 a_1245_303.t4 365.917
R148 a_1245_303.n3 a_1245_303.n2 352.126
R149 a_1245_303.n2 a_1245_303.n1 177.291
R150 a_1245_303.n0 a_1245_303.t5 158.39
R151 a_1245_303.n2 a_1245_303.n0 151.67
R152 a_1245_303.n3 a_1245_303.t3 72.702
R153 a_1245_303.n1 a_1245_303.t0 63.333
R154 a_1245_303.t1 a_1245_303.n3 50.422
R155 a_1245_303.n1 a_1245_303.t2 26.77
R156 a_1592_47.n1 a_1592_47.t5 1025.84
R157 a_1592_47.n1 a_1592_47.t4 412.282
R158 a_1592_47.n3 a_1592_47.n2 342.717
R159 a_1592_47.n2 a_1592_47.n0 210.387
R160 a_1592_47.n2 a_1592_47.n1 144.894
R161 a_1592_47.n0 a_1592_47.t1 70
R162 a_1592_47.n3 a_1592_47.t2 68.011
R163 a_1592_47.t0 a_1592_47.n3 63.321
R164 a_1592_47.n0 a_1592_47.t3 61.666
R165 a_1767_21.n4 a_1767_21.t8 1015.03
R166 a_1767_21.n7 a_1767_21.n6 499.934
R167 a_1767_21.n2 a_1767_21.t5 257.066
R168 a_1767_21.n0 a_1767_21.t10 212.079
R169 a_1767_21.n1 a_1767_21.t6 212.079
R170 a_1767_21.n5 a_1767_21.n4 181.032
R171 a_1767_21.n4 a_1767_21.t4 178.584
R172 a_1767_21.n3 a_1767_21.t9 176.733
R173 a_1767_21.n0 a_1767_21.t3 139.779
R174 a_1767_21.n1 a_1767_21.t7 139.779
R175 a_1767_21.n5 a_1767_21.t2 131.071
R176 a_1767_21.n6 a_1767_21.n3 102.396
R177 a_1767_21.n6 a_1767_21.n5 72.423
R178 a_1767_21.n2 a_1767_21.n1 69.378
R179 a_1767_21.n1 a_1767_21.n0 67.187
R180 a_1767_21.n7 a_1767_21.t1 63.321
R181 a_1767_21.t0 a_1767_21.n7 63.321
R182 a_1767_21.n3 a_1767_21.n2 0.73
R183 Q Q.n0 310.785
R184 Q Q.n1 110.054
R185 Q.n0 Q.t1 34.475
R186 Q.n1 Q.t2 32.307
R187 Q.n0 Q.t0 26.595
R188 Q.n1 Q.t3 24.923
R189 VGND.n48 VGND.t13 159.774
R190 VGND.n50 VGND.t4 149.495
R191 VGND.n37 VGND.t11 148.719
R192 VGND.n1 VGND.n0 128.641
R193 VGND.n16 VGND.t1 117.142
R194 VGND.n2 VGND.t3 115.662
R195 VGND.n17 VGND.n16 113.205
R196 VGND.n6 VGND.n5 110.187
R197 VGND.n27 VGND.n26 107.239
R198 VGND.n57 VGND.n56 107.239
R199 VGND.n26 VGND.t0 72.857
R200 VGND.n26 VGND.t9 60.579
R201 VGND.n16 VGND.t5 52.857
R202 VGND.n5 VGND.t6 48.571
R203 VGND.n5 VGND.t7 32.571
R204 VGND.n0 VGND.t8 30.461
R205 VGND.n0 VGND.t2 24.923
R206 VGND.n56 VGND.t12 24.923
R207 VGND.n56 VGND.t10 24.923
R208 VGND.n18 VGND.n17 15.058
R209 VGND.n4 VGND.n3 4.65
R210 VGND.n7 VGND.n6 4.65
R211 VGND.n9 VGND.n8 4.65
R212 VGND.n11 VGND.n10 4.65
R213 VGND.n13 VGND.n12 4.65
R214 VGND.n15 VGND.n14 4.65
R215 VGND.n19 VGND.n18 4.65
R216 VGND.n21 VGND.n20 4.65
R217 VGND.n23 VGND.n22 4.65
R218 VGND.n25 VGND.n24 4.65
R219 VGND.n28 VGND.n27 4.65
R220 VGND.n30 VGND.n29 4.65
R221 VGND.n32 VGND.n31 4.65
R222 VGND.n34 VGND.n33 4.65
R223 VGND.n36 VGND.n35 4.65
R224 VGND.n39 VGND.n38 4.65
R225 VGND.n41 VGND.n40 4.65
R226 VGND.n43 VGND.n42 4.65
R227 VGND.n45 VGND.n44 4.65
R228 VGND.n47 VGND.n46 4.65
R229 VGND.n49 VGND.n48 4.65
R230 VGND.n51 VGND.n50 4.65
R231 VGND.n53 VGND.n52 4.65
R232 VGND.n55 VGND.n54 4.65
R233 VGND.n38 VGND.n37 4.141
R234 VGND.n2 VGND.n1 4.062
R235 VGND.n58 VGND.n57 3.932
R236 VGND.n4 VGND.n2 0.211
R237 VGND.n58 VGND.n55 0.137
R238 VGND.n7 VGND.n4 0.119
R239 VGND.n9 VGND.n7 0.119
R240 VGND.n11 VGND.n9 0.119
R241 VGND.n13 VGND.n11 0.119
R242 VGND.n15 VGND.n13 0.119
R243 VGND.n19 VGND.n15 0.119
R244 VGND.n21 VGND.n19 0.119
R245 VGND.n23 VGND.n21 0.119
R246 VGND.n25 VGND.n23 0.119
R247 VGND.n28 VGND.n25 0.119
R248 VGND.n30 VGND.n28 0.119
R249 VGND.n32 VGND.n30 0.119
R250 VGND.n34 VGND.n32 0.119
R251 VGND.n36 VGND.n34 0.119
R252 VGND.n39 VGND.n36 0.119
R253 VGND.n41 VGND.n39 0.119
R254 VGND.n43 VGND.n41 0.119
R255 VGND.n45 VGND.n43 0.119
R256 VGND.n47 VGND.n45 0.119
R257 VGND.n49 VGND.n47 0.119
R258 VGND.n51 VGND.n49 0.119
R259 VGND.n53 VGND.n51 0.119
R260 VGND.n55 VGND.n53 0.119
R261 VGND VGND.n58 0.11
R262 VNB VNB.t15 26484.6
R263 VNB.t16 VNB.t19 6619.1
R264 VNB.t2 VNB.t8 6211.76
R265 VNB.t5 VNB.t21 6123.67
R266 VNB.t20 VNB.t5 5321.88
R267 VNB.t10 VNB.t1 4820.59
R268 VNB.t6 VNB.t16 3558.82
R269 VNB.t0 VNB.t14 3550.91
R270 VNB.t19 VNB.t13 3548.39
R271 VNB.t12 VNB.t18 3526.47
R272 VNB.t13 VNB.t17 3476.38
R273 VNB.t18 VNB.t10 3105.88
R274 VNB.t7 VNB.t6 2863.63
R275 VNB.t1 VNB.t2 2555.88
R276 VNB.t17 VNB.t0 2329.41
R277 VNB.t21 VNB.t7 2329.41
R278 VNB.t14 VNB.t12 2280.14
R279 VNB.t8 VNB.t9 2279.52
R280 VNB.t9 VNB.t11 2224.18
R281 VNB.t11 VNB.t3 2175.82
R282 VNB.t3 VNB.t4 2030.77
R283 VNB.t15 VNB.t20 2030.77
R284 a_1701_47.t0 a_1701_47.t1 93.516
R285 a_1758_413.t0 a_1758_413.t1 121.952
R286 a_1946_47.t0 a_1946_47.t1 70
R287 a_2135_47.n2 a_2135_47.t1 251.659
R288 a_2135_47.t0 a_2135_47.n2 242.552
R289 a_2135_47.n1 a_2135_47.t4 212.079
R290 a_2135_47.n0 a_2135_47.t3 212.079
R291 a_2135_47.n2 a_2135_47.n1 177.562
R292 a_2135_47.n1 a_2135_47.t2 139.779
R293 a_2135_47.n0 a_2135_47.t5 139.779
R294 a_2135_47.n1 a_2135_47.n0 61.345
R295 SCD.n0 SCD.t0 248.765
R296 SCD.n0 SCD.t1 191.996
R297 SCD SCD.n0 79.072
R298 a_817_66.t1 a_817_66.t0 60
R299 SCE.t2 SCE.t3 729.319
R300 SCE.n0 SCE.t0 273.133
R301 SCE.n1 SCE.t2 215.9
R302 SCE.n1 SCE.n0 145.294
R303 SCE.n0 SCE.t1 138.173
R304 SCE SCE.n1 83.053
R305  SCE 34.974
R306 a_538_389.t0 a_538_389.t1 94.851
R307 RESET_B.n6 RESET_B.t0 2023.69
R308 RESET_B.n2 RESET_B.t2 396.265
R309 RESET_B.n6 RESET_B.t3 205.8
R310 RESET_B.n3 RESET_B.t1 126.39
R311 RESET_B.n3 RESET_B.n2 12.45
R312 RESET_B.n9 RESET_B 11.255
R313 RESET_B.n7 RESET_B.n6 9.81
R314 RESET_B.n4 RESET_B.n3 9.3
R315 RESET_B.n7 RESET_B 5.451
R316 RESET_B.n9 RESET_B.n8 4.659
R317 RESET_B.n5 RESET_B.n4 3.772
R318 RESET_B RESET_B.n9 3.751
R319 RESET_B.n4 RESET_B.n1 3.2
R320 RESET_B.n8 RESET_B.n5 2.364
R321 RESET_B.n8 RESET_B.n7 1.73
R322 RESET_B.n1 RESET_B.n0 0.685
R323 D.n0 D.t0 234.941
R324 D.n0 D.t1 164.248
R325 D.n1 D.n0 76
R326  D.n1 22.551
R327 D.n1 D 5.818
R328 a_569_119.t0 a_569_119.t1 60
R329 a_1187_47.t1 a_1187_47.t0 111.393
R330 a_1293_47.t0 a_1293_47.t1 60
R331 a_1191_413.t0 a_1191_413.n0 738.672
R332 a_1191_413.n0 a_1191_413.t1 63.321
R333 a_1191_413.n0 a_1191_413.t2 63.321
R334 Q_N Q_N.n0 141.505
R335 Q_N Q_N.n1 70.257
R336 Q_N.n0 Q_N.t1 26.595
R337 Q_N.n0 Q_N.t0 26.595
R338 Q_N.n1 Q_N.t2 24.923
R339 Q_N.n1 Q_N.t3 24.923
R340 CLK.n0 CLK.t0 428.577
R341 CLK.n0 CLK.t1 426.167
R342 CLK.n1 CLK.n0 76
R343 CLK.n1 CLK 10.422
R344 CLK CLK.n1 2.011
C0 VPWR Q_N 0.23fF
C1 SCD VGND 0.11fF
C2 VPB VPWR 0.27fF
C3 VGND Q 0.15fF
C4 VPWR VGND 0.14fF
C5 VGND Q_N 0.24fF
C6 RESET_B VGND 0.35fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__sdfrtn_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__sdfrtn_1 VPWR VGND SCE SCD D RESET_B CLK_N Q VNB VPB
X0 a_193_47.t1 a_27_47.t2 VPWR.t10 VPB.t16 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_780_389.t1 a_299_66.t2 a_620_389.t2 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=540000u l=150000u
X2 a_1245_303.t1 a_1079_413.t4 VPWR.t3 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X3 VPWR.t6 a_1592_47.t4 a_1767_21.t2 VPB.t7 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 VGND.t7 a_1767_21.t3 a_1701_47.t0 VNB.t9 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 a_1758_413.t1 a_27_47.t3 a_1592_47.t2 VPB.t15 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 a_1767_21.t1 a_1592_47.t5 a_1946_47.t1 VNB.t17 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7 VGND.t0 SCD.t0 a_817_66.t1 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=180000u
X8 a_538_389.t0 SCE.t0 VPWR.t11 VPB.t17 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=540000u l=150000u
X9 VPWR.t4 SCD.t1 a_780_389.t0 VPB.t5 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=540000u l=150000u
X10 VPWR.t5 SCE.t1 a_299_66.t0 VPB.t6 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=540000u l=150000u
X11 a_1767_21.t0 RESET_B.t0 VPWR.t7 VPB.t8 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12 a_193_47.t0 a_27_47.t4 VGND.t9 VNB.t15 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 a_620_389.t5 D.t0 a_569_119.t0 VNB.t16 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14 a_1187_47.t1 a_27_47.t5 a_1079_413.t3 VNB.t14 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X15 a_1293_47.t0 a_1245_303.t4 a_1187_47.t0 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16 VPWR.t2 a_1245_303.t5 a_1191_413.t0 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17 a_620_389.t1 D.t1 a_538_389.t1 VPB.t10 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=540000u l=150000u
X18 a_1191_413.t2 a_193_47.t2 a_1079_413.t1 VPB.t13 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19 a_569_119.t1 a_299_66.t3 VGND.t8 VNB.t10 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20 VPWR.t0 a_1767_21.t4 a_1758_413.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21 VGND.t3 RESET_B.t1 a_1293_47.t1 VNB.t5 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22 Q.t1 a_1767_21.t5 VPWR.t1 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X23 Q.t0 a_1767_21.t6 VGND.t6 VNB.t8 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X24 a_1079_413.t0 a_193_47.t3 a_620_389.t3 VNB.t12 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X25 a_1191_413.t1 RESET_B.t2 VPWR.t8 VPB.t9 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X26 a_1701_47.t1 a_193_47.t4 a_1592_47.t1 VNB.t11 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X27 a_1946_47.t0 RESET_B.t3 VGND.t4 VNB.t6 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X28 a_1592_47.t3 a_27_47.t6 a_1245_303.t3 VNB.t13 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X29 VGND.t1 SCE.t2 a_299_66.t1 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X30 a_1592_47.t0 a_193_47.t5 a_1245_303.t2 VPB.t12 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X31 a_1245_303.t0 a_1079_413.t5 VGND.t2 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X32 a_1079_413.t2 a_27_47.t7 a_620_389.t4 VPB.t14 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X33 VPWR.t9 CLK_N.t0 a_27_47.t1 VPB.t11 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X34 a_817_66.t0 SCE.t3 a_620_389.t0 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=500000u
X35 VGND.t5 CLK_N.t1 a_27_47.t0 VNB.t7 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
R0 a_27_47.n1 a_27_47.t6 266.53
R1 a_27_47.n0 a_27_47.t5 265.71
R2 a_27_47.n3 a_27_47.t2 241.534
R3 a_27_47.n1 a_27_47.t3 231.814
R4 a_27_47.t1 a_27_47.n5 205.348
R5 a_27_47.n4 a_27_47.t0 178.71
R6 a_27_47.n3 a_27_47.t4 169.234
R7 a_27_47.n0 a_27_47.t7 146.401
R8 a_27_47.n4 a_27_47.n3 76
R9 a_27_47.n5 a_27_47.n4 40.733
R10 a_27_47.n5 a_27_47.n2 8.697
R11 a_27_47.n2 a_27_47.n1 7.332
R12 a_27_47.n2 a_27_47.n0 3.302
R13 VPWR.n13 VPWR.t3 514.01
R14 VPWR.n29 VPWR.t4 408.48
R15 VPWR.n0 VPWR.t6 370.56
R16 VPWR.n38 VPWR.n37 323.37
R17 VPWR.n48 VPWR.n47 311.893
R18 VPWR.n5 VPWR.n4 310.932
R19 VPWR.n18 VPWR.n17 292.5
R20 VPWR.n1 VPWR.t1 155.579
R21 VPWR.n4 VPWR.t0 114.916
R22 VPWR.n17 VPWR.t8 103.19
R23 VPWR.n17 VPWR.t2 93.809
R24 VPWR.n4 VPWR.t7 63.321
R25 VPWR.n37 VPWR.t11 49.25
R26 VPWR.n37 VPWR.t5 49.25
R27 VPWR.n47 VPWR.t9 29.55
R28 VPWR.n47 VPWR.t10 26.595
R29 VPWR.n39 VPWR.n38 9.411
R30 VPWR.n3 VPWR.n2 4.65
R31 VPWR.n6 VPWR.n5 4.65
R32 VPWR.n8 VPWR.n7 4.65
R33 VPWR.n10 VPWR.n9 4.65
R34 VPWR.n12 VPWR.n11 4.65
R35 VPWR.n14 VPWR.n13 4.65
R36 VPWR.n16 VPWR.n15 4.65
R37 VPWR.n20 VPWR.n19 4.65
R38 VPWR.n22 VPWR.n21 4.65
R39 VPWR.n24 VPWR.n23 4.65
R40 VPWR.n26 VPWR.n25 4.65
R41 VPWR.n28 VPWR.n27 4.65
R42 VPWR.n30 VPWR.n29 4.65
R43 VPWR.n32 VPWR.n31 4.65
R44 VPWR.n34 VPWR.n33 4.65
R45 VPWR.n36 VPWR.n35 4.65
R46 VPWR.n40 VPWR.n39 4.65
R47 VPWR.n42 VPWR.n41 4.65
R48 VPWR.n44 VPWR.n43 4.65
R49 VPWR.n46 VPWR.n45 4.65
R50 VPWR.n49 VPWR.n48 3.958
R51 VPWR.n1 VPWR.n0 3.252
R52 VPWR.n19 VPWR.n18 2.702
R53 VPWR.n3 VPWR.n1 0.774
R54 VPWR.n49 VPWR.n46 0.137
R55 VPWR VPWR.n49 0.121
R56 VPWR.n6 VPWR.n3 0.119
R57 VPWR.n8 VPWR.n6 0.119
R58 VPWR.n10 VPWR.n8 0.119
R59 VPWR.n12 VPWR.n10 0.119
R60 VPWR.n14 VPWR.n12 0.119
R61 VPWR.n16 VPWR.n14 0.119
R62 VPWR.n20 VPWR.n16 0.119
R63 VPWR.n22 VPWR.n20 0.119
R64 VPWR.n24 VPWR.n22 0.119
R65 VPWR.n26 VPWR.n24 0.119
R66 VPWR.n28 VPWR.n26 0.119
R67 VPWR.n30 VPWR.n28 0.119
R68 VPWR.n32 VPWR.n30 0.119
R69 VPWR.n34 VPWR.n32 0.119
R70 VPWR.n36 VPWR.n34 0.119
R71 VPWR.n40 VPWR.n36 0.119
R72 VPWR.n42 VPWR.n40 0.119
R73 VPWR.n44 VPWR.n42 0.119
R74 VPWR.n46 VPWR.n44 0.119
R75 a_193_47.n1 a_193_47.t2 534.047
R76 a_193_47.n0 a_193_47.t5 489.903
R77 a_193_47.n1 a_193_47.t3 276.816
R78 a_193_47.t1 a_193_47.n3 232.909
R79 a_193_47.n0 a_193_47.t4 204.42
R80 a_193_47.n3 a_193_47.t0 163.239
R81 a_193_47.n2 a_193_47.n0 14.808
R82 a_193_47.n2 a_193_47.n1 11.633
R83 a_193_47.n3 a_193_47.n2 7.904
R84 VPB.t16 VPB.t6 774.312
R85 VPB.t5 VPB.t14 637.547
R86 VPB.t7 VPB.t2 556.386
R87 VPB.t9 VPB.t4 556.386
R88 VPB.t10 VPB.t1 511.784
R89 VPB.t3 VPB.t9 337.383
R90 VPB.t14 VPB.t13 331.464
R91 VPB.t0 VPB.t8 313.707
R92 VPB.t4 VPB.t12 281.152
R93 VPB.t1 VPB.t5 275.084
R94 VPB.t6 VPB.t17 268.686
R95 VPB.t17 VPB.t10 262.289
R96 VPB.t11 VPB.t16 257.476
R97 VPB.t12 VPB.t15 254.517
R98 VPB.t8 VPB.t7 248.598
R99 VPB.t13 VPB.t3 248.598
R100 VPB.t15 VPB.t0 242.679
R101 VPB VPB.t11 177.57
R102 a_299_66.n0 a_299_66.t2 1032.99
R103 a_299_66.t0 a_299_66.n0 408.174
R104 a_299_66.n0 a_299_66.t3 270.218
R105 a_299_66.n0 a_299_66.t1 195.971
R106 a_620_389.n0 a_620_389.t4 393.588
R107 a_620_389.n3 a_620_389.n2 307.182
R108 a_620_389.n0 a_620_389.t3 267.547
R109 a_620_389.n2 a_620_389.n1 184.051
R110 a_620_389.t1 a_620_389.n3 162.342
R111 a_620_389.n1 a_620_389.t0 106.635
R112 a_620_389.n2 a_620_389.n0 83.2
R113 a_620_389.n3 a_620_389.t2 74.787
R114 a_620_389.n1 a_620_389.t5 38.572
R115 a_780_389.t0 a_780_389.t1 102.148
R116 a_1079_413.n3 a_1079_413.n2 393.455
R117 a_1079_413.n1 a_1079_413.t4 339.006
R118 a_1079_413.n2 a_1079_413.n0 193.393
R119 a_1079_413.n1 a_1079_413.t5 168.699
R120 a_1079_413.n2 a_1079_413.n1 157.693
R121 a_1079_413.n3 a_1079_413.t2 128.988
R122 a_1079_413.n0 a_1079_413.t0 71.666
R123 a_1079_413.t1 a_1079_413.n3 63.321
R124 a_1079_413.n0 a_1079_413.t3 45
R125 a_1245_303.n0 a_1245_303.t4 365.917
R126 a_1245_303.n3 a_1245_303.n2 352.126
R127 a_1245_303.n2 a_1245_303.n1 177.291
R128 a_1245_303.n0 a_1245_303.t5 158.39
R129 a_1245_303.n2 a_1245_303.n0 151.67
R130 a_1245_303.n3 a_1245_303.t2 72.702
R131 a_1245_303.n1 a_1245_303.t3 63.333
R132 a_1245_303.t1 a_1245_303.n3 50.422
R133 a_1245_303.n1 a_1245_303.t0 26.77
R134 a_1592_47.n1 a_1592_47.t5 1025.84
R135 a_1592_47.n1 a_1592_47.t4 412.282
R136 a_1592_47.n3 a_1592_47.n2 342.717
R137 a_1592_47.n2 a_1592_47.n0 210.387
R138 a_1592_47.n2 a_1592_47.n1 144.894
R139 a_1592_47.n0 a_1592_47.t3 70
R140 a_1592_47.t0 a_1592_47.n3 68.011
R141 a_1592_47.n3 a_1592_47.t2 63.321
R142 a_1592_47.n0 a_1592_47.t1 61.666
R143 a_1767_21.n1 a_1767_21.t4 1015.03
R144 a_1767_21.n4 a_1767_21.n3 491.4
R145 a_1767_21.n0 a_1767_21.t5 239.503
R146 a_1767_21.n2 a_1767_21.n1 181.032
R147 a_1767_21.n1 a_1767_21.t3 178.584
R148 a_1767_21.n0 a_1767_21.t6 167.203
R149 a_1767_21.n2 a_1767_21.t1 131.071
R150 a_1767_21.n3 a_1767_21.n0 86.24
R151 a_1767_21.n3 a_1767_21.n2 64.011
R152 a_1767_21.n4 a_1767_21.t2 63.321
R153 a_1767_21.t0 a_1767_21.n4 63.321
R154 a_1701_47.t0 a_1701_47.t1 93.516
R155 VGND.n0 VGND.t6 202.156
R156 VGND.n33 VGND.t8 159.774
R157 VGND.n35 VGND.t1 149.495
R158 VGND.n22 VGND.t0 148.719
R159 VGND.n1 VGND.t4 117.142
R160 VGND.n2 VGND.n1 113.205
R161 VGND.n12 VGND.n11 107.239
R162 VGND.n42 VGND.n41 107.239
R163 VGND.n11 VGND.t3 72.857
R164 VGND.n11 VGND.t2 60.579
R165 VGND.n1 VGND.t7 52.857
R166 VGND.n41 VGND.t9 24.923
R167 VGND.n41 VGND.t5 24.923
R168 VGND.n3 VGND.n2 15.058
R169 VGND.n4 VGND.n3 4.65
R170 VGND.n6 VGND.n5 4.65
R171 VGND.n8 VGND.n7 4.65
R172 VGND.n10 VGND.n9 4.65
R173 VGND.n13 VGND.n12 4.65
R174 VGND.n15 VGND.n14 4.65
R175 VGND.n17 VGND.n16 4.65
R176 VGND.n19 VGND.n18 4.65
R177 VGND.n21 VGND.n20 4.65
R178 VGND.n24 VGND.n23 4.65
R179 VGND.n26 VGND.n25 4.65
R180 VGND.n28 VGND.n27 4.65
R181 VGND.n30 VGND.n29 4.65
R182 VGND.n32 VGND.n31 4.65
R183 VGND.n34 VGND.n33 4.65
R184 VGND.n36 VGND.n35 4.65
R185 VGND.n38 VGND.n37 4.65
R186 VGND.n40 VGND.n39 4.65
R187 VGND.n23 VGND.n22 4.141
R188 VGND.n43 VGND.n42 3.932
R189 VGND.n4 VGND.n0 0.139
R190 VGND.n43 VGND.n40 0.137
R191 VGND.n6 VGND.n4 0.119
R192 VGND.n8 VGND.n6 0.119
R193 VGND.n10 VGND.n8 0.119
R194 VGND.n13 VGND.n10 0.119
R195 VGND.n15 VGND.n13 0.119
R196 VGND.n17 VGND.n15 0.119
R197 VGND.n19 VGND.n17 0.119
R198 VGND.n21 VGND.n19 0.119
R199 VGND.n24 VGND.n21 0.119
R200 VGND.n26 VGND.n24 0.119
R201 VGND.n28 VGND.n26 0.119
R202 VGND.n30 VGND.n28 0.119
R203 VGND.n32 VGND.n30 0.119
R204 VGND.n34 VGND.n32 0.119
R205 VGND.n36 VGND.n34 0.119
R206 VGND.n38 VGND.n36 0.119
R207 VGND.n40 VGND.n38 0.119
R208 VGND VGND.n43 0.11
R209 VNB VNB.t7 26484.6
R210 VNB.t0 VNB.t12 6619.1
R211 VNB.t2 VNB.t10 6123.67
R212 VNB.t17 VNB.t8 5483.65
R213 VNB.t15 VNB.t2 5321.88
R214 VNB.t9 VNB.t6 4820.59
R215 VNB.t1 VNB.t0 3558.82
R216 VNB.t5 VNB.t3 3550.91
R217 VNB.t12 VNB.t14 3548.39
R218 VNB.t13 VNB.t11 3526.47
R219 VNB.t14 VNB.t4 3476.38
R220 VNB.t11 VNB.t9 3105.88
R221 VNB.t16 VNB.t1 2863.63
R222 VNB.t6 VNB.t17 2555.88
R223 VNB.t4 VNB.t5 2329.41
R224 VNB.t10 VNB.t16 2329.41
R225 VNB.t3 VNB.t13 2280.14
R226 VNB.t7 VNB.t15 2030.77
R227 a_1758_413.t0 a_1758_413.t1 121.952
R228 a_1946_47.t0 a_1946_47.t1 70
R229 SCD.n0 SCD.t0 248.765
R230 SCD.n0 SCD.t1 191.996
R231 SCD SCD.n0 79.072
R232 a_817_66.t1 a_817_66.t0 60
R233 SCE.t2 SCE.t3 729.319
R234 SCE.n0 SCE.t0 273.133
R235 SCE.n1 SCE.t2 215.9
R236 SCE.n1 SCE.n0 145.294
R237 SCE.n0 SCE.t1 138.173
R238 SCE SCE.n1 83.053
R239  SCE 34.974
R240 a_538_389.t0 a_538_389.t1 94.851
R241 RESET_B.n6 RESET_B.t0 2023.69
R242 RESET_B.n2 RESET_B.t2 396.265
R243 RESET_B.n6 RESET_B.t3 205.8
R244 RESET_B.n3 RESET_B.t1 126.39
R245 RESET_B.n3 RESET_B.n2 12.45
R246 RESET_B.n9 RESET_B 11.255
R247 RESET_B.n7 RESET_B.n6 9.81
R248 RESET_B.n4 RESET_B.n3 9.3
R249 RESET_B.n7 RESET_B 5.451
R250 RESET_B.n9 RESET_B.n8 4.659
R251 RESET_B.n5 RESET_B.n4 3.772
R252 RESET_B RESET_B.n9 3.751
R253 RESET_B.n4 RESET_B.n1 3.2
R254 RESET_B.n8 RESET_B.n5 2.364
R255 RESET_B.n8 RESET_B.n7 1.73
R256 RESET_B.n1 RESET_B.n0 0.685
R257 D.n0 D.t0 234.941
R258 D.n0 D.t1 164.248
R259 D.n1 D.n0 76
R260  D.n1 22.551
R261 D.n1 D 5.818
R262 a_569_119.t0 a_569_119.t1 60
R263 a_1187_47.t0 a_1187_47.t1 111.393
R264 a_1293_47.t0 a_1293_47.t1 60
R265 a_1191_413.n0 a_1191_413.t1 738.672
R266 a_1191_413.t0 a_1191_413.n0 63.321
R267 a_1191_413.n0 a_1191_413.t2 63.321
R268 Q.n2 Q.t1 207.372
R269 Q.n0 Q.t0 117.423
R270 Q.n1 Q 89.6
R271 Q.n1 Q.n0 64.808
R272 Q Q.n1 16
R273 Q.n0 Q 10.092
R274 Q.n2 Q 9.019
R275 Q Q.n2 7.458
R276 Q.n1 Q 0.738
R277 CLK_N.n0 CLK_N.t0 428.577
R278 CLK_N.n0 CLK_N.t1 426.167
R279 CLK_N.n1 CLK_N.n0 76
R280 CLK_N.n1 CLK_N 10.422
R281 CLK_N CLK_N.n1 2.011
C0 VPWR Q 0.11fF
C1 RESET_B VGND 0.34fF
C2 SCD VGND 0.11fF
C3 VPB VPWR 0.23fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__sdfrtp_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__sdfrtp_1 VPWR VGND SCE SCD D RESET_B CLK Q VNB VPB
X0 a_193_47.t1 a_27_47.t2 VPWR.t0 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_780_389.t1 a_299_66.t2 a_620_389.t5 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=540000u l=150000u
X2 a_1245_303.t3 a_1079_413.t4 VPWR.t10 VPB.t16 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X3 VPWR.t3 a_1592_47.t4 a_1767_21.t2 VPB.t6 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 VGND.t6 a_1767_21.t3 a_1701_47.t1 VNB.t12 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 a_1758_413.t0 a_193_47.t2 a_1592_47.t2 VPB.t12 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 a_1767_21.t1 a_1592_47.t5 a_1946_47.t1 VNB.t13 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7 VGND.t2 SCD.t0 a_817_66.t1 VNB.t5 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=180000u
X8 a_538_389.t1 SCE.t0 VPWR.t1 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=540000u l=150000u
X9 VPWR.t6 SCD.t1 a_780_389.t0 VPB.t9 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=540000u l=150000u
X10 VPWR.t2 SCE.t1 a_299_66.t0 VPB.t5 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=540000u l=150000u
X11 a_1767_21.t0 RESET_B.t0 VPWR.t8 VPB.t13 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12 a_193_47.t0 a_27_47.t3 VGND.t0 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 a_620_389.t4 D.t0 a_569_119.t1 VNB.t10 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14 a_1187_47.t0 a_193_47.t3 a_1079_413.t2 VNB.t7 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X15 a_1293_47.t0 a_1245_303.t4 a_1187_47.t1 VNB.t14 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16 VPWR.t7 a_1245_303.t5 a_1191_413.t1 VPB.t10 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17 a_620_389.t3 D.t1 a_538_389.t0 VPB.t15 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=540000u l=150000u
X18 a_1191_413.t0 a_27_47.t4 a_1079_413.t1 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19 a_569_119.t0 a_299_66.t3 VGND.t7 VNB.t15 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20 VPWR.t4 a_1767_21.t4 a_1758_413.t1 VPB.t7 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21 VGND.t3 RESET_B.t1 a_1293_47.t1 VNB.t8 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22 Q.t0 a_1767_21.t5 VPWR.t5 VPB.t8 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X23 Q.t1 a_1767_21.t6 VGND.t5 VNB.t11 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X24 a_1079_413.t0 a_27_47.t5 a_620_389.t0 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X25 a_1191_413.t2 RESET_B.t2 VPWR.t9 VPB.t14 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X26 a_1701_47.t0 a_27_47.t6 a_1592_47.t0 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X27 a_1946_47.t0 RESET_B.t3 VGND.t4 VNB.t9 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X28 a_1592_47.t3 a_193_47.t4 a_1245_303.t1 VNB.t6 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X29 VGND.t1 SCE.t2 a_299_66.t1 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X30 a_1592_47.t1 a_27_47.t7 a_1245_303.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X31 a_1245_303.t2 a_1079_413.t5 VGND.t9 VNB.t17 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X32 a_1079_413.t3 a_193_47.t5 a_620_389.t2 VPB.t11 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X33 VPWR.t11 CLK.t0 a_27_47.t0 VPB.t17 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X34 a_817_66.t0 SCE.t3 a_620_389.t1 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=500000u
X35 VGND.t8 CLK.t1 a_27_47.t1 VNB.t16 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
R0 a_27_47.n1 a_27_47.t4 534.047
R1 a_27_47.n0 a_27_47.t7 489.903
R2 a_27_47.n1 a_27_47.t5 276.816
R3 a_27_47.t0 a_27_47.n9 243.743
R4 a_27_47.n7 a_27_47.t2 238.856
R5 a_27_47.n0 a_27_47.t6 204.42
R6 a_27_47.n3 a_27_47.t1 175.866
R7 a_27_47.n5 a_27_47.t3 156.738
R8 a_27_47.n2 a_27_47.n0 14.808
R9 a_27_47.n6 a_27_47.n5 12.496
R10 a_27_47.n2 a_27_47.n1 11.633
R11 a_27_47.n8 a_27_47.n7 9.3
R12 a_27_47.n9 a_27_47.n2 6.029
R13 a_27_47.n4 a_27_47.n3 2.844
R14 a_27_47.n7 a_27_47.n6 2.677
R15 a_27_47.n9 a_27_47.n8 1.13
R16 a_27_47.n8 a_27_47.n4 0.609
R17 VPWR.n13 VPWR.t10 514.01
R18 VPWR.n29 VPWR.t6 408.48
R19 VPWR.n0 VPWR.t3 370.56
R20 VPWR.n38 VPWR.n37 323.37
R21 VPWR.n48 VPWR.n47 311.893
R22 VPWR.n5 VPWR.n4 310.932
R23 VPWR.n18 VPWR.n17 292.5
R24 VPWR.n1 VPWR.t5 155.579
R25 VPWR.n4 VPWR.t4 114.916
R26 VPWR.n17 VPWR.t9 103.19
R27 VPWR.n17 VPWR.t7 93.809
R28 VPWR.n4 VPWR.t8 63.321
R29 VPWR.n37 VPWR.t1 49.25
R30 VPWR.n37 VPWR.t2 49.25
R31 VPWR.n47 VPWR.t11 29.55
R32 VPWR.n47 VPWR.t0 26.595
R33 VPWR.n39 VPWR.n38 9.411
R34 VPWR.n3 VPWR.n2 4.65
R35 VPWR.n6 VPWR.n5 4.65
R36 VPWR.n8 VPWR.n7 4.65
R37 VPWR.n10 VPWR.n9 4.65
R38 VPWR.n12 VPWR.n11 4.65
R39 VPWR.n14 VPWR.n13 4.65
R40 VPWR.n16 VPWR.n15 4.65
R41 VPWR.n20 VPWR.n19 4.65
R42 VPWR.n22 VPWR.n21 4.65
R43 VPWR.n24 VPWR.n23 4.65
R44 VPWR.n26 VPWR.n25 4.65
R45 VPWR.n28 VPWR.n27 4.65
R46 VPWR.n30 VPWR.n29 4.65
R47 VPWR.n32 VPWR.n31 4.65
R48 VPWR.n34 VPWR.n33 4.65
R49 VPWR.n36 VPWR.n35 4.65
R50 VPWR.n40 VPWR.n39 4.65
R51 VPWR.n42 VPWR.n41 4.65
R52 VPWR.n44 VPWR.n43 4.65
R53 VPWR.n46 VPWR.n45 4.65
R54 VPWR.n49 VPWR.n48 3.958
R55 VPWR.n1 VPWR.n0 3.252
R56 VPWR.n19 VPWR.n18 2.702
R57 VPWR.n3 VPWR.n1 0.774
R58 VPWR.n49 VPWR.n46 0.137
R59 VPWR VPWR.n49 0.121
R60 VPWR.n6 VPWR.n3 0.119
R61 VPWR.n8 VPWR.n6 0.119
R62 VPWR.n10 VPWR.n8 0.119
R63 VPWR.n12 VPWR.n10 0.119
R64 VPWR.n14 VPWR.n12 0.119
R65 VPWR.n16 VPWR.n14 0.119
R66 VPWR.n20 VPWR.n16 0.119
R67 VPWR.n22 VPWR.n20 0.119
R68 VPWR.n24 VPWR.n22 0.119
R69 VPWR.n26 VPWR.n24 0.119
R70 VPWR.n28 VPWR.n26 0.119
R71 VPWR.n30 VPWR.n28 0.119
R72 VPWR.n32 VPWR.n30 0.119
R73 VPWR.n34 VPWR.n32 0.119
R74 VPWR.n36 VPWR.n34 0.119
R75 VPWR.n40 VPWR.n36 0.119
R76 VPWR.n42 VPWR.n40 0.119
R77 VPWR.n44 VPWR.n42 0.119
R78 VPWR.n46 VPWR.n44 0.119
R79 a_193_47.n1 a_193_47.t4 266.53
R80 a_193_47.n0 a_193_47.t3 265.71
R81 a_193_47.n1 a_193_47.t2 231.814
R82 a_193_47.n3 a_193_47.t0 210.139
R83 a_193_47.n0 a_193_47.t5 146.401
R84 a_193_47.t1 a_193_47.n3 38.199
R85 a_193_47.n2 a_193_47.n1 7.332
R86 a_193_47.n3 a_193_47.n2 6.062
R87 a_193_47.n2 a_193_47.n0 3.302
R88 VPB.t2 VPB.t5 774.312
R89 VPB.t9 VPB.t11 637.547
R90 VPB.t6 VPB.t8 556.386
R91 VPB.t14 VPB.t16 556.386
R92 VPB.t15 VPB.t3 511.784
R93 VPB.t10 VPB.t14 337.383
R94 VPB.t11 VPB.t1 331.464
R95 VPB.t7 VPB.t13 313.707
R96 VPB.t16 VPB.t0 281.152
R97 VPB.t3 VPB.t9 275.084
R98 VPB.t5 VPB.t4 268.686
R99 VPB.t4 VPB.t15 262.289
R100 VPB.t17 VPB.t2 257.476
R101 VPB.t0 VPB.t12 254.517
R102 VPB.t13 VPB.t6 248.598
R103 VPB.t1 VPB.t10 248.598
R104 VPB.t12 VPB.t7 242.679
R105 VPB VPB.t17 177.57
R106 a_299_66.n0 a_299_66.t2 1032.99
R107 a_299_66.t0 a_299_66.n0 408.174
R108 a_299_66.n0 a_299_66.t3 270.218
R109 a_299_66.n0 a_299_66.t1 195.971
R110 a_620_389.n0 a_620_389.t2 393.588
R111 a_620_389.n3 a_620_389.n2 307.182
R112 a_620_389.n0 a_620_389.t0 267.547
R113 a_620_389.n2 a_620_389.n1 184.051
R114 a_620_389.t3 a_620_389.n3 162.342
R115 a_620_389.n1 a_620_389.t1 106.635
R116 a_620_389.n2 a_620_389.n0 83.2
R117 a_620_389.n3 a_620_389.t5 74.787
R118 a_620_389.n1 a_620_389.t4 38.572
R119 a_780_389.t0 a_780_389.t1 102.148
R120 a_1079_413.n3 a_1079_413.n2 393.455
R121 a_1079_413.n1 a_1079_413.t4 339.006
R122 a_1079_413.n2 a_1079_413.n0 193.393
R123 a_1079_413.n1 a_1079_413.t5 168.699
R124 a_1079_413.n2 a_1079_413.n1 157.693
R125 a_1079_413.n3 a_1079_413.t3 128.988
R126 a_1079_413.n0 a_1079_413.t0 71.666
R127 a_1079_413.t1 a_1079_413.n3 63.321
R128 a_1079_413.n0 a_1079_413.t2 45
R129 a_1245_303.n0 a_1245_303.t4 365.917
R130 a_1245_303.n3 a_1245_303.n2 352.126
R131 a_1245_303.n2 a_1245_303.n1 177.291
R132 a_1245_303.n0 a_1245_303.t5 158.39
R133 a_1245_303.n2 a_1245_303.n0 151.67
R134 a_1245_303.n3 a_1245_303.t0 72.702
R135 a_1245_303.n1 a_1245_303.t1 63.333
R136 a_1245_303.t3 a_1245_303.n3 50.422
R137 a_1245_303.n1 a_1245_303.t2 26.77
R138 a_1592_47.n1 a_1592_47.t5 1025.84
R139 a_1592_47.n1 a_1592_47.t4 412.282
R140 a_1592_47.n3 a_1592_47.n2 342.717
R141 a_1592_47.n2 a_1592_47.n0 210.387
R142 a_1592_47.n2 a_1592_47.n1 144.894
R143 a_1592_47.n0 a_1592_47.t3 70
R144 a_1592_47.t1 a_1592_47.n3 68.011
R145 a_1592_47.n3 a_1592_47.t2 63.321
R146 a_1592_47.n0 a_1592_47.t0 61.666
R147 a_1767_21.n1 a_1767_21.t4 1015.03
R148 a_1767_21.n4 a_1767_21.n3 491.4
R149 a_1767_21.n0 a_1767_21.t5 239.503
R150 a_1767_21.n2 a_1767_21.n1 181.032
R151 a_1767_21.n1 a_1767_21.t3 178.584
R152 a_1767_21.n0 a_1767_21.t6 167.203
R153 a_1767_21.n2 a_1767_21.t1 131.071
R154 a_1767_21.n3 a_1767_21.n0 86.24
R155 a_1767_21.n3 a_1767_21.n2 64.011
R156 a_1767_21.n4 a_1767_21.t2 63.321
R157 a_1767_21.t0 a_1767_21.n4 63.321
R158 a_1701_47.t1 a_1701_47.t0 93.516
R159 VGND.n0 VGND.t5 202.156
R160 VGND.n33 VGND.t7 159.774
R161 VGND.n35 VGND.t1 149.495
R162 VGND.n22 VGND.t2 148.719
R163 VGND.n1 VGND.t4 117.142
R164 VGND.n2 VGND.n1 113.205
R165 VGND.n12 VGND.n11 107.239
R166 VGND.n42 VGND.n41 107.239
R167 VGND.n11 VGND.t3 72.857
R168 VGND.n11 VGND.t9 60.579
R169 VGND.n1 VGND.t6 52.857
R170 VGND.n41 VGND.t0 24.923
R171 VGND.n41 VGND.t8 24.923
R172 VGND.n3 VGND.n2 15.058
R173 VGND.n4 VGND.n3 4.65
R174 VGND.n6 VGND.n5 4.65
R175 VGND.n8 VGND.n7 4.65
R176 VGND.n10 VGND.n9 4.65
R177 VGND.n13 VGND.n12 4.65
R178 VGND.n15 VGND.n14 4.65
R179 VGND.n17 VGND.n16 4.65
R180 VGND.n19 VGND.n18 4.65
R181 VGND.n21 VGND.n20 4.65
R182 VGND.n24 VGND.n23 4.65
R183 VGND.n26 VGND.n25 4.65
R184 VGND.n28 VGND.n27 4.65
R185 VGND.n30 VGND.n29 4.65
R186 VGND.n32 VGND.n31 4.65
R187 VGND.n34 VGND.n33 4.65
R188 VGND.n36 VGND.n35 4.65
R189 VGND.n38 VGND.n37 4.65
R190 VGND.n40 VGND.n39 4.65
R191 VGND.n23 VGND.n22 4.141
R192 VGND.n43 VGND.n42 3.932
R193 VGND.n4 VGND.n0 0.139
R194 VGND.n43 VGND.n40 0.137
R195 VGND.n6 VGND.n4 0.119
R196 VGND.n8 VGND.n6 0.119
R197 VGND.n10 VGND.n8 0.119
R198 VGND.n13 VGND.n10 0.119
R199 VGND.n15 VGND.n13 0.119
R200 VGND.n17 VGND.n15 0.119
R201 VGND.n19 VGND.n17 0.119
R202 VGND.n21 VGND.n19 0.119
R203 VGND.n24 VGND.n21 0.119
R204 VGND.n26 VGND.n24 0.119
R205 VGND.n28 VGND.n26 0.119
R206 VGND.n30 VGND.n28 0.119
R207 VGND.n32 VGND.n30 0.119
R208 VGND.n34 VGND.n32 0.119
R209 VGND.n36 VGND.n34 0.119
R210 VGND.n38 VGND.n36 0.119
R211 VGND.n40 VGND.n38 0.119
R212 VGND VGND.n43 0.11
R213 VNB VNB.t16 26484.6
R214 VNB.t5 VNB.t1 6619.1
R215 VNB.t3 VNB.t15 6123.67
R216 VNB.t13 VNB.t11 5483.65
R217 VNB.t2 VNB.t3 5321.88
R218 VNB.t12 VNB.t9 4820.59
R219 VNB.t4 VNB.t5 3558.82
R220 VNB.t8 VNB.t17 3550.91
R221 VNB.t1 VNB.t7 3548.39
R222 VNB.t6 VNB.t0 3526.47
R223 VNB.t7 VNB.t14 3476.38
R224 VNB.t0 VNB.t12 3105.88
R225 VNB.t10 VNB.t4 2863.63
R226 VNB.t9 VNB.t13 2555.88
R227 VNB.t14 VNB.t8 2329.41
R228 VNB.t15 VNB.t10 2329.41
R229 VNB.t17 VNB.t6 2280.14
R230 VNB.t16 VNB.t2 2030.77
R231 a_1758_413.t0 a_1758_413.t1 121.952
R232 a_1946_47.t0 a_1946_47.t1 70
R233 SCD.n0 SCD.t0 248.765
R234 SCD.n0 SCD.t1 191.996
R235 SCD SCD.n0 79.072
R236 a_817_66.t1 a_817_66.t0 60
R237 SCE.t2 SCE.t3 729.319
R238 SCE.n0 SCE.t0 273.133
R239 SCE.n1 SCE.t2 215.9
R240 SCE.n1 SCE.n0 145.294
R241 SCE.n0 SCE.t1 138.173
R242 SCE SCE.n1 83.053
R243  SCE 34.974
R244 a_538_389.t0 a_538_389.t1 94.851
R245 RESET_B.n6 RESET_B.t0 2023.69
R246 RESET_B.n2 RESET_B.t2 396.265
R247 RESET_B.n6 RESET_B.t3 205.8
R248 RESET_B.n3 RESET_B.t1 126.39
R249 RESET_B.n3 RESET_B.n2 12.45
R250 RESET_B.n9 RESET_B 11.255
R251 RESET_B.n7 RESET_B.n6 9.81
R252 RESET_B.n4 RESET_B.n3 9.3
R253 RESET_B.n7 RESET_B 5.451
R254 RESET_B.n9 RESET_B.n8 4.659
R255 RESET_B.n5 RESET_B.n4 3.772
R256 RESET_B RESET_B.n9 3.751
R257 RESET_B.n4 RESET_B.n1 3.2
R258 RESET_B.n8 RESET_B.n5 2.364
R259 RESET_B.n8 RESET_B.n7 1.73
R260 RESET_B.n1 RESET_B.n0 0.685
R261 D.n0 D.t0 234.941
R262 D.n0 D.t1 164.248
R263 D.n1 D.n0 76
R264  D.n1 22.551
R265 D.n1 D 5.818
R266 a_569_119.t0 a_569_119.t1 60
R267 a_1187_47.t1 a_1187_47.t0 111.393
R268 a_1293_47.t0 a_1293_47.t1 60
R269 a_1191_413.n0 a_1191_413.t2 738.672
R270 a_1191_413.n0 a_1191_413.t1 63.321
R271 a_1191_413.t0 a_1191_413.n0 63.321
R272 Q.n2 Q.t0 207.372
R273 Q.n0 Q.t1 117.423
R274 Q.n1 Q 89.6
R275 Q.n1 Q.n0 64.808
R276 Q Q.n1 16
R277 Q.n0 Q 10.092
R278 Q.n2 Q 9.019
R279 Q Q.n2 7.458
R280 Q.n1 Q 0.738
R281 CLK.n0 CLK.t0 428.577
R282 CLK.n0 CLK.t1 426.167
R283 CLK.n1 CLK.n0 76
R284 CLK.n1 CLK 10.422
R285 CLK CLK.n1 2.011
C0 SCD VGND 0.11fF
C1 VPB VPWR 0.23fF
C2 RESET_B VGND 0.34fF
C3 VPWR Q 0.11fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__sdfrtp_2.ext - technology: sky130A

.subckt sky130_fd_sc_hd__sdfrtp_2 VPWR VGND SCE SCD D RESET_B CLK Q VNB VPB
X0 a_193_47.t1 a_27_47.t2 VPWR.t6 VPB.t9 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_780_389.t0 a_299_66.t2 a_620_389.t2 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=540000u l=150000u
X2 a_1245_303.t2 a_1079_413.t4 VPWR.t10 VPB.t13 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X3 VPWR.t5 a_1592_47.t4 a_1767_21.t2 VPB.t6 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 VGND.t3 a_1767_21.t3 a_1701_47.t1 VNB.t8 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 a_1758_413.t1 a_193_47.t2 a_1592_47.t3 VPB.t18 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 a_1767_21.t1 a_1592_47.t5 a_1946_47.t1 VNB.t5 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7 VGND.t9 SCD.t0 a_817_66.t1 VNB.t15 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=180000u
X8 a_538_389.t1 SCE.t0 VPWR.t7 VPB.t10 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=540000u l=150000u
X9 VPWR.t12 SCD.t1 a_780_389.t1 VPB.t15 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=540000u l=150000u
X10 VPWR.t8 SCE.t1 a_299_66.t0 VPB.t11 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=540000u l=150000u
X11 a_1767_21.t0 RESET_B.t0 VPWR.t1 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12 a_193_47.t0 a_27_47.t3 VGND.t2 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 a_620_389.t3 D.t0 a_569_119.t1 VNB.t14 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14 a_1187_47.t1 a_193_47.t3 a_1079_413.t2 VNB.t18 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X15 VGND.t5 a_1767_21.t4 Q.t3 VNB.t7 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X16 a_1293_47.t0 a_1245_303.t4 a_1187_47.t0 VNB.t10 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17 VPWR.t3 a_1767_21.t5 Q.t1 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X18 VPWR.t0 a_1245_303.t5 a_1191_413.t1 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19 a_620_389.t4 D.t1 a_538_389.t0 VPB.t16 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=540000u l=150000u
X20 a_1191_413.t0 a_27_47.t4 a_1079_413.t0 VPB.t8 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21 a_569_119.t0 a_299_66.t3 VGND.t7 VNB.t12 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22 VPWR.t4 a_1767_21.t6 a_1758_413.t0 VPB.t5 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23 VGND.t0 RESET_B.t1 a_1293_47.t1 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24 Q.t0 a_1767_21.t7 VPWR.t9 VPB.t12 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X25 Q.t2 a_1767_21.t8 VGND.t4 VNB.t6 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X26 a_1079_413.t1 a_27_47.t5 a_620_389.t0 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X27 a_1191_413.t2 RESET_B.t2 VPWR.t2 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X28 a_1701_47.t0 a_27_47.t6 a_1592_47.t1 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X29 a_1946_47.t0 RESET_B.t3 VGND.t1 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X30 a_1592_47.t2 a_193_47.t4 a_1245_303.t3 VNB.t17 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X31 VGND.t6 SCE.t2 a_299_66.t1 VNB.t9 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X32 a_1592_47.t0 a_27_47.t7 a_1245_303.t0 VPB.t7 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X33 a_1245_303.t1 a_1079_413.t5 VGND.t8 VNB.t13 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X34 a_1079_413.t3 a_193_47.t5 a_620_389.t5 VPB.t17 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X35 VPWR.t11 CLK.t0 a_27_47.t0 VPB.t14 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X36 a_817_66.t0 SCE.t3 a_620_389.t1 VNB.t11 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=500000u
X37 VGND.t10 CLK.t1 a_27_47.t1 VNB.t16 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
R0 a_27_47.n1 a_27_47.t4 534.047
R1 a_27_47.n0 a_27_47.t7 489.903
R2 a_27_47.n1 a_27_47.t5 276.816
R3 a_27_47.t0 a_27_47.n9 243.743
R4 a_27_47.n7 a_27_47.t2 238.856
R5 a_27_47.n0 a_27_47.t6 204.42
R6 a_27_47.n3 a_27_47.t1 175.866
R7 a_27_47.n5 a_27_47.t3 156.738
R8 a_27_47.n2 a_27_47.n0 14.808
R9 a_27_47.n6 a_27_47.n5 12.496
R10 a_27_47.n2 a_27_47.n1 11.633
R11 a_27_47.n8 a_27_47.n7 9.3
R12 a_27_47.n9 a_27_47.n2 6.029
R13 a_27_47.n4 a_27_47.n3 2.844
R14 a_27_47.n7 a_27_47.n6 2.677
R15 a_27_47.n9 a_27_47.n8 1.13
R16 a_27_47.n8 a_27_47.n4 0.609
R17 VPWR.n15 VPWR.t10 514.01
R18 VPWR.n31 VPWR.t12 408.48
R19 VPWR.n2 VPWR.t5 370.56
R20 VPWR.n40 VPWR.n39 323.37
R21 VPWR.n50 VPWR.n49 311.893
R22 VPWR.n7 VPWR.n6 310.932
R23 VPWR.n20 VPWR.n19 292.5
R24 VPWR.n1 VPWR.t3 158.724
R25 VPWR.n0 VPWR.t9 152.716
R26 VPWR.n6 VPWR.t4 114.916
R27 VPWR.n19 VPWR.t2 103.19
R28 VPWR.n19 VPWR.t0 93.809
R29 VPWR.n6 VPWR.t1 63.321
R30 VPWR.n39 VPWR.t7 49.25
R31 VPWR.n39 VPWR.t8 49.25
R32 VPWR.n49 VPWR.t11 29.55
R33 VPWR.n49 VPWR.t6 26.595
R34 VPWR.n41 VPWR.n40 9.411
R35 VPWR.n3 VPWR.n2 4.65
R36 VPWR.n5 VPWR.n4 4.65
R37 VPWR.n8 VPWR.n7 4.65
R38 VPWR.n10 VPWR.n9 4.65
R39 VPWR.n12 VPWR.n11 4.65
R40 VPWR.n14 VPWR.n13 4.65
R41 VPWR.n16 VPWR.n15 4.65
R42 VPWR.n18 VPWR.n17 4.65
R43 VPWR.n22 VPWR.n21 4.65
R44 VPWR.n24 VPWR.n23 4.65
R45 VPWR.n26 VPWR.n25 4.65
R46 VPWR.n28 VPWR.n27 4.65
R47 VPWR.n30 VPWR.n29 4.65
R48 VPWR.n32 VPWR.n31 4.65
R49 VPWR.n34 VPWR.n33 4.65
R50 VPWR.n36 VPWR.n35 4.65
R51 VPWR.n38 VPWR.n37 4.65
R52 VPWR.n42 VPWR.n41 4.65
R53 VPWR.n44 VPWR.n43 4.65
R54 VPWR.n46 VPWR.n45 4.65
R55 VPWR.n48 VPWR.n47 4.65
R56 VPWR.n51 VPWR.n50 3.958
R57 VPWR.n1 VPWR.n0 3.84
R58 VPWR.n21 VPWR.n20 2.702
R59 VPWR.n3 VPWR.n1 0.24
R60 VPWR.n51 VPWR.n48 0.137
R61 VPWR VPWR.n51 0.121
R62 VPWR.n5 VPWR.n3 0.119
R63 VPWR.n8 VPWR.n5 0.119
R64 VPWR.n10 VPWR.n8 0.119
R65 VPWR.n12 VPWR.n10 0.119
R66 VPWR.n14 VPWR.n12 0.119
R67 VPWR.n16 VPWR.n14 0.119
R68 VPWR.n18 VPWR.n16 0.119
R69 VPWR.n22 VPWR.n18 0.119
R70 VPWR.n24 VPWR.n22 0.119
R71 VPWR.n26 VPWR.n24 0.119
R72 VPWR.n28 VPWR.n26 0.119
R73 VPWR.n30 VPWR.n28 0.119
R74 VPWR.n32 VPWR.n30 0.119
R75 VPWR.n34 VPWR.n32 0.119
R76 VPWR.n36 VPWR.n34 0.119
R77 VPWR.n38 VPWR.n36 0.119
R78 VPWR.n42 VPWR.n38 0.119
R79 VPWR.n44 VPWR.n42 0.119
R80 VPWR.n46 VPWR.n44 0.119
R81 VPWR.n48 VPWR.n46 0.119
R82 a_193_47.n1 a_193_47.t4 266.53
R83 a_193_47.n0 a_193_47.t3 265.71
R84 a_193_47.n1 a_193_47.t2 231.814
R85 a_193_47.n3 a_193_47.t0 210.139
R86 a_193_47.n0 a_193_47.t5 146.401
R87 a_193_47.t1 a_193_47.n3 38.199
R88 a_193_47.n2 a_193_47.n1 7.332
R89 a_193_47.n3 a_193_47.n2 6.062
R90 a_193_47.n2 a_193_47.n0 3.302
R91 VPB.t9 VPB.t11 774.312
R92 VPB.t15 VPB.t17 637.547
R93 VPB.t6 VPB.t12 556.386
R94 VPB.t3 VPB.t13 556.386
R95 VPB.t16 VPB.t1 511.784
R96 VPB.t0 VPB.t3 337.383
R97 VPB.t17 VPB.t8 331.464
R98 VPB.t5 VPB.t2 313.707
R99 VPB.t13 VPB.t7 281.152
R100 VPB.t1 VPB.t15 275.084
R101 VPB.t11 VPB.t10 268.686
R102 VPB.t10 VPB.t16 262.289
R103 VPB.t14 VPB.t9 257.476
R104 VPB.t7 VPB.t18 254.517
R105 VPB.t12 VPB.t4 248.598
R106 VPB.t2 VPB.t6 248.598
R107 VPB.t8 VPB.t0 248.598
R108 VPB.t18 VPB.t5 242.679
R109 VPB VPB.t14 177.57
R110 a_299_66.n0 a_299_66.t2 1032.99
R111 a_299_66.t0 a_299_66.n0 408.174
R112 a_299_66.n0 a_299_66.t3 270.218
R113 a_299_66.n0 a_299_66.t1 195.971
R114 a_620_389.n0 a_620_389.t5 393.588
R115 a_620_389.n3 a_620_389.n2 307.182
R116 a_620_389.n0 a_620_389.t0 267.547
R117 a_620_389.n2 a_620_389.n1 184.051
R118 a_620_389.n3 a_620_389.t4 162.342
R119 a_620_389.n1 a_620_389.t1 106.635
R120 a_620_389.n2 a_620_389.n0 83.2
R121 a_620_389.t2 a_620_389.n3 74.787
R122 a_620_389.n1 a_620_389.t3 38.572
R123 a_780_389.t0 a_780_389.t1 102.148
R124 a_1079_413.n3 a_1079_413.n2 393.455
R125 a_1079_413.n1 a_1079_413.t4 339.006
R126 a_1079_413.n2 a_1079_413.n0 193.393
R127 a_1079_413.n1 a_1079_413.t5 168.699
R128 a_1079_413.n2 a_1079_413.n1 157.693
R129 a_1079_413.n3 a_1079_413.t3 128.988
R130 a_1079_413.n0 a_1079_413.t1 71.666
R131 a_1079_413.t0 a_1079_413.n3 63.321
R132 a_1079_413.n0 a_1079_413.t2 45
R133 a_1245_303.n0 a_1245_303.t4 365.917
R134 a_1245_303.n3 a_1245_303.n2 352.126
R135 a_1245_303.n2 a_1245_303.n1 177.291
R136 a_1245_303.n0 a_1245_303.t5 158.39
R137 a_1245_303.n2 a_1245_303.n0 151.67
R138 a_1245_303.n3 a_1245_303.t0 72.702
R139 a_1245_303.n1 a_1245_303.t3 63.333
R140 a_1245_303.t2 a_1245_303.n3 50.422
R141 a_1245_303.n1 a_1245_303.t1 26.77
R142 a_1592_47.n1 a_1592_47.t5 1025.84
R143 a_1592_47.n1 a_1592_47.t4 412.282
R144 a_1592_47.n3 a_1592_47.n2 342.717
R145 a_1592_47.n2 a_1592_47.n0 210.387
R146 a_1592_47.n2 a_1592_47.n1 144.894
R147 a_1592_47.n0 a_1592_47.t2 70
R148 a_1592_47.t0 a_1592_47.n3 68.011
R149 a_1592_47.n3 a_1592_47.t3 63.321
R150 a_1592_47.n0 a_1592_47.t1 61.666
R151 a_1767_21.n2 a_1767_21.t6 1015.03
R152 a_1767_21.n5 a_1767_21.n4 491.4
R153 a_1767_21.n0 a_1767_21.t5 212.079
R154 a_1767_21.n1 a_1767_21.t7 212.079
R155 a_1767_21.n3 a_1767_21.n2 181.032
R156 a_1767_21.n2 a_1767_21.t3 178.584
R157 a_1767_21.n0 a_1767_21.t4 139.779
R158 a_1767_21.n1 a_1767_21.t8 139.779
R159 a_1767_21.n3 a_1767_21.t1 131.071
R160 a_1767_21.n4 a_1767_21.n1 97.924
R161 a_1767_21.n4 a_1767_21.n3 64.011
R162 a_1767_21.n5 a_1767_21.t2 63.321
R163 a_1767_21.t0 a_1767_21.n5 63.321
R164 a_1767_21.n1 a_1767_21.n0 61.345
R165 a_1701_47.t1 a_1701_47.t0 93.516
R166 VGND.n1 VGND.t5 202.621
R167 VGND.n0 VGND.t4 197.787
R168 VGND.n40 VGND.t7 159.774
R169 VGND.n42 VGND.t6 149.495
R170 VGND.n29 VGND.t9 148.719
R171 VGND.n8 VGND.t1 117.142
R172 VGND.n9 VGND.n8 113.205
R173 VGND.n19 VGND.n18 107.239
R174 VGND.n49 VGND.n48 107.239
R175 VGND.n18 VGND.t0 72.857
R176 VGND.n18 VGND.t8 60.579
R177 VGND.n8 VGND.t3 52.857
R178 VGND.n48 VGND.t2 24.923
R179 VGND.n48 VGND.t10 24.923
R180 VGND.n10 VGND.n9 15.058
R181 VGND.n3 VGND.n2 4.65
R182 VGND.n5 VGND.n4 4.65
R183 VGND.n7 VGND.n6 4.65
R184 VGND.n11 VGND.n10 4.65
R185 VGND.n13 VGND.n12 4.65
R186 VGND.n15 VGND.n14 4.65
R187 VGND.n17 VGND.n16 4.65
R188 VGND.n20 VGND.n19 4.65
R189 VGND.n22 VGND.n21 4.65
R190 VGND.n24 VGND.n23 4.65
R191 VGND.n26 VGND.n25 4.65
R192 VGND.n28 VGND.n27 4.65
R193 VGND.n31 VGND.n30 4.65
R194 VGND.n33 VGND.n32 4.65
R195 VGND.n35 VGND.n34 4.65
R196 VGND.n37 VGND.n36 4.65
R197 VGND.n39 VGND.n38 4.65
R198 VGND.n41 VGND.n40 4.65
R199 VGND.n43 VGND.n42 4.65
R200 VGND.n45 VGND.n44 4.65
R201 VGND.n47 VGND.n46 4.65
R202 VGND.n1 VGND.n0 4.4
R203 VGND.n30 VGND.n29 4.141
R204 VGND.n50 VGND.n49 3.932
R205 VGND.n3 VGND.n1 0.25
R206 VGND.n50 VGND.n47 0.137
R207 VGND.n5 VGND.n3 0.119
R208 VGND.n7 VGND.n5 0.119
R209 VGND.n11 VGND.n7 0.119
R210 VGND.n13 VGND.n11 0.119
R211 VGND.n15 VGND.n13 0.119
R212 VGND.n17 VGND.n15 0.119
R213 VGND.n20 VGND.n17 0.119
R214 VGND.n22 VGND.n20 0.119
R215 VGND.n24 VGND.n22 0.119
R216 VGND.n26 VGND.n24 0.119
R217 VGND.n28 VGND.n26 0.119
R218 VGND.n31 VGND.n28 0.119
R219 VGND.n33 VGND.n31 0.119
R220 VGND.n35 VGND.n33 0.119
R221 VGND.n37 VGND.n35 0.119
R222 VGND.n39 VGND.n37 0.119
R223 VGND.n41 VGND.n39 0.119
R224 VGND.n43 VGND.n41 0.119
R225 VGND.n45 VGND.n43 0.119
R226 VGND.n47 VGND.n45 0.119
R227 VGND VGND.n50 0.11
R228 VNB VNB.t16 26484.6
R229 VNB.t15 VNB.t3 6619.1
R230 VNB.t9 VNB.t12 6123.67
R231 VNB.t5 VNB.t6 5483.65
R232 VNB.t4 VNB.t9 5321.88
R233 VNB.t8 VNB.t1 4820.59
R234 VNB.t11 VNB.t15 3558.82
R235 VNB.t0 VNB.t13 3550.91
R236 VNB.t3 VNB.t18 3548.39
R237 VNB.t17 VNB.t2 3526.47
R238 VNB.t18 VNB.t10 3476.38
R239 VNB.t2 VNB.t8 3105.88
R240 VNB.t14 VNB.t11 2863.63
R241 VNB.t1 VNB.t5 2555.88
R242 VNB.t10 VNB.t0 2329.41
R243 VNB.t12 VNB.t14 2329.41
R244 VNB.t13 VNB.t17 2280.14
R245 VNB.t6 VNB.t7 2030.77
R246 VNB.t16 VNB.t4 2030.77
R247 a_1758_413.t0 a_1758_413.t1 121.952
R248 a_1946_47.t0 a_1946_47.t1 70
R249 SCD.n0 SCD.t0 248.765
R250 SCD.n0 SCD.t1 191.996
R251 SCD SCD.n0 79.072
R252 a_817_66.t1 a_817_66.t0 60
R253 SCE.t2 SCE.t3 729.319
R254 SCE.n0 SCE.t0 273.133
R255 SCE.n1 SCE.t2 215.9
R256 SCE.n1 SCE.n0 145.294
R257 SCE.n0 SCE.t1 138.173
R258 SCE SCE.n1 83.053
R259  SCE 34.974
R260 a_538_389.t0 a_538_389.t1 94.851
R261 RESET_B.n6 RESET_B.t0 2023.69
R262 RESET_B.n2 RESET_B.t2 396.265
R263 RESET_B.n6 RESET_B.t3 205.8
R264 RESET_B.n3 RESET_B.t1 126.39
R265 RESET_B.n3 RESET_B.n2 12.45
R266 RESET_B.n9 RESET_B 11.255
R267 RESET_B.n7 RESET_B.n6 9.81
R268 RESET_B.n4 RESET_B.n3 9.3
R269 RESET_B.n7 RESET_B 5.451
R270 RESET_B.n9 RESET_B.n8 4.659
R271 RESET_B.n5 RESET_B.n4 3.772
R272 RESET_B RESET_B.n9 3.751
R273 RESET_B.n4 RESET_B.n1 3.2
R274 RESET_B.n8 RESET_B.n5 2.364
R275 RESET_B.n8 RESET_B.n7 1.73
R276 RESET_B.n1 RESET_B.n0 0.685
R277 D.n0 D.t0 234.941
R278 D.n0 D.t1 164.248
R279 D.n1 D.n0 76
R280  D.n1 22.551
R281 D.n1 D 5.818
R282 a_569_119.t0 a_569_119.t1 60
R283 a_1187_47.t0 a_1187_47.t1 111.393
R284 Q.n4 Q.n3 143.02
R285 Q.n1 Q.n0 92.5
R286 Q.n2 Q 89.6
R287 Q.n2 Q.n1 64.808
R288 Q.n3 Q.t1 26.595
R289 Q.n3 Q.t0 26.595
R290 Q.n0 Q.t3 24.923
R291 Q.n0 Q.t2 24.923
R292 Q Q.n2 16
R293 Q.n1 Q 10.092
R294 Q.n4 Q 9.022
R295 Q Q.n4 7.342
R296 Q.n2 Q 0.738
R297 a_1293_47.t0 a_1293_47.t1 60
R298 a_1191_413.n0 a_1191_413.t2 738.672
R299 a_1191_413.n0 a_1191_413.t1 63.321
R300 a_1191_413.t0 a_1191_413.n0 63.321
R301 CLK.n0 CLK.t0 428.577
R302 CLK.n0 CLK.t1 426.167
R303 CLK.n1 CLK.n0 76
R304 CLK.n1 CLK 10.422
R305 CLK CLK.n1 2.011
C0 RESET_B VGND 0.35fF
C1 VPWR Q 0.24fF
C2 SCD VGND 0.11fF
C3 VPB VPWR 0.24fF
C4 VGND Q 0.11fF
C5 VPWR VGND 0.11fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__sdfrtp_4.ext - technology: sky130A

.subckt sky130_fd_sc_hd__sdfrtp_4 VPWR VGND SCE SCD D RESET_B CLK Q VNB VPB
X0 a_193_47.t0 a_27_47.t2 VPWR.t1 VPB.t5 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_780_389.t1 a_299_66.t2 a_620_389.t2 VPB.t14 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=540000u l=150000u
X2 a_1245_303.t2 a_1079_413.t4 VPWR.t9 VPB.t13 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X3 VPWR.t6 a_1592_47.t4 a_1767_21.t2 VPB.t10 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 VGND.t8 a_1767_21.t3 a_1701_47.t1 VNB.t13 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 a_1758_413.t0 a_193_47.t2 a_1592_47.t0 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 a_1767_21.t1 a_1592_47.t5 a_1946_47.t1 VNB.t20 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7 VGND.t0 SCD.t0 a_817_66.t0 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=180000u
X8 a_538_389.t0 SCE.t0 VPWR.t13 VPB.t19 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=540000u l=150000u
X9 VPWR.t0 SCD.t1 a_780_389.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=540000u l=150000u
X10 VGND.t7 a_1767_21.t4 Q.t7 VNB.t12 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 VPWR.t14 SCE.t1 a_299_66.t1 VPB.t20 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=540000u l=150000u
X12 a_1767_21.t0 RESET_B.t0 VPWR.t7 VPB.t11 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13 a_193_47.t1 a_27_47.t3 VGND.t1 VNB.t5 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14 a_620_389.t4 D.t0 a_569_119.t1 VNB.t18 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15 a_1187_47.t0 a_193_47.t3 a_1079_413.t1 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X16 VGND.t6 a_1767_21.t5 Q.t6 VNB.t11 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X17 a_1293_47.t0 a_1245_303.t4 a_1187_47.t1 VNB.t6 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18 VPWR.t11 a_1767_21.t6 Q.t3 VPB.t17 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X19 VPWR.t2 a_1245_303.t5 a_1191_413.t1 VPB.t6 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20 a_620_389.t5 D.t1 a_538_389.t1 VPB.t15 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=540000u l=150000u
X21 Q.t5 a_1767_21.t7 VGND.t5 VNB.t10 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X22 a_1191_413.t0 a_27_47.t4 a_1079_413.t3 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23 a_569_119.t0 a_299_66.t3 VGND.t9 VNB.t14 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24 VPWR.t4 a_1767_21.t8 a_1758_413.t1 VPB.t8 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X25 VGND.t2 RESET_B.t1 a_1293_47.t1 VNB.t7 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X26 Q.t2 a_1767_21.t9 VPWR.t5 VPB.t9 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X27 Q.t4 a_1767_21.t10 VGND.t4 VNB.t9 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X28 a_1079_413.t2 a_27_47.t5 a_620_389.t1 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X29 a_1191_413.t2 RESET_B.t2 VPWR.t8 VPB.t12 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X30 VPWR.t3 a_1767_21.t11 Q.t1 VPB.t7 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X31 a_1701_47.t0 a_27_47.t6 a_1592_47.t3 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X32 a_1946_47.t0 RESET_B.t3 VGND.t3 VNB.t8 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X33 a_1592_47.t1 a_193_47.t4 a_1245_303.t0 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X34 Q.t0 a_1767_21.t12 VPWR.t12 VPB.t18 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X35 VGND.t10 SCE.t2 a_299_66.t0 VNB.t15 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X36 a_1592_47.t2 a_27_47.t7 a_1245_303.t1 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X37 a_1245_303.t3 a_1079_413.t5 VGND.t12 VNB.t19 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X38 a_1079_413.t0 a_193_47.t5 a_620_389.t0 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X39 VPWR.t10 CLK.t0 a_27_47.t1 VPB.t16 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X40 a_817_66.t1 SCE.t3 a_620_389.t3 VNB.t16 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=500000u
X41 VGND.t11 CLK.t1 a_27_47.t0 VNB.t17 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
R0 a_27_47.n1 a_27_47.t4 534.047
R1 a_27_47.n0 a_27_47.t7 489.903
R2 a_27_47.n1 a_27_47.t5 276.816
R3 a_27_47.t1 a_27_47.n9 243.743
R4 a_27_47.n7 a_27_47.t2 238.856
R5 a_27_47.n0 a_27_47.t6 204.42
R6 a_27_47.n3 a_27_47.t0 175.866
R7 a_27_47.n5 a_27_47.t3 156.738
R8 a_27_47.n2 a_27_47.n0 14.808
R9 a_27_47.n6 a_27_47.n5 12.496
R10 a_27_47.n2 a_27_47.n1 11.633
R11 a_27_47.n8 a_27_47.n7 9.3
R12 a_27_47.n9 a_27_47.n2 6.029
R13 a_27_47.n4 a_27_47.n3 2.844
R14 a_27_47.n7 a_27_47.n6 2.677
R15 a_27_47.n9 a_27_47.n8 1.13
R16 a_27_47.n8 a_27_47.n4 0.609
R17 VPWR.n20 VPWR.t9 514.01
R18 VPWR.n36 VPWR.t0 408.48
R19 VPWR.n7 VPWR.t6 370.56
R20 VPWR.n45 VPWR.n44 323.37
R21 VPWR.n55 VPWR.n54 311.893
R22 VPWR.n12 VPWR.n11 310.932
R23 VPWR.n25 VPWR.n24 292.5
R24 VPWR.n2 VPWR.t3 156.581
R25 VPWR.n5 VPWR.t5 152.716
R26 VPWR.n1 VPWR.n0 126.121
R27 VPWR.n11 VPWR.t4 114.916
R28 VPWR.n24 VPWR.t8 103.19
R29 VPWR.n24 VPWR.t2 93.809
R30 VPWR.n11 VPWR.t7 63.321
R31 VPWR.n44 VPWR.t13 49.25
R32 VPWR.n44 VPWR.t14 49.25
R33 VPWR.n54 VPWR.t10 29.55
R34 VPWR.n0 VPWR.t11 28.565
R35 VPWR.n0 VPWR.t12 26.595
R36 VPWR.n54 VPWR.t1 26.595
R37 VPWR.n46 VPWR.n45 9.411
R38 VPWR.n4 VPWR.n3 4.65
R39 VPWR.n6 VPWR.n5 4.65
R40 VPWR.n8 VPWR.n7 4.65
R41 VPWR.n10 VPWR.n9 4.65
R42 VPWR.n13 VPWR.n12 4.65
R43 VPWR.n15 VPWR.n14 4.65
R44 VPWR.n17 VPWR.n16 4.65
R45 VPWR.n19 VPWR.n18 4.65
R46 VPWR.n21 VPWR.n20 4.65
R47 VPWR.n23 VPWR.n22 4.65
R48 VPWR.n27 VPWR.n26 4.65
R49 VPWR.n29 VPWR.n28 4.65
R50 VPWR.n31 VPWR.n30 4.65
R51 VPWR.n33 VPWR.n32 4.65
R52 VPWR.n35 VPWR.n34 4.65
R53 VPWR.n37 VPWR.n36 4.65
R54 VPWR.n39 VPWR.n38 4.65
R55 VPWR.n41 VPWR.n40 4.65
R56 VPWR.n43 VPWR.n42 4.65
R57 VPWR.n47 VPWR.n46 4.65
R58 VPWR.n49 VPWR.n48 4.65
R59 VPWR.n51 VPWR.n50 4.65
R60 VPWR.n53 VPWR.n52 4.65
R61 VPWR.n56 VPWR.n55 3.958
R62 VPWR.n2 VPWR.n1 3.933
R63 VPWR.n26 VPWR.n25 2.702
R64 VPWR.n4 VPWR.n2 0.244
R65 VPWR.n56 VPWR.n53 0.137
R66 VPWR VPWR.n56 0.121
R67 VPWR.n6 VPWR.n4 0.119
R68 VPWR.n8 VPWR.n6 0.119
R69 VPWR.n10 VPWR.n8 0.119
R70 VPWR.n13 VPWR.n10 0.119
R71 VPWR.n15 VPWR.n13 0.119
R72 VPWR.n17 VPWR.n15 0.119
R73 VPWR.n19 VPWR.n17 0.119
R74 VPWR.n21 VPWR.n19 0.119
R75 VPWR.n23 VPWR.n21 0.119
R76 VPWR.n27 VPWR.n23 0.119
R77 VPWR.n29 VPWR.n27 0.119
R78 VPWR.n31 VPWR.n29 0.119
R79 VPWR.n33 VPWR.n31 0.119
R80 VPWR.n35 VPWR.n33 0.119
R81 VPWR.n37 VPWR.n35 0.119
R82 VPWR.n39 VPWR.n37 0.119
R83 VPWR.n41 VPWR.n39 0.119
R84 VPWR.n43 VPWR.n41 0.119
R85 VPWR.n47 VPWR.n43 0.119
R86 VPWR.n49 VPWR.n47 0.119
R87 VPWR.n51 VPWR.n49 0.119
R88 VPWR.n53 VPWR.n51 0.119
R89 a_193_47.n1 a_193_47.t4 266.53
R90 a_193_47.n0 a_193_47.t3 265.71
R91 a_193_47.n1 a_193_47.t2 231.814
R92 a_193_47.n3 a_193_47.t1 210.139
R93 a_193_47.n0 a_193_47.t5 146.401
R94 a_193_47.t0 a_193_47.n3 38.199
R95 a_193_47.n2 a_193_47.n1 7.332
R96 a_193_47.n3 a_193_47.n2 6.062
R97 a_193_47.n2 a_193_47.n0 3.302
R98 VPB.t5 VPB.t20 774.312
R99 VPB.t0 VPB.t1 637.547
R100 VPB.t10 VPB.t9 556.386
R101 VPB.t12 VPB.t13 556.386
R102 VPB.t15 VPB.t14 511.784
R103 VPB.t6 VPB.t12 337.383
R104 VPB.t1 VPB.t4 331.464
R105 VPB.t8 VPB.t11 313.707
R106 VPB.t13 VPB.t3 281.152
R107 VPB.t14 VPB.t0 275.084
R108 VPB.t20 VPB.t19 268.686
R109 VPB.t19 VPB.t15 262.289
R110 VPB.t16 VPB.t5 257.476
R111 VPB.t17 VPB.t18 254.517
R112 VPB.t3 VPB.t2 254.517
R113 VPB.t18 VPB.t7 248.598
R114 VPB.t9 VPB.t17 248.598
R115 VPB.t11 VPB.t10 248.598
R116 VPB.t4 VPB.t6 248.598
R117 VPB.t2 VPB.t8 242.679
R118 VPB VPB.t16 177.57
R119 a_299_66.n0 a_299_66.t2 1032.99
R120 a_299_66.t1 a_299_66.n0 408.174
R121 a_299_66.n0 a_299_66.t3 270.218
R122 a_299_66.n0 a_299_66.t0 195.971
R123 a_620_389.n0 a_620_389.t0 393.588
R124 a_620_389.n3 a_620_389.n2 307.182
R125 a_620_389.n0 a_620_389.t1 267.547
R126 a_620_389.n2 a_620_389.n1 184.051
R127 a_620_389.n3 a_620_389.t5 162.342
R128 a_620_389.n1 a_620_389.t3 106.635
R129 a_620_389.n2 a_620_389.n0 83.2
R130 a_620_389.t2 a_620_389.n3 74.787
R131 a_620_389.n1 a_620_389.t4 38.572
R132 a_780_389.t0 a_780_389.t1 102.148
R133 a_1079_413.n3 a_1079_413.n2 393.455
R134 a_1079_413.n1 a_1079_413.t4 339.006
R135 a_1079_413.n2 a_1079_413.n0 193.393
R136 a_1079_413.n1 a_1079_413.t5 168.699
R137 a_1079_413.n2 a_1079_413.n1 157.693
R138 a_1079_413.t0 a_1079_413.n3 128.988
R139 a_1079_413.n0 a_1079_413.t2 71.666
R140 a_1079_413.n3 a_1079_413.t3 63.321
R141 a_1079_413.n0 a_1079_413.t1 45
R142 a_1245_303.n0 a_1245_303.t4 365.917
R143 a_1245_303.n3 a_1245_303.n2 352.126
R144 a_1245_303.n2 a_1245_303.n1 177.291
R145 a_1245_303.n0 a_1245_303.t5 158.39
R146 a_1245_303.n2 a_1245_303.n0 151.67
R147 a_1245_303.n3 a_1245_303.t1 72.702
R148 a_1245_303.n1 a_1245_303.t0 63.333
R149 a_1245_303.t2 a_1245_303.n3 50.422
R150 a_1245_303.n1 a_1245_303.t3 26.77
R151 a_1592_47.n1 a_1592_47.t5 1025.84
R152 a_1592_47.n1 a_1592_47.t4 412.282
R153 a_1592_47.n3 a_1592_47.n2 342.717
R154 a_1592_47.n2 a_1592_47.n0 210.387
R155 a_1592_47.n2 a_1592_47.n1 144.894
R156 a_1592_47.n0 a_1592_47.t1 70
R157 a_1592_47.n3 a_1592_47.t2 68.011
R158 a_1592_47.t0 a_1592_47.n3 63.321
R159 a_1592_47.n0 a_1592_47.t3 61.666
R160 a_1767_21.n4 a_1767_21.t8 1015.03
R161 a_1767_21.n7 a_1767_21.n6 491.4
R162 a_1767_21.n0 a_1767_21.t11 212.079
R163 a_1767_21.n1 a_1767_21.t12 212.079
R164 a_1767_21.n2 a_1767_21.t6 212.079
R165 a_1767_21.n3 a_1767_21.t9 212.079
R166 a_1767_21.n5 a_1767_21.n4 181.032
R167 a_1767_21.n4 a_1767_21.t3 178.584
R168 a_1767_21.n0 a_1767_21.t4 139.779
R169 a_1767_21.n1 a_1767_21.t7 139.779
R170 a_1767_21.n2 a_1767_21.t5 139.779
R171 a_1767_21.n3 a_1767_21.t10 139.779
R172 a_1767_21.n5 a_1767_21.t1 131.071
R173 a_1767_21.n6 a_1767_21.n3 97.924
R174 a_1767_21.n6 a_1767_21.n5 64.011
R175 a_1767_21.n7 a_1767_21.t2 63.321
R176 a_1767_21.t0 a_1767_21.n7 63.321
R177 a_1767_21.n2 a_1767_21.n1 62.806
R178 a_1767_21.n1 a_1767_21.n0 61.345
R179 a_1767_21.n3 a_1767_21.n2 61.345
R180 a_1701_47.t1 a_1701_47.t0 93.516
R181 VGND.n2 VGND.t7 207.936
R182 VGND.n5 VGND.t4 197.787
R183 VGND.n46 VGND.t9 159.774
R184 VGND.n48 VGND.t10 149.495
R185 VGND.n35 VGND.t0 148.719
R186 VGND.n14 VGND.t3 117.142
R187 VGND.n1 VGND.n0 114.711
R188 VGND.n15 VGND.n14 113.205
R189 VGND.n25 VGND.n24 107.239
R190 VGND.n55 VGND.n54 107.239
R191 VGND.n24 VGND.t2 72.857
R192 VGND.n24 VGND.t12 60.579
R193 VGND.n14 VGND.t8 52.857
R194 VGND.n0 VGND.t6 26.769
R195 VGND.n0 VGND.t5 24.923
R196 VGND.n54 VGND.t1 24.923
R197 VGND.n54 VGND.t11 24.923
R198 VGND.n16 VGND.n15 15.058
R199 VGND.n2 VGND.n1 9.603
R200 VGND.n4 VGND.n3 4.65
R201 VGND.n7 VGND.n6 4.65
R202 VGND.n9 VGND.n8 4.65
R203 VGND.n11 VGND.n10 4.65
R204 VGND.n13 VGND.n12 4.65
R205 VGND.n17 VGND.n16 4.65
R206 VGND.n19 VGND.n18 4.65
R207 VGND.n21 VGND.n20 4.65
R208 VGND.n23 VGND.n22 4.65
R209 VGND.n26 VGND.n25 4.65
R210 VGND.n28 VGND.n27 4.65
R211 VGND.n30 VGND.n29 4.65
R212 VGND.n32 VGND.n31 4.65
R213 VGND.n34 VGND.n33 4.65
R214 VGND.n37 VGND.n36 4.65
R215 VGND.n39 VGND.n38 4.65
R216 VGND.n41 VGND.n40 4.65
R217 VGND.n43 VGND.n42 4.65
R218 VGND.n45 VGND.n44 4.65
R219 VGND.n47 VGND.n46 4.65
R220 VGND.n49 VGND.n48 4.65
R221 VGND.n51 VGND.n50 4.65
R222 VGND.n53 VGND.n52 4.65
R223 VGND.n36 VGND.n35 4.141
R224 VGND.n56 VGND.n55 3.932
R225 VGND.n6 VGND.n5 0.376
R226 VGND.n4 VGND.n2 0.317
R227 VGND.n56 VGND.n53 0.137
R228 VGND.n7 VGND.n4 0.119
R229 VGND.n9 VGND.n7 0.119
R230 VGND.n11 VGND.n9 0.119
R231 VGND.n13 VGND.n11 0.119
R232 VGND.n17 VGND.n13 0.119
R233 VGND.n19 VGND.n17 0.119
R234 VGND.n21 VGND.n19 0.119
R235 VGND.n23 VGND.n21 0.119
R236 VGND.n26 VGND.n23 0.119
R237 VGND.n28 VGND.n26 0.119
R238 VGND.n30 VGND.n28 0.119
R239 VGND.n32 VGND.n30 0.119
R240 VGND.n34 VGND.n32 0.119
R241 VGND.n37 VGND.n34 0.119
R242 VGND.n39 VGND.n37 0.119
R243 VGND.n41 VGND.n39 0.119
R244 VGND.n43 VGND.n41 0.119
R245 VGND.n45 VGND.n43 0.119
R246 VGND.n47 VGND.n45 0.119
R247 VGND.n49 VGND.n47 0.119
R248 VGND.n51 VGND.n49 0.119
R249 VGND.n53 VGND.n51 0.119
R250 VGND VGND.n56 0.11
R251 VNB VNB.t17 26484.6
R252 VNB.t0 VNB.t4 6619.1
R253 VNB.t15 VNB.t14 6123.67
R254 VNB.t20 VNB.t9 5483.65
R255 VNB.t5 VNB.t15 5321.88
R256 VNB.t13 VNB.t8 4820.59
R257 VNB.t16 VNB.t0 3558.82
R258 VNB.t7 VNB.t19 3550.91
R259 VNB.t4 VNB.t2 3548.39
R260 VNB.t1 VNB.t3 3526.47
R261 VNB.t2 VNB.t6 3476.38
R262 VNB.t3 VNB.t13 3105.88
R263 VNB.t18 VNB.t16 2863.63
R264 VNB.t8 VNB.t20 2555.88
R265 VNB.t6 VNB.t7 2329.41
R266 VNB.t14 VNB.t18 2329.41
R267 VNB.t19 VNB.t1 2280.14
R268 VNB.t11 VNB.t10 2079.12
R269 VNB.t10 VNB.t12 2030.77
R270 VNB.t9 VNB.t11 2030.77
R271 VNB.t17 VNB.t5 2030.77
R272 a_1758_413.t0 a_1758_413.t1 121.952
R273 a_1946_47.t0 a_1946_47.t1 70
R274 SCD.n0 SCD.t0 248.765
R275 SCD.n0 SCD.t1 191.996
R276 SCD SCD.n0 79.072
R277 a_817_66.t0 a_817_66.t1 60
R278 SCE.t2 SCE.t3 729.319
R279 SCE.n0 SCE.t0 273.133
R280 SCE.n1 SCE.t2 215.9
R281 SCE.n1 SCE.n0 145.294
R282 SCE.n0 SCE.t1 138.173
R283 SCE SCE.n1 83.053
R284  SCE 34.974
R285 a_538_389.t0 a_538_389.t1 94.851
R286 Q.n4 Q.n2 175.821
R287 Q.n8 Q.n7 143.02
R288 Q.n4 Q.n3 111.188
R289 Q.n1 Q.n0 92.5
R290 Q.n6 Q 89.6
R291 Q.n5 Q.n4 31.806
R292 Q.n7 Q.t3 26.595
R293 Q.n7 Q.t2 26.595
R294 Q.n2 Q.t1 26.595
R295 Q.n2 Q.t0 26.595
R296 Q.n0 Q.t6 24.923
R297 Q.n0 Q.t4 24.923
R298 Q.n3 Q.t7 24.923
R299 Q.n3 Q.t5 24.923
R300 Q.n6 Q.n5 24.38
R301 Q.n5 Q.n1 20.313
R302 Q Q.n6 16
R303 Q.n1 Q 10.092
R304 Q.n8 Q 9.022
R305 Q Q.n8 7.342
R306 Q.n6 Q 0.738
R307 RESET_B.n6 RESET_B.t0 2023.69
R308 RESET_B.n2 RESET_B.t2 396.265
R309 RESET_B.n6 RESET_B.t3 205.8
R310 RESET_B.n3 RESET_B.t1 126.39
R311 RESET_B.n3 RESET_B.n2 12.45
R312 RESET_B.n9 RESET_B 11.255
R313 RESET_B.n7 RESET_B.n6 9.81
R314 RESET_B.n4 RESET_B.n3 9.3
R315 RESET_B.n7 RESET_B 5.451
R316 RESET_B.n9 RESET_B.n8 4.659
R317 RESET_B.n5 RESET_B.n4 3.772
R318 RESET_B RESET_B.n9 3.751
R319 RESET_B.n4 RESET_B.n1 3.2
R320 RESET_B.n8 RESET_B.n5 2.364
R321 RESET_B.n8 RESET_B.n7 1.73
R322 RESET_B.n1 RESET_B.n0 0.685
R323 D.n0 D.t0 234.941
R324 D.n0 D.t1 164.248
R325 D.n1 D.n0 76
R326  D.n1 22.551
R327 D.n1 D 5.818
R328 a_569_119.t0 a_569_119.t1 60
R329 a_1187_47.t1 a_1187_47.t0 111.393
R330 a_1293_47.t0 a_1293_47.t1 60
R331 a_1191_413.n0 a_1191_413.t2 738.672
R332 a_1191_413.n0 a_1191_413.t1 63.321
R333 a_1191_413.t0 a_1191_413.n0 63.321
R334 CLK.n0 CLK.t0 428.577
R335 CLK.n0 CLK.t1 426.167
R336 CLK.n1 CLK.n0 76
R337 CLK.n1 CLK 10.422
R338 CLK CLK.n1 2.011
C0 VGND Q 0.25fF
C1 VPWR VGND 0.13fF
C2 RESET_B VGND 0.35fF
C3 VPWR Q 0.55fF
C4 SCD VGND 0.11fF
C5 VPB VPWR 0.26fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__sdfsbp_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__sdfsbp_1 SCD CLK Q_N D SET_B SCE Q VPWR VGND VNB VPB
X0 Q.t1 a_2412_47.t2 VGND.t12 VNB.t20 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 a_1129_21.t2 a_997_413.t4 VPWR.t14 VPB.t20 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 VPWR.t2 SCD.t0 a_27_369.t1 VPB.t5 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X3 a_1081_413.t0 a_643_369.t2 a_997_413.t2 VPB.t6 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 a_1587_329.t4 SET_B.t0 VPWR.t8 VPB.t12 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 a_809_369.t1 a_643_369.t3 VGND.t2 VNB.t6 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 a_997_413.t0 a_809_369.t2 a_181_47.t5 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7 a_1347_47.t1 a_997_413.t5 a_1129_21.t1 VNB.t15 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 VPWR.t4 a_1129_21.t3 a_1081_413.t1 VPB.t16 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9 a_1770_295.t0 a_1587_329.t5 VPWR.t5 VPB.t9 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10 Q_N.t0 a_1587_329.t6 VPWR.t6 VPB.t10 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 a_1807_47.t0 a_643_369.t4 a_1587_329.t0 VNB.t7 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12 VPWR.t9 SET_B.t1 a_1129_21.t0 VPB.t13 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13 Q_N.t1 a_1587_329.t7 VGND.t4 VNB.t10 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14 a_181_47.t3 SCE.t0 a_109_47.t1 VNB.t18 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15 a_1514_47.t1 a_997_413.t6 VGND.t9 VNB.t16 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X16 a_1587_329.t2 a_809_369.t3 a_1514_47.t0 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X17 VPWR.t1 a_1770_295.t2 a_1712_413.t0 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18 VGND.t7 SET_B.t2 a_1347_47.t0 VNB.t13 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19 Q.t0 a_2412_47.t3 VPWR.t12 VPB.t18 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X20 a_1879_47.t0 a_1770_295.t3 a_1807_47.t1 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21 a_27_369.t0 a_319_21.t2 a_181_47.t4 VPB.t15 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X22 VGND.t11 SCE.t1 a_319_21.t1 VNB.t19 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23 a_181_47.t1 D.t0 a_193_369.t1 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X24 a_265_47.t0 D.t1 a_181_47.t2 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X25 a_997_413.t3 a_643_369.t5 a_181_47.t0 VNB.t8 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X26 VGND.t5 a_1587_329.t8 a_2412_47.t0 VNB.t11 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X27 a_1087_47.t0 a_809_369.t4 a_997_413.t1 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X28 a_193_369.t0 SCE.t2 VPWR.t10 VPB.t14 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X29 a_809_369.t0 a_643_369.t6 VPWR.t3 VPB.t7 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X30 VPWR.t0 SCE.t3 a_319_21.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X31 VGND.t8 SET_B.t3 a_1879_47.t1 VNB.t14 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X32 VPWR.t7 a_1587_329.t9 a_2412_47.t1 VPB.t11 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X33 VPWR.t11 CLK.t0 a_643_369.t1 VPB.t17 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X34 a_1514_329.t1 a_997_413.t7 VPWR.t13 VPB.t19 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X35 a_1587_329.t1 a_643_369.t7 a_1514_329.t0 VPB.t8 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X36 a_1712_413.t1 a_809_369.t5 a_1587_329.t3 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X37 VGND.t1 a_319_21.t3 a_265_47.t1 VNB.t5 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X38 VGND.t3 a_1129_21.t4 a_1087_47.t1 VNB.t9 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X39 VGND.t10 CLK.t1 a_643_369.t0 VNB.t17 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X40 a_1770_295.t1 a_1587_329.t10 VGND.t6 VNB.t12 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X41 a_109_47.t0 SCD.t1 VGND.t0 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
R0 a_2412_47.t1 a_2412_47.n1 252.48
R1 a_2412_47.n0 a_2412_47.t3 241.534
R2 a_2412_47.n0 a_2412_47.t2 169.234
R3 a_2412_47.n1 a_2412_47.t0 164.899
R4 a_2412_47.n1 a_2412_47.n0 101.212
R5 VGND.n47 VGND.t1 166.664
R6 VGND.n43 VGND.t11 145.376
R7 VGND.n56 VGND.t0 145.005
R8 VGND.n29 VGND.t3 131.071
R9 VGND.n2 VGND.n0 123.241
R10 VGND.n1 VGND.t4 113.732
R11 VGND.n6 VGND.n5 113.205
R12 VGND.n39 VGND.n38 107.364
R13 VGND.n22 VGND.n21 92.5
R14 VGND.n5 VGND.t8 77.142
R15 VGND.n0 VGND.t5 54.285
R16 VGND.n21 VGND.t9 42.008
R17 VGND.n21 VGND.t7 38.571
R18 VGND.n5 VGND.t6 38.571
R19 VGND.n38 VGND.t2 38.571
R20 VGND.n38 VGND.t10 38.571
R21 VGND.n0 VGND.t12 25.934
R22 VGND.n48 VGND.n47 4.894
R23 VGND.n57 VGND.n56 4.65
R24 VGND.n4 VGND.n3 4.65
R25 VGND.n8 VGND.n7 4.65
R26 VGND.n10 VGND.n9 4.65
R27 VGND.n12 VGND.n11 4.65
R28 VGND.n14 VGND.n13 4.65
R29 VGND.n16 VGND.n15 4.65
R30 VGND.n18 VGND.n17 4.65
R31 VGND.n20 VGND.n19 4.65
R32 VGND.n24 VGND.n23 4.65
R33 VGND.n26 VGND.n25 4.65
R34 VGND.n28 VGND.n27 4.65
R35 VGND.n31 VGND.n30 4.65
R36 VGND.n33 VGND.n32 4.65
R37 VGND.n35 VGND.n34 4.65
R38 VGND.n37 VGND.n36 4.65
R39 VGND.n40 VGND.n39 4.65
R40 VGND.n42 VGND.n41 4.65
R41 VGND.n44 VGND.n43 4.65
R42 VGND.n46 VGND.n45 4.65
R43 VGND.n49 VGND.n48 4.65
R44 VGND.n51 VGND.n50 4.65
R45 VGND.n53 VGND.n52 4.65
R46 VGND.n55 VGND.n54 4.65
R47 VGND.n30 VGND.n29 4.189
R48 VGND.n2 VGND.n1 4.074
R49 VGND.n7 VGND.n6 3.388
R50 VGND.n23 VGND.n22 1.438
R51 VGND.n4 VGND.n2 0.142
R52 VGND.n8 VGND.n4 0.119
R53 VGND.n10 VGND.n8 0.119
R54 VGND.n12 VGND.n10 0.119
R55 VGND.n14 VGND.n12 0.119
R56 VGND.n16 VGND.n14 0.119
R57 VGND.n18 VGND.n16 0.119
R58 VGND.n20 VGND.n18 0.119
R59 VGND.n24 VGND.n20 0.119
R60 VGND.n26 VGND.n24 0.119
R61 VGND.n28 VGND.n26 0.119
R62 VGND.n31 VGND.n28 0.119
R63 VGND.n33 VGND.n31 0.119
R64 VGND.n35 VGND.n33 0.119
R65 VGND.n37 VGND.n35 0.119
R66 VGND.n40 VGND.n37 0.119
R67 VGND.n42 VGND.n40 0.119
R68 VGND.n44 VGND.n42 0.119
R69 VGND.n46 VGND.n44 0.119
R70 VGND.n49 VGND.n46 0.119
R71 VGND.n51 VGND.n49 0.119
R72 VGND.n53 VGND.n51 0.119
R73 VGND.n55 VGND.n53 0.119
R74 VGND.n57 VGND.n55 0.119
R75 VGND VGND.n57 0.02
R76 Q.n2 Q.n1 292.5
R77 Q.n1 Q.n0 147.08
R78 Q.n5 Q.t1 82.802
R79 Q.n1 Q.t0 26.595
R80 Q.n4 Q 19.372
R81 Q.n0 Q 10.397
R82 Q Q.n5 6.811
R83 Q.n3 Q.n2 6.211
R84 Q.n5 Q 5.593
R85 Q.n2 Q 4.705
R86 Q.n4 Q 4.151
R87 Q Q.n3 3.459
R88 Q.n0 Q 2.366
R89 Q Q.n4 2.258
R90 Q.n3 Q 1.882
R91 VNB VNB.t2 6438.23
R92 VNB.t5 VNB.t19 6276.47
R93 VNB.t9 VNB.t15 6082.35
R94 VNB.t6 VNB.t8 6082.35
R95 VNB.t19 VNB.t17 6082.35
R96 VNB.t12 VNB.t10 5321.88
R97 VNB.t10 VNB.t11 4545.05
R98 VNB.t3 VNB.t14 4141.18
R99 VNB.t16 VNB.t0 4131.11
R100 VNB.t14 VNB.t12 3591.18
R101 VNB.t0 VNB.t7 3292.09
R102 VNB.t8 VNB.t1 2717.65
R103 VNB.t17 VNB.t6 2717.65
R104 VNB.t4 VNB.t5 2717.65
R105 VNB.t18 VNB.t4 2717.65
R106 VNB.t7 VNB.t3 2329.41
R107 VNB.t15 VNB.t13 2329.41
R108 VNB.t1 VNB.t9 2329.41
R109 VNB.t2 VNB.t18 2329.41
R110 VNB.t11 VNB.t20 2296.7
R111 VNB.t13 VNB.t16 2280.14
R112 a_997_413.n1 a_997_413.t4 583.073
R113 a_997_413.n5 a_997_413.n4 369.55
R114 a_997_413.n0 a_997_413.t7 267.241
R115 a_997_413.n1 a_997_413.t5 251.077
R116 a_997_413.n0 a_997_413.t6 170.841
R117 a_997_413.n4 a_997_413.n3 141.906
R118 a_997_413.n2 a_997_413.n0 120.616
R119 a_997_413.n2 a_997_413.n1 76
R120 a_997_413.n5 a_997_413.t2 63.321
R121 a_997_413.t0 a_997_413.n5 63.321
R122 a_997_413.n4 a_997_413.n2 46.717
R123 a_997_413.n3 a_997_413.t1 38.571
R124 a_997_413.n3 a_997_413.t3 38.571
R125 VPWR.n42 VPWR.t0 439.401
R126 VPWR.n5 VPWR.t5 370.56
R127 VPWR.n53 VPWR.n52 310.932
R128 VPWR.n10 VPWR.n9 306.463
R129 VPWR.n27 VPWR.n26 306.463
R130 VPWR.n38 VPWR.n37 306.463
R131 VPWR.n21 VPWR.n20 292.5
R132 VPWR.n2 VPWR.n0 186.79
R133 VPWR.n9 VPWR.t1 168.857
R134 VPWR.n1 VPWR.t6 158.058
R135 VPWR.n26 VPWR.t14 114.916
R136 VPWR.n26 VPWR.t4 91.464
R137 VPWR.n20 VPWR.t13 87.945
R138 VPWR.n20 VPWR.t9 84.428
R139 VPWR.n9 VPWR.t8 63.321
R140 VPWR.n0 VPWR.t7 58.484
R141 VPWR.n37 VPWR.t3 41.554
R142 VPWR.n37 VPWR.t11 41.554
R143 VPWR.n52 VPWR.t10 41.554
R144 VPWR.n52 VPWR.t2 41.554
R145 VPWR.n0 VPWR.t12 31.662
R146 VPWR.n4 VPWR.n3 4.65
R147 VPWR.n6 VPWR.n5 4.65
R148 VPWR.n8 VPWR.n7 4.65
R149 VPWR.n11 VPWR.n10 4.65
R150 VPWR.n13 VPWR.n12 4.65
R151 VPWR.n15 VPWR.n14 4.65
R152 VPWR.n17 VPWR.n16 4.65
R153 VPWR.n19 VPWR.n18 4.65
R154 VPWR.n23 VPWR.n22 4.65
R155 VPWR.n25 VPWR.n24 4.65
R156 VPWR.n28 VPWR.n27 4.65
R157 VPWR.n30 VPWR.n29 4.65
R158 VPWR.n32 VPWR.n31 4.65
R159 VPWR.n34 VPWR.n33 4.65
R160 VPWR.n36 VPWR.n35 4.65
R161 VPWR.n39 VPWR.n38 4.65
R162 VPWR.n41 VPWR.n40 4.65
R163 VPWR.n43 VPWR.n42 4.65
R164 VPWR.n45 VPWR.n44 4.65
R165 VPWR.n47 VPWR.n46 4.65
R166 VPWR.n49 VPWR.n48 4.65
R167 VPWR.n51 VPWR.n50 4.65
R168 VPWR.n2 VPWR.n1 4.075
R169 VPWR.n54 VPWR.n53 3.932
R170 VPWR.n22 VPWR.n21 0.752
R171 VPWR.n4 VPWR.n2 0.141
R172 VPWR.n54 VPWR.n51 0.137
R173 VPWR VPWR.n54 0.121
R174 VPWR.n6 VPWR.n4 0.119
R175 VPWR.n8 VPWR.n6 0.119
R176 VPWR.n11 VPWR.n8 0.119
R177 VPWR.n13 VPWR.n11 0.119
R178 VPWR.n15 VPWR.n13 0.119
R179 VPWR.n17 VPWR.n15 0.119
R180 VPWR.n19 VPWR.n17 0.119
R181 VPWR.n23 VPWR.n19 0.119
R182 VPWR.n25 VPWR.n23 0.119
R183 VPWR.n28 VPWR.n25 0.119
R184 VPWR.n30 VPWR.n28 0.119
R185 VPWR.n32 VPWR.n30 0.119
R186 VPWR.n34 VPWR.n32 0.119
R187 VPWR.n36 VPWR.n34 0.119
R188 VPWR.n39 VPWR.n36 0.119
R189 VPWR.n41 VPWR.n39 0.119
R190 VPWR.n43 VPWR.n41 0.119
R191 VPWR.n45 VPWR.n43 0.119
R192 VPWR.n47 VPWR.n45 0.119
R193 VPWR.n49 VPWR.n47 0.119
R194 VPWR.n51 VPWR.n49 0.119
R195 a_1129_21.n2 a_1129_21.n1 439.616
R196 a_1129_21.n0 a_1129_21.t1 247.361
R197 a_1129_21.n1 a_1129_21.n0 204.526
R198 a_1129_21.n1 a_1129_21.t3 139.821
R199 a_1129_21.n0 a_1129_21.t4 132.184
R200 a_1129_21.t0 a_1129_21.n2 84.428
R201 a_1129_21.n2 a_1129_21.t2 72.702
R202 VPB.t9 VPB.t10 559.345
R203 VPB.t10 VPB.t11 556.386
R204 VPB.t12 VPB.t9 556.386
R205 VPB.t7 VPB.t3 556.386
R206 VPB.t0 VPB.t17 556.386
R207 VPB.t15 VPB.t0 556.386
R208 VPB.t2 VPB.t12 381.775
R209 VPB.t8 VPB.t4 369.937
R210 VPB.t16 VPB.t20 349.221
R211 VPB.t13 VPB.t19 343.302
R212 VPB.t6 VPB.t16 301.869
R213 VPB.t20 VPB.t13 287.071
R214 VPB.t11 VPB.t18 281.152
R215 VPB.t4 VPB.t2 260.436
R216 VPB.t3 VPB.t6 248.598
R217 VPB.t17 VPB.t7 248.598
R218 VPB.t1 VPB.t15 248.598
R219 VPB.t5 VPB.t14 248.598
R220 VPB.t19 VPB.t8 216.043
R221 VPB.t14 VPB.t1 213.084
R222 VPB VPB.t5 189.408
R223 SCD.n0 SCD.t0 297.824
R224 SCD.n0 SCD.t1 204.638
R225 SCD.n1 SCD.n0 76
R226 SCD.n1 SCD 19.446
R227 SCD SCD.n1 14.03
R228 a_27_369.t0 a_27_369.t1 883.532
R229 a_643_369.n2 a_643_369.t5 393.633
R230 a_643_369.t1 a_643_369.n5 377.577
R231 a_643_369.n0 a_643_369.t4 348.718
R232 a_643_369.n0 a_643_369.t7 343.241
R233 a_643_369.n3 a_643_369.t6 267.297
R234 a_643_369.n4 a_643_369.t0 199.461
R235 a_643_369.n1 a_643_369.t2 147.521
R236 a_643_369.n3 a_643_369.n2 100.205
R237 a_643_369.n2 a_643_369.t3 91.58
R238 a_643_369.n4 a_643_369.n3 76
R239 a_643_369.n1 a_643_369.n0 37.716
R240 a_643_369.n5 a_643_369.n4 30.03
R241 a_643_369.n5 a_643_369.n1 6.022
R242 a_1081_413.t0 a_1081_413.t1 168.857
R243 SET_B.n0 SET_B.t3 350.788
R244 SET_B.n1 SET_B.t2 340.969
R245 SET_B.n0 SET_B.t0 209.401
R246 SET_B.n1 SET_B.t1 177.067
R247 SET_B.n2 SET_B.n0 140.657
R248 SET_B.n2 SET_B.n1 7.848
R249 SET_B SET_B.n2 3.774
R250 a_1587_329.n7 a_1587_329.n6 384.902
R251 a_1587_329.n6 a_1587_329.t4 373.979
R252 a_1587_329.n3 a_1587_329.n2 334.522
R253 a_1587_329.n0 a_1587_329.t9 247.426
R254 a_1587_329.n1 a_1587_329.t6 212.079
R255 a_1587_329.n0 a_1587_329.t8 176.733
R256 a_1587_329.n5 a_1587_329.t5 154.759
R257 a_1587_329.n1 a_1587_329.t7 139.779
R258 a_1587_329.n1 a_1587_329.n0 137.296
R259 a_1587_329.n4 a_1587_329.n1 126.342
R260 a_1587_329.n3 a_1587_329.t10 125.878
R261 a_1587_329.n6 a_1587_329.n5 118.095
R262 a_1587_329.t1 a_1587_329.n7 102.017
R263 a_1587_329.n7 a_1587_329.t3 91.464
R264 a_1587_329.n2 a_1587_329.t0 88.571
R265 a_1587_329.n5 a_1587_329.n4 74.796
R266 a_1587_329.n2 a_1587_329.t2 33.437
R267 a_1587_329.n4 a_1587_329.n3 32.133
R268 a_809_369.n2 a_809_369.t4 433.507
R269 a_809_369.n0 a_809_369.t3 383.456
R270 a_809_369.t0 a_809_369.n3 380.975
R271 a_809_369.n2 a_809_369.t2 321.333
R272 a_809_369.n1 a_809_369.t1 182.04
R273 a_809_369.n0 a_809_369.t5 148.348
R274 a_809_369.n1 a_809_369.n0 116.617
R275 a_809_369.n3 a_809_369.n2 38.615
R276 a_809_369.n3 a_809_369.n1 1.197
R277 a_181_47.n0 a_181_47.t5 399.999
R278 a_181_47.n3 a_181_47.n2 324.146
R279 a_181_47.n2 a_181_47.n1 322.769
R280 a_181_47.n0 a_181_47.t0 196.303
R281 a_181_47.n3 a_181_47.t4 41.554
R282 a_181_47.t1 a_181_47.n3 41.554
R283 a_181_47.n1 a_181_47.t2 38.571
R284 a_181_47.n1 a_181_47.t3 38.571
R285 a_181_47.n2 a_181_47.n0 13.323
R286 a_1347_47.t0 a_1347_47.t1 60
R287 a_1770_295.n0 a_1770_295.t2 458.433
R288 a_1770_295.t0 a_1770_295.n1 405.79
R289 a_1770_295.n1 a_1770_295.t1 185.706
R290 a_1770_295.n1 a_1770_295.n0 182.379
R291 a_1770_295.n0 a_1770_295.t3 161.201
R292 Q_N.n2 Q_N.n1 292.5
R293 Q_N.n1 Q_N.n0 147.009
R294 Q_N.n3 Q_N.t1 83.064
R295 Q_N.n1 Q_N.t0 26.595
R296 Q_N.n0 Q_N 10.611
R297 Q_N Q_N.n2 8.145
R298 Q_N.n3 Q_N 7.105
R299 Q_N Q_N.n3 5.714
R300 Q_N.n2 Q_N 5.042
R301 Q_N.n0 Q_N 2.535
R302 a_1807_47.t0 a_1807_47.t1 60
R303 SCE.n0 SCE.t3 293.601
R304 SCE.n1 SCE.t2 290.645
R305 SCE.n1 SCE.t0 227.906
R306 SCE.n0 SCE.t1 202.561
R307 SCE.n2 SCE.n0 12.836
R308 SCE.n2 SCE.n1 8.407
R309 SCE SCE.n2 3.384
R310 a_109_47.t0 a_109_47.t1 60
R311 a_1514_47.t0 a_1514_47.t1 130.312
R312 a_1712_413.t0 a_1712_413.t1 136.023
R313 a_1879_47.t0 a_1879_47.t1 140
R314 a_319_21.t0 a_319_21.n1 462.451
R315 a_319_21.n0 a_319_21.t2 284.379
R316 a_319_21.n0 a_319_21.t3 191.193
R317 a_319_21.n1 a_319_21.t1 167.058
R318 a_319_21.n1 a_319_21.n0 76
R319 D.n0 D.t0 373.281
R320 D.n0 D.t1 132.281
R321 D.n1 D.n0 76
R322 D.n1 D 23.542
R323 D D.n1 7.542
R324 a_193_369.t0 a_193_369.t1 64.64
R325 a_265_47.t0 a_265_47.t1 77.142
R326 a_1087_47.t0 a_1087_47.t1 60
R327 CLK.n0 CLK.t0 255.075
R328 CLK.n0 CLK.t1 218.64
R329 CLK.n1 CLK.n0 76
R330 CLK.n1 CLK 20.362
R331 CLK CLK.n1 2.909
R332 a_1514_329.t0 a_1514_329.t1 50.422
C0 VPWR Q 0.17fF
C1 VGND Q_N 0.16fF
C2 SCE VGND 0.14fF
C3 SCE CLK 0.10fF
C4 VPB VPWR 0.27fF
C5 SCD SCE 0.21fF
C6 VGND Q 0.12fF
C7 VPWR VGND 0.17fF
C8 VPWR Q_N 0.15fF
C9 SCE D 0.17fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__sdfsbp_2.ext - technology: sky130A

.subckt sky130_fd_sc_hd__sdfsbp_2 SCD CLK Q_N D SET_B SCE Q VPWR VGND VNB VPB
X0 a_1006_47.t2 a_818_47.t2 a_181_47.t4 VPB.t19 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1 a_1781_295.t0 a_1597_329.t5 VPWR.t6 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 VGND.t14 a_328_21.t2 a_265_47.t1 VNB.t22 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3 Q_N.t1 a_1597_329.t6 VGND.t3 VNB.t6 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 a_818_47.t0 a_652_47.t2 VGND.t10 VNB.t12 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 VPWR.t9 a_2501_47.t2 Q.t3 VPB.t9 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 a_1090_47.t1 a_818_47.t3 a_1006_47.t3 VNB.t18 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7 VPWR.t1 SCD.t0 a_27_369.t0 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X8 Q.t2 a_2501_47.t3 VPWR.t10 VPB.t10 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 VPWR.t8 SET_B.t0 a_1132_21.t0 VPB.t8 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10 a_1517_47.t1 a_1006_47.t4 VGND.t13 VNB.t21 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X11 VGND.t9 a_1132_21.t3 a_1090_47.t0 VNB.t11 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12 VGND.t4 a_1597_329.t7 a_2501_47.t0 VNB.t5 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13 a_181_47.t2 SCE.t0 a_109_47.t1 VNB.t15 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14 VPWR.t2 a_1781_295.t2 a_1723_413.t0 VPB.t6 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15 VGND.t11 SCE.t1 a_328_21.t0 VNB.t16 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16 a_1006_47.t0 a_652_47.t3 a_181_47.t1 VNB.t13 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17 VGND.t7 a_2501_47.t4 Q.t1 VNB.t9 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X18 a_818_47.t1 a_652_47.t4 VPWR.t12 VPB.t12 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X19 VGND.t5 SET_B.t1 a_1885_47.t1 VNB.t7 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20 VPWR.t13 SCE.t2 a_328_21.t1 VPB.t15 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X21 a_1597_329.t4 a_818_47.t4 a_1517_47.t0 VNB.t17 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X22 a_181_47.t3 D.t0 a_193_369.t0 VPB.t17 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X23 a_27_369.t1 a_328_21.t3 a_181_47.t5 VPB.t20 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X24 a_1597_329.t1 a_652_47.t5 a_1525_329.t0 VPB.t13 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X25 a_265_47.t0 D.t1 a_181_47.t0 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X26 a_1781_295.t1 a_1597_329.t8 VGND.t1 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X27 a_1813_47.t1 a_652_47.t6 a_1597_329.t2 VNB.t14 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X28 a_1350_47.t1 a_1006_47.t5 a_1132_21.t1 VNB.t20 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X29 Q.t0 a_2501_47.t5 VGND.t8 VNB.t10 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X30 a_193_369.t1 SCE.t3 VPWR.t14 VPB.t16 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X31 a_1525_329.t1 a_1006_47.t6 VPWR.t15 VPB.t22 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X32 a_1723_413.t1 a_818_47.t5 a_1597_329.t3 VPB.t18 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X33 a_1885_47.t0 a_1781_295.t3 a_1813_47.t0 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X34 VPWR.t4 a_1597_329.t9 Q_N.t3 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X35 VGND.t12 CLK.t0 a_652_47.t1 VNB.t19 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X36 VPWR.t0 CLK.t1 a_652_47.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X37 VPWR.t11 a_1132_21.t4 a_1102_413.t0 VPB.t11 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X38 a_1132_21.t2 a_1006_47.t7 VPWR.t16 VPB.t21 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X39 VGND.t6 SET_B.t2 a_1350_47.t0 VNB.t8 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X40 VGND.t2 a_1597_329.t10 Q_N.t0 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X41 a_1102_413.t1 a_652_47.t7 a_1006_47.t1 VPB.t14 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X42 Q_N.t2 a_1597_329.t11 VPWR.t3 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X43 VPWR.t5 a_1597_329.t12 a_2501_47.t1 VPB.t5 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X44 a_1597_329.t0 SET_B.t3 VPWR.t7 VPB.t7 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X45 a_109_47.t0 SCD.t1 VGND.t0 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
R0 a_818_47.n0 a_818_47.t4 385.062
R1 a_818_47.n2 a_818_47.t3 383.313
R2 a_818_47.t1 a_818_47.n3 382.013
R3 a_818_47.n2 a_818_47.t2 319.726
R4 a_818_47.n1 a_818_47.t0 182.04
R5 a_818_47.n0 a_818_47.t5 148.348
R6 a_818_47.n1 a_818_47.n0 116.666
R7 a_818_47.n3 a_818_47.n2 46.649
R8 a_818_47.n3 a_818_47.n1 1.197
R9 a_181_47.n0 a_181_47.t4 399.073
R10 a_181_47.n3 a_181_47.n2 318.426
R11 a_181_47.n0 a_181_47.t1 193.322
R12 a_181_47.n2 a_181_47.n1 175.878
R13 a_181_47.t3 a_181_47.n3 60.023
R14 a_181_47.n3 a_181_47.t5 41.554
R15 a_181_47.n1 a_181_47.t0 38.571
R16 a_181_47.n1 a_181_47.t2 38.571
R17 a_181_47.n2 a_181_47.n0 12.398
R18 a_1006_47.n4 a_1006_47.n0 367.417
R19 a_1006_47.n1 a_1006_47.t7 312.131
R20 a_1006_47.n2 a_1006_47.t6 263.861
R21 a_1006_47.n1 a_1006_47.t5 243.044
R22 a_1006_47.n2 a_1006_47.t4 167.461
R23 a_1006_47.n5 a_1006_47.n4 149.577
R24 a_1006_47.n3 a_1006_47.n2 125.108
R25 a_1006_47.n0 a_1006_47.t2 89.119
R26 a_1006_47.n3 a_1006_47.n1 76
R27 a_1006_47.n0 a_1006_47.t1 63.321
R28 a_1006_47.n4 a_1006_47.n3 50.07
R29 a_1006_47.n5 a_1006_47.t3 38.571
R30 a_1006_47.t0 a_1006_47.n5 38.571
R31 VPB.t3 VPB.t5 594.859
R32 VPB.t2 VPB.t4 556.386
R33 VPB.t7 VPB.t2 556.386
R34 VPB.t12 VPB.t19 556.386
R35 VPB.t15 VPB.t0 556.386
R36 VPB.t20 VPB.t15 550.467
R37 VPB.t13 VPB.t18 372.897
R38 VPB.t11 VPB.t21 352.18
R39 VPB.t8 VPB.t22 343.302
R40 VPB.t6 VPB.t7 328.504
R41 VPB.t21 VPB.t8 290.031
R42 VPB.t17 VPB.t20 284.112
R43 VPB.t5 VPB.t10 281.152
R44 VPB.t19 VPB.t14 281.152
R45 VPB.t14 VPB.t11 266.355
R46 VPB.t18 VPB.t6 260.436
R47 VPB.t10 VPB.t9 248.598
R48 VPB.t4 VPB.t3 248.598
R49 VPB.t0 VPB.t12 248.598
R50 VPB.t1 VPB.t16 248.598
R51 VPB.t22 VPB.t13 213.084
R52 VPB.t16 VPB.t17 213.084
R53 VPB VPB.t1 192.367
R54 a_1597_329.n8 a_1597_329.n7 378.126
R55 a_1597_329.n7 a_1597_329.t0 370.28
R56 a_1597_329.n4 a_1597_329.n3 301.205
R57 a_1597_329.n0 a_1597_329.t12 249.032
R58 a_1597_329.n1 a_1597_329.t9 212.079
R59 a_1597_329.n2 a_1597_329.t11 212.079
R60 a_1597_329.n0 a_1597_329.t7 176.733
R61 a_1597_329.n6 a_1597_329.t5 167.037
R62 a_1597_329.n5 a_1597_329.n2 147.521
R63 a_1597_329.n1 a_1597_329.n0 146.79
R64 a_1597_329.n1 a_1597_329.t10 139.779
R65 a_1597_329.n2 a_1597_329.t6 139.779
R66 a_1597_329.n4 a_1597_329.t8 132.281
R67 a_1597_329.t1 a_1597_329.n8 104.362
R68 a_1597_329.n7 a_1597_329.n6 100.597
R69 a_1597_329.n8 a_1597_329.t3 91.464
R70 a_1597_329.n3 a_1597_329.t2 81.428
R71 a_1597_329.n2 a_1597_329.n1 61.345
R72 a_1597_329.n6 a_1597_329.n5 60.665
R73 a_1597_329.n3 a_1597_329.t4 34.865
R74 a_1597_329.n5 a_1597_329.n4 13.063
R75 VPWR.n50 VPWR.t13 425.096
R76 VPWR.n13 VPWR.t6 370.56
R77 VPWR.n18 VPWR.n17 306.463
R78 VPWR.n35 VPWR.n34 306.463
R79 VPWR.n46 VPWR.n45 306.463
R80 VPWR.n62 VPWR.n61 306.463
R81 VPWR.n29 VPWR.n28 292.5
R82 VPWR.n1 VPWR.n0 165.298
R83 VPWR.n2 VPWR.t9 165.091
R84 VPWR.n5 VPWR.t4 161.63
R85 VPWR.n9 VPWR.t3 158.058
R86 VPWR.n17 VPWR.t2 126.642
R87 VPWR.n34 VPWR.t16 112.571
R88 VPWR.n34 VPWR.t11 96.154
R89 VPWR.n28 VPWR.t15 87.945
R90 VPWR.n28 VPWR.t8 84.428
R91 VPWR.n17 VPWR.t7 63.321
R92 VPWR.n0 VPWR.t5 56.945
R93 VPWR.n45 VPWR.t12 41.554
R94 VPWR.n45 VPWR.t0 41.554
R95 VPWR.n61 VPWR.t14 41.554
R96 VPWR.n61 VPWR.t1 41.554
R97 VPWR.n0 VPWR.t10 33.109
R98 VPWR.n4 VPWR.n3 4.65
R99 VPWR.n6 VPWR.n5 4.65
R100 VPWR.n8 VPWR.n7 4.65
R101 VPWR.n10 VPWR.n9 4.65
R102 VPWR.n12 VPWR.n11 4.65
R103 VPWR.n14 VPWR.n13 4.65
R104 VPWR.n16 VPWR.n15 4.65
R105 VPWR.n19 VPWR.n18 4.65
R106 VPWR.n21 VPWR.n20 4.65
R107 VPWR.n23 VPWR.n22 4.65
R108 VPWR.n25 VPWR.n24 4.65
R109 VPWR.n27 VPWR.n26 4.65
R110 VPWR.n31 VPWR.n30 4.65
R111 VPWR.n33 VPWR.n32 4.65
R112 VPWR.n36 VPWR.n35 4.65
R113 VPWR.n38 VPWR.n37 4.65
R114 VPWR.n40 VPWR.n39 4.65
R115 VPWR.n42 VPWR.n41 4.65
R116 VPWR.n44 VPWR.n43 4.65
R117 VPWR.n47 VPWR.n46 4.65
R118 VPWR.n49 VPWR.n48 4.65
R119 VPWR.n52 VPWR.n51 4.65
R120 VPWR.n54 VPWR.n53 4.65
R121 VPWR.n56 VPWR.n55 4.65
R122 VPWR.n58 VPWR.n57 4.65
R123 VPWR.n60 VPWR.n59 4.65
R124 VPWR.n63 VPWR.n62 3.932
R125 VPWR.n2 VPWR.n1 3.904
R126 VPWR.n51 VPWR.n50 2.309
R127 VPWR.n30 VPWR.n29 1.788
R128 VPWR.n4 VPWR.n2 0.224
R129 VPWR.n63 VPWR.n60 0.137
R130 VPWR VPWR.n63 0.123
R131 VPWR.n6 VPWR.n4 0.119
R132 VPWR.n8 VPWR.n6 0.119
R133 VPWR.n10 VPWR.n8 0.119
R134 VPWR.n12 VPWR.n10 0.119
R135 VPWR.n14 VPWR.n12 0.119
R136 VPWR.n16 VPWR.n14 0.119
R137 VPWR.n19 VPWR.n16 0.119
R138 VPWR.n21 VPWR.n19 0.119
R139 VPWR.n23 VPWR.n21 0.119
R140 VPWR.n25 VPWR.n23 0.119
R141 VPWR.n27 VPWR.n25 0.119
R142 VPWR.n31 VPWR.n27 0.119
R143 VPWR.n33 VPWR.n31 0.119
R144 VPWR.n36 VPWR.n33 0.119
R145 VPWR.n38 VPWR.n36 0.119
R146 VPWR.n40 VPWR.n38 0.119
R147 VPWR.n42 VPWR.n40 0.119
R148 VPWR.n44 VPWR.n42 0.119
R149 VPWR.n47 VPWR.n44 0.119
R150 VPWR.n49 VPWR.n47 0.119
R151 VPWR.n52 VPWR.n49 0.119
R152 VPWR.n54 VPWR.n52 0.119
R153 VPWR.n56 VPWR.n54 0.119
R154 VPWR.n58 VPWR.n56 0.119
R155 VPWR.n60 VPWR.n58 0.119
R156 a_1781_295.n0 a_1781_295.t2 448.369
R157 a_1781_295.t0 a_1781_295.n1 404.408
R158 a_1781_295.n1 a_1781_295.t1 193.167
R159 a_1781_295.n1 a_1781_295.n0 180.642
R160 a_1781_295.n0 a_1781_295.t3 159.17
R161 a_328_21.n2 a_328_21.n1 336.204
R162 a_328_21.n0 a_328_21.t3 269.919
R163 a_328_21.n0 a_328_21.t2 178.923
R164 a_328_21.n1 a_328_21.t0 167.863
R165 a_328_21.n2 a_328_21.t1 129.49
R166 a_328_21.n1 a_328_21.n0 124.93
R167 a_328_21.n3 a_328_21.n2 3.788
R168 a_265_47.t0 a_265_47.t1 90
R169 VGND.n57 VGND.t14 150.527
R170 VGND.n65 VGND.t0 131.071
R171 VGND.n52 VGND.t11 131.071
R172 VGND.n38 VGND.t9 131.071
R173 VGND.n9 VGND.t3 113.911
R174 VGND.n15 VGND.n14 110.932
R175 VGND.n48 VGND.n47 107.86
R176 VGND.n2 VGND.t7 106.649
R177 VGND.n1 VGND.n0 105.48
R178 VGND.n5 VGND.t2 103.416
R179 VGND.n31 VGND.n30 92.5
R180 VGND.n14 VGND.t5 55.714
R181 VGND.n0 VGND.t4 45.714
R182 VGND.n30 VGND.t13 42.008
R183 VGND.n14 VGND.t1 40
R184 VGND.n30 VGND.t6 38.571
R185 VGND.n47 VGND.t10 38.571
R186 VGND.n47 VGND.t12 38.571
R187 VGND.n0 VGND.t8 34.505
R188 VGND.n66 VGND.n65 5.214
R189 VGND.n10 VGND.n9 4.894
R190 VGND.n16 VGND.n15 4.894
R191 VGND.n4 VGND.n3 4.65
R192 VGND.n6 VGND.n5 4.65
R193 VGND.n8 VGND.n7 4.65
R194 VGND.n11 VGND.n10 4.65
R195 VGND.n13 VGND.n12 4.65
R196 VGND.n17 VGND.n16 4.65
R197 VGND.n19 VGND.n18 4.65
R198 VGND.n21 VGND.n20 4.65
R199 VGND.n23 VGND.n22 4.65
R200 VGND.n25 VGND.n24 4.65
R201 VGND.n27 VGND.n26 4.65
R202 VGND.n29 VGND.n28 4.65
R203 VGND.n33 VGND.n32 4.65
R204 VGND.n35 VGND.n34 4.65
R205 VGND.n37 VGND.n36 4.65
R206 VGND.n40 VGND.n39 4.65
R207 VGND.n42 VGND.n41 4.65
R208 VGND.n44 VGND.n43 4.65
R209 VGND.n46 VGND.n45 4.65
R210 VGND.n49 VGND.n48 4.65
R211 VGND.n51 VGND.n50 4.65
R212 VGND.n54 VGND.n53 4.65
R213 VGND.n56 VGND.n55 4.65
R214 VGND.n58 VGND.n57 4.65
R215 VGND.n60 VGND.n59 4.65
R216 VGND.n62 VGND.n61 4.65
R217 VGND.n64 VGND.n63 4.65
R218 VGND.n39 VGND.n38 4.538
R219 VGND.n2 VGND.n1 3.904
R220 VGND.n53 VGND.n52 2.5
R221 VGND.n32 VGND.n31 1.653
R222 VGND.n4 VGND.n2 0.224
R223 VGND.n6 VGND.n4 0.119
R224 VGND.n8 VGND.n6 0.119
R225 VGND.n11 VGND.n8 0.119
R226 VGND.n13 VGND.n11 0.119
R227 VGND.n17 VGND.n13 0.119
R228 VGND.n19 VGND.n17 0.119
R229 VGND.n21 VGND.n19 0.119
R230 VGND.n23 VGND.n21 0.119
R231 VGND.n25 VGND.n23 0.119
R232 VGND.n27 VGND.n25 0.119
R233 VGND.n29 VGND.n27 0.119
R234 VGND.n33 VGND.n29 0.119
R235 VGND.n35 VGND.n33 0.119
R236 VGND.n37 VGND.n35 0.119
R237 VGND.n40 VGND.n37 0.119
R238 VGND.n42 VGND.n40 0.119
R239 VGND.n44 VGND.n42 0.119
R240 VGND.n46 VGND.n44 0.119
R241 VGND.n49 VGND.n46 0.119
R242 VGND.n51 VGND.n49 0.119
R243 VGND.n54 VGND.n51 0.119
R244 VGND.n56 VGND.n54 0.119
R245 VGND.n58 VGND.n56 0.119
R246 VGND.n60 VGND.n58 0.119
R247 VGND.n62 VGND.n60 0.119
R248 VGND.n64 VGND.n62 0.119
R249 VGND.n66 VGND.n64 0.119
R250 VGND VGND.n66 0.022
R251 VNB VNB.t2 6470.59
R252 VNB.t4 VNB.t6 6227.76
R253 VNB.t11 VNB.t20 6082.35
R254 VNB.t12 VNB.t13 6082.35
R255 VNB.t16 VNB.t19 6082.35
R256 VNB.t22 VNB.t16 6082.35
R257 VNB.t3 VNB.t5 4859.34
R258 VNB.t21 VNB.t17 4302.22
R259 VNB.t1 VNB.t7 3235.29
R260 VNB.t17 VNB.t14 3162.68
R261 VNB.t7 VNB.t4 3138.24
R262 VNB.t0 VNB.t22 3008.82
R263 VNB.t13 VNB.t18 2717.65
R264 VNB.t19 VNB.t12 2717.65
R265 VNB.t15 VNB.t0 2717.65
R266 VNB.t14 VNB.t1 2329.41
R267 VNB.t20 VNB.t8 2329.41
R268 VNB.t18 VNB.t11 2329.41
R269 VNB.t2 VNB.t15 2329.41
R270 VNB.t5 VNB.t10 2296.7
R271 VNB.t8 VNB.t21 2280.14
R272 VNB.t10 VNB.t9 2030.77
R273 VNB.t6 VNB.t3 2030.77
R274 Q_N.n2 Q_N.n1 292.5
R275 Q_N.n1 Q_N.n0 146.887
R276 Q_N Q_N.n4 93.958
R277 Q_N.n1 Q_N.t3 26.595
R278 Q_N.n1 Q_N.t2 26.595
R279 Q_N.n4 Q_N.t0 24.923
R280 Q_N.n4 Q_N.t1 24.923
R281 Q_N Q_N.n3 9.559
R282 Q_N.n0 Q_N 8.873
R283 Q_N Q_N.n2 6.805
R284 Q_N.n2 Q_N 4.212
R285 Q_N.n0 Q_N 2.116
R286 Q_N.n3 Q_N 1.458
R287 a_652_47.n2 a_652_47.t3 393.633
R288 a_652_47.t0 a_652_47.n5 371.142
R289 a_652_47.n0 a_652_47.t6 353.209
R290 a_652_47.n0 a_652_47.t5 343.241
R291 a_652_47.n3 a_652_47.t4 249.394
R292 a_652_47.n4 a_652_47.t1 196.463
R293 a_652_47.n1 a_652_47.t7 147.445
R294 a_652_47.n3 a_652_47.n2 105.025
R295 a_652_47.n2 a_652_47.t2 91.58
R296 a_652_47.n4 a_652_47.n3 76
R297 a_652_47.n1 a_652_47.n0 64.281
R298 a_652_47.n5 a_652_47.n4 30.276
R299 a_652_47.n5 a_652_47.n1 5.824
R300 a_2501_47.t1 a_2501_47.n2 258.462
R301 a_2501_47.n0 a_2501_47.t2 212.079
R302 a_2501_47.n1 a_2501_47.t3 212.079
R303 a_2501_47.n2 a_2501_47.t0 169.471
R304 a_2501_47.n0 a_2501_47.t4 139.779
R305 a_2501_47.n1 a_2501_47.t5 139.779
R306 a_2501_47.n2 a_2501_47.n1 108.857
R307 a_2501_47.n1 a_2501_47.n0 61.345
R308 Q.n1 Q.n0 146.061
R309 Q.n5 Q.n4 92.5
R310 Q.n0 Q.t3 26.595
R311 Q.n0 Q.t2 26.595
R312 Q.n4 Q.t1 24.923
R313 Q.n4 Q.t0 24.923
R314 Q.n3 Q 15.928
R315 Q Q.n5 12.606
R316 Q.n2 Q 11.248
R317 Q Q.n1 9.62
R318 Q.n1 Q 3.486
R319 Q.n3 Q 3.413
R320 Q Q.n2 2.844
R321 Q Q.n3 2.327
R322 Q.n2 Q 1.939
R323 Q.n5 Q 0.581
R324 a_1090_47.t0 a_1090_47.t1 60
R325 SCD.n0 SCD.t0 299.43
R326 SCD.n0 SCD.t1 206.244
R327 SCD.n1 SCD.n0 76
R328 SCD.n1 SCD 19.827
R329 SCD SCD.n1 14.305
R330 a_27_369.t0 a_27_369.t1 784.249
R331 SET_B.n1 SET_B.t1 358.397
R332 SET_B.n0 SET_B.t2 357.656
R333 SET_B.n1 SET_B.t3 170.194
R334 SET_B.n0 SET_B.t0 166.576
R335 SET_B.n2 SET_B.n1 134.344
R336 SET_B.n2 SET_B.n0 83
R337 SET_B SET_B.n2 3.4
R338 a_1132_21.n2 a_1132_21.n1 439.993
R339 a_1132_21.n0 a_1132_21.t1 251.077
R340 a_1132_21.n1 a_1132_21.n0 201.407
R341 a_1132_21.n1 a_1132_21.t4 139.55
R342 a_1132_21.n0 a_1132_21.t3 129.336
R343 a_1132_21.t0 a_1132_21.n2 84.428
R344 a_1132_21.n2 a_1132_21.t2 75.047
R345 a_1517_47.t0 a_1517_47.t1 136.875
R346 SCE.n0 SCE.t2 294.778
R347 SCE.n1 SCE.t3 292.153
R348 SCE.n1 SCE.t0 227.541
R349 SCE.n0 SCE.t1 203.815
R350 SCE.n2 SCE.n0 13.068
R351 SCE.n2 SCE.n1 8.415
R352 SCE SCE.n2 3.384
R353 a_109_47.t0 a_109_47.t1 60
R354 a_1723_413.t0 a_1723_413.t1 136.023
R355 a_1885_47.t0 a_1885_47.t1 100
R356 D.n0 D.t0 373.281
R357 D.n0 D.t1 132.281
R358 D.n1 D.n0 76
R359 D.n1 D 23.129
R360 D D.n1 7.41
R361 a_193_369.t0 a_193_369.t1 64.64
R362 a_1525_329.t0 a_1525_329.t1 49.25
R363 a_1813_47.t0 a_1813_47.t1 60
R364 a_1350_47.t0 a_1350_47.t1 60
R365 CLK.n0 CLK.t1 248.454
R366 CLK.n0 CLK.t0 216.867
R367 CLK.n1 CLK.n0 76
R368 CLK.n1 CLK 18.139
R369 CLK CLK.n1 2.909
R370 a_1102_413.t0 a_1102_413.t1 140.714
C0 VPWR Q_N 0.32fF
C1 SCE D 0.17fF
C2 VGND Q_N 0.28fF
C3 VPWR Q 0.32fF
C4 SCE VGND 0.16fF
C5 SCE CLK 0.11fF
C6 VPB VPWR 0.30fF
C7 SCD SCE 0.21fF
C8 VGND Q 0.22fF
C9 VPWR VGND 0.22fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__sdfstp_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__sdfstp_1 SCD CLK D SET_B SCE Q VPWR VGND VNB VPB
X0 VPWR.t0 a_1597_329.t5 a_2227_47.t0 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1 Q.t0 a_2227_47.t2 VGND.t3 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 a_1597_329.t2 SET_B.t0 VPWR.t6 VPB.t8 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3 VPWR.t3 SCD.t0 a_27_369.t1 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X4 a_1081_413.t0 a_643_369.t2 a_997_413.t1 VPB.t17 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 a_809_369.t0 a_643_369.t3 VGND.t11 VNB.t17 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 VGND.t0 a_1597_329.t6 a_2227_47.t1 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7 a_997_413.t3 a_809_369.t2 a_181_47.t2 VPB.t10 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 VPWR.t7 SET_B.t1 a_1129_21.t2 VPB.t9 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9 a_1347_47.t0 a_997_413.t4 a_1129_21.t0 VNB.t7 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10 VPWR.t8 a_1129_21.t3 a_1081_413.t1 VPB.t11 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11 a_181_47.t0 SCE.t0 a_109_47.t0 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12 a_1514_47.t0 a_997_413.t5 VGND.t4 VNB.t8 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X13 VPWR.t9 a_1781_295.t2 a_1723_413.t1 VPB.t12 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14 VGND.t5 SET_B.t2 a_1347_47.t1 VNB.t9 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15 a_27_369.t0 a_319_21.t2 a_181_47.t4 VPB.t13 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X16 VGND.t10 SCE.t1 a_319_21.t0 VNB.t15 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17 a_1597_329.t0 a_809_369.t3 a_1514_47.t1 VNB.t5 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X18 a_1815_47.t0 a_643_369.t4 a_1597_329.t3 VNB.t18 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19 a_181_47.t1 D.t0 a_193_369.t1 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X20 VGND.t6 SET_B.t3 a_1887_47.t0 VNB.t10 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21 a_1597_329.t4 a_643_369.t5 a_1525_329.t1 VPB.t18 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X22 a_265_47.t1 D.t1 a_181_47.t5 VNB.t16 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23 a_997_413.t0 a_643_369.t6 a_181_47.t3 VNB.t19 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24 a_1781_295.t0 a_1597_329.t7 VGND.t1 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X25 a_1887_47.t1 a_1781_295.t3 a_1815_47.t1 VNB.t13 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X26 a_1087_47.t0 a_809_369.t4 a_997_413.t2 VNB.t6 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X27 a_193_369.t0 SCE.t2 VPWR.t10 VPB.t14 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X28 a_809_369.t1 a_643_369.t7 VPWR.t13 VPB.t19 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X29 a_1525_329.t0 a_997_413.t6 VPWR.t4 VPB.t6 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X30 a_1723_413.t0 a_809_369.t5 a_1597_329.t1 VPB.t5 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X31 VPWR.t11 SCE.t3 a_319_21.t1 VPB.t15 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X32 Q.t1 a_2227_47.t3 VPWR.t2 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X33 VPWR.t12 CLK.t0 a_643_369.t1 VPB.t16 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X34 a_1129_21.t1 a_997_413.t7 VPWR.t5 VPB.t7 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X35 VGND.t9 a_319_21.t3 a_265_47.t0 VNB.t14 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X36 VGND.t8 a_1129_21.t4 a_1087_47.t1 VNB.t12 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X37 VGND.t2 CLK.t1 a_643_369.t0 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X38 a_1781_295.t1 a_1597_329.t8 VPWR.t1 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X39 a_109_47.t1 SCD.t1 VGND.t7 VNB.t11 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
R0 a_1597_329.n6 a_1597_329.n5 381.354
R1 a_1597_329.n2 a_1597_329.t6 356.68
R2 a_1597_329.n5 a_1597_329.t2 355.821
R3 a_1597_329.n3 a_1597_329.n2 291.341
R4 a_1597_329.n1 a_1597_329.n0 269.852
R5 a_1597_329.n3 a_1597_329.t8 144.6
R6 a_1597_329.n2 a_1597_329.t5 133.352
R7 a_1597_329.n1 a_1597_329.t7 132.281
R8 a_1597_329.n4 a_1597_329.n1 111.574
R9 a_1597_329.n5 a_1597_329.n4 110.713
R10 a_1597_329.t4 a_1597_329.n6 104.362
R11 a_1597_329.n6 a_1597_329.t1 91.464
R12 a_1597_329.n0 a_1597_329.t3 84.285
R13 a_1597_329.n0 a_1597_329.t0 34.865
R14 a_1597_329.n4 a_1597_329.n3 32.133
R15 a_2227_47.t0 a_2227_47.n1 245.338
R16 a_2227_47.n0 a_2227_47.t3 241.534
R17 a_2227_47.n0 a_2227_47.t2 169.234
R18 a_2227_47.n1 a_2227_47.t1 158.394
R19 a_2227_47.n1 a_2227_47.n0 102.181
R20 VPWR.n39 VPWR.t11 441.584
R21 VPWR.n0 VPWR.t1 370.56
R22 VPWR.n51 VPWR.n50 309.566
R23 VPWR.n6 VPWR.n5 306.463
R24 VPWR.n35 VPWR.n34 306.463
R25 VPWR.n17 VPWR.n16 292.5
R26 VPWR.n23 VPWR.n22 292.5
R27 VPWR.n2 VPWR.n1 170.964
R28 VPWR.n22 VPWR.t5 138.369
R29 VPWR.n5 VPWR.t9 126.642
R30 VPWR.n22 VPWR.t8 91.464
R31 VPWR.n5 VPWR.t6 89.119
R32 VPWR.n16 VPWR.t4 87.945
R33 VPWR.n16 VPWR.t7 84.428
R34 VPWR.n1 VPWR.t0 60.023
R35 VPWR.n34 VPWR.t13 41.554
R36 VPWR.n34 VPWR.t12 41.554
R37 VPWR.n50 VPWR.t10 41.554
R38 VPWR.n50 VPWR.t3 41.554
R39 VPWR.n1 VPWR.t2 31.137
R40 VPWR.n4 VPWR.n3 4.65
R41 VPWR.n7 VPWR.n6 4.65
R42 VPWR.n9 VPWR.n8 4.65
R43 VPWR.n11 VPWR.n10 4.65
R44 VPWR.n13 VPWR.n12 4.65
R45 VPWR.n15 VPWR.n14 4.65
R46 VPWR.n19 VPWR.n18 4.65
R47 VPWR.n21 VPWR.n20 4.65
R48 VPWR.n25 VPWR.n24 4.65
R49 VPWR.n27 VPWR.n26 4.65
R50 VPWR.n29 VPWR.n28 4.65
R51 VPWR.n31 VPWR.n30 4.65
R52 VPWR.n33 VPWR.n32 4.65
R53 VPWR.n36 VPWR.n35 4.65
R54 VPWR.n38 VPWR.n37 4.65
R55 VPWR.n41 VPWR.n40 4.65
R56 VPWR.n43 VPWR.n42 4.65
R57 VPWR.n45 VPWR.n44 4.65
R58 VPWR.n47 VPWR.n46 4.65
R59 VPWR.n49 VPWR.n48 4.65
R60 VPWR.n2 VPWR.n0 3.974
R61 VPWR.n52 VPWR.n51 3.932
R62 VPWR.n24 VPWR.n23 2.415
R63 VPWR.n18 VPWR.n17 1.788
R64 VPWR.n40 VPWR.n39 0.376
R65 VPWR.n4 VPWR.n2 0.149
R66 VPWR.n52 VPWR.n49 0.137
R67 VPWR VPWR.n52 0.123
R68 VPWR.n7 VPWR.n4 0.119
R69 VPWR.n9 VPWR.n7 0.119
R70 VPWR.n11 VPWR.n9 0.119
R71 VPWR.n13 VPWR.n11 0.119
R72 VPWR.n15 VPWR.n13 0.119
R73 VPWR.n19 VPWR.n15 0.119
R74 VPWR.n21 VPWR.n19 0.119
R75 VPWR.n25 VPWR.n21 0.119
R76 VPWR.n27 VPWR.n25 0.119
R77 VPWR.n29 VPWR.n27 0.119
R78 VPWR.n31 VPWR.n29 0.119
R79 VPWR.n33 VPWR.n31 0.119
R80 VPWR.n36 VPWR.n33 0.119
R81 VPWR.n38 VPWR.n36 0.119
R82 VPWR.n41 VPWR.n38 0.119
R83 VPWR.n43 VPWR.n41 0.119
R84 VPWR.n45 VPWR.n43 0.119
R85 VPWR.n47 VPWR.n45 0.119
R86 VPWR.n49 VPWR.n47 0.119
R87 VPB.t0 VPB.t1 556.386
R88 VPB.t8 VPB.t0 556.386
R89 VPB.t19 VPB.t10 556.386
R90 VPB.t15 VPB.t16 556.386
R91 VPB.t13 VPB.t15 556.386
R92 VPB.t11 VPB.t7 378.816
R93 VPB.t18 VPB.t5 372.897
R94 VPB.t12 VPB.t8 361.059
R95 VPB.t9 VPB.t6 343.302
R96 VPB.t17 VPB.t11 301.869
R97 VPB.t7 VPB.t9 290.031
R98 VPB.t1 VPB.t2 284.112
R99 VPB.t5 VPB.t12 260.436
R100 VPB.t10 VPB.t17 248.598
R101 VPB.t16 VPB.t19 248.598
R102 VPB.t3 VPB.t13 248.598
R103 VPB.t4 VPB.t14 248.598
R104 VPB.t6 VPB.t18 213.084
R105 VPB.t14 VPB.t3 213.084
R106 VPB VPB.t4 192.367
R107 VGND.n43 VGND.t9 157.996
R108 VGND.n51 VGND.t7 131.071
R109 VGND.n38 VGND.t10 131.071
R110 VGND.n24 VGND.t8 131.071
R111 VGND.n3 VGND.n0 111.107
R112 VGND.n2 VGND.n1 110.932
R113 VGND.n34 VGND.n33 106.463
R114 VGND.n17 VGND.n16 92.5
R115 VGND.n1 VGND.t6 81.428
R116 VGND.n0 VGND.t0 55.714
R117 VGND.n16 VGND.t5 41.428
R118 VGND.n16 VGND.t4 39.151
R119 VGND.n1 VGND.t1 38.571
R120 VGND.n33 VGND.t11 38.571
R121 VGND.n33 VGND.t2 38.571
R122 VGND.n0 VGND.t3 25.934
R123 VGND.n52 VGND.n51 5.214
R124 VGND.n5 VGND.n4 4.65
R125 VGND.n7 VGND.n6 4.65
R126 VGND.n9 VGND.n8 4.65
R127 VGND.n11 VGND.n10 4.65
R128 VGND.n13 VGND.n12 4.65
R129 VGND.n15 VGND.n14 4.65
R130 VGND.n19 VGND.n18 4.65
R131 VGND.n21 VGND.n20 4.65
R132 VGND.n23 VGND.n22 4.65
R133 VGND.n26 VGND.n25 4.65
R134 VGND.n28 VGND.n27 4.65
R135 VGND.n30 VGND.n29 4.65
R136 VGND.n32 VGND.n31 4.65
R137 VGND.n35 VGND.n34 4.65
R138 VGND.n37 VGND.n36 4.65
R139 VGND.n40 VGND.n39 4.65
R140 VGND.n42 VGND.n41 4.65
R141 VGND.n44 VGND.n43 4.65
R142 VGND.n46 VGND.n45 4.65
R143 VGND.n48 VGND.n47 4.65
R144 VGND.n50 VGND.n49 4.65
R145 VGND.n25 VGND.n24 4.189
R146 VGND.n3 VGND.n2 4.118
R147 VGND.n39 VGND.n38 2.8
R148 VGND.n18 VGND.n17 1.582
R149 VGND.n5 VGND.n3 0.142
R150 VGND.n7 VGND.n5 0.119
R151 VGND.n9 VGND.n7 0.119
R152 VGND.n11 VGND.n9 0.119
R153 VGND.n13 VGND.n11 0.119
R154 VGND.n15 VGND.n13 0.119
R155 VGND.n19 VGND.n15 0.119
R156 VGND.n21 VGND.n19 0.119
R157 VGND.n23 VGND.n21 0.119
R158 VGND.n26 VGND.n23 0.119
R159 VGND.n28 VGND.n26 0.119
R160 VGND.n30 VGND.n28 0.119
R161 VGND.n32 VGND.n30 0.119
R162 VGND.n35 VGND.n32 0.119
R163 VGND.n37 VGND.n35 0.119
R164 VGND.n40 VGND.n37 0.119
R165 VGND.n42 VGND.n40 0.119
R166 VGND.n44 VGND.n42 0.119
R167 VGND.n46 VGND.n44 0.119
R168 VGND.n48 VGND.n46 0.119
R169 VGND.n50 VGND.n48 0.119
R170 VGND.n52 VGND.n50 0.119
R171 VGND VGND.n52 0.022
R172 Q.n0 Q.t1 172.661
R173 Q.n3 Q.t0 117.423
R174 Q.n2 Q 18.863
R175 Q Q.n3 12.235
R176 Q.n1 Q 10.917
R177 Q Q.n0 9.339
R178 Q.n2 Q 4.042
R179 Q.n0 Q 3.384
R180 Q Q.n1 3.368
R181 Q Q.n2 2.258
R182 Q.n1 Q 1.882
R183 Q.n3 Q 0.564
R184 VNB.t0 VNB.t1 6858.82
R185 VNB VNB.t11 6470.59
R186 VNB.t14 VNB.t15 6276.47
R187 VNB.t12 VNB.t7 6082.35
R188 VNB.t17 VNB.t19 6082.35
R189 VNB.t15 VNB.t2 6082.35
R190 VNB.t8 VNB.t5 4375.56
R191 VNB.t10 VNB.t0 3688.24
R192 VNB.t5 VNB.t18 3227.39
R193 VNB.t13 VNB.t10 3105.88
R194 VNB.t19 VNB.t6 2717.65
R195 VNB.t2 VNB.t17 2717.65
R196 VNB.t16 VNB.t14 2717.65
R197 VNB.t4 VNB.t16 2717.65
R198 VNB.t18 VNB.t13 2329.41
R199 VNB.t7 VNB.t9 2329.41
R200 VNB.t6 VNB.t12 2329.41
R201 VNB.t11 VNB.t4 2329.41
R202 VNB.t9 VNB.t8 2280.14
R203 VNB.t1 VNB.t3 2269.18
R204 SET_B.n0 SET_B.t2 360.179
R205 SET_B.n1 SET_B.t3 357.215
R206 SET_B.n0 SET_B.t1 166.576
R207 SET_B.n1 SET_B.t0 161.029
R208 SET_B.n2 SET_B.n1 137.809
R209 SET_B.n2 SET_B.n0 83
R210 SET_B SET_B.n2 3.4
R211 SCD.n0 SCD.t0 299.43
R212 SCD.n0 SCD.t1 206.244
R213 SCD.n1 SCD.n0 76
R214 SCD.n1 SCD 19.827
R215 SCD SCD.n1 14.305
R216 a_27_369.t0 a_27_369.t1 883.735
R217 a_643_369.n2 a_643_369.t6 393.633
R218 a_643_369.t1 a_643_369.n5 377.811
R219 a_643_369.n0 a_643_369.t5 343.241
R220 a_643_369.n0 a_643_369.t4 337.584
R221 a_643_369.n3 a_643_369.t7 267.297
R222 a_643_369.n4 a_643_369.t0 199.461
R223 a_643_369.n1 a_643_369.t2 147.521
R224 a_643_369.n3 a_643_369.n2 100.205
R225 a_643_369.n2 a_643_369.t3 91.58
R226 a_643_369.n4 a_643_369.n3 76
R227 a_643_369.n1 a_643_369.n0 49.157
R228 a_643_369.n5 a_643_369.n4 30.276
R229 a_643_369.n5 a_643_369.n1 5.776
R230 a_997_413.n4 a_997_413.n0 369.55
R231 a_997_413.n1 a_997_413.t7 312.131
R232 a_997_413.n2 a_997_413.t6 262.639
R233 a_997_413.n1 a_997_413.t4 238.224
R234 a_997_413.n2 a_997_413.t5 166.239
R235 a_997_413.n5 a_997_413.n4 141.906
R236 a_997_413.n3 a_997_413.n2 124.559
R237 a_997_413.n3 a_997_413.n1 76
R238 a_997_413.n0 a_997_413.t1 63.321
R239 a_997_413.n0 a_997_413.t3 63.321
R240 a_997_413.n4 a_997_413.n3 53.834
R241 a_997_413.n5 a_997_413.t2 38.571
R242 a_997_413.t0 a_997_413.n5 38.571
R243 a_1081_413.t0 a_1081_413.t1 168.857
R244 a_809_369.n2 a_809_369.t4 433.507
R245 a_809_369.n0 a_809_369.t3 385.062
R246 a_809_369.t1 a_809_369.n3 380.975
R247 a_809_369.n2 a_809_369.t2 321.333
R248 a_809_369.n1 a_809_369.t0 182.711
R249 a_809_369.n0 a_809_369.t5 148.348
R250 a_809_369.n1 a_809_369.n0 117.346
R251 a_809_369.n3 a_809_369.n2 38.615
R252 a_809_369.n3 a_809_369.n1 1.197
R253 a_181_47.n2 a_181_47.n1 481.592
R254 a_181_47.n0 a_181_47.t2 400.951
R255 a_181_47.n3 a_181_47.n2 321.187
R256 a_181_47.n0 a_181_47.t3 196.304
R257 a_181_47.n3 a_181_47.t4 41.554
R258 a_181_47.t1 a_181_47.n3 41.554
R259 a_181_47.n1 a_181_47.t5 38.571
R260 a_181_47.n1 a_181_47.t0 38.571
R261 a_181_47.n2 a_181_47.n0 13.323
R262 a_1129_21.n1 a_1129_21.n0 443.758
R263 a_1129_21.t0 a_1129_21.n2 249.309
R264 a_1129_21.n2 a_1129_21.n1 204.526
R265 a_1129_21.n1 a_1129_21.t3 139.821
R266 a_1129_21.n2 a_1129_21.t4 132.184
R267 a_1129_21.n0 a_1129_21.t2 84.428
R268 a_1129_21.n0 a_1129_21.t1 75.047
R269 a_1347_47.t0 a_1347_47.t1 60
R270 SCE.n0 SCE.t3 293.601
R271 SCE.n1 SCE.t2 292.153
R272 SCE.n1 SCE.t0 227.541
R273 SCE.n0 SCE.t1 202.561
R274 SCE.n2 SCE.n0 12.84
R275 SCE.n2 SCE.n1 8.415
R276 SCE SCE.n2 3.384
R277 a_109_47.t0 a_109_47.t1 60
R278 a_1514_47.t0 a_1514_47.t1 139.687
R279 a_1781_295.n0 a_1781_295.t2 453.613
R280 a_1781_295.n1 a_1781_295.t1 405.297
R281 a_1781_295.t0 a_1781_295.n1 209.699
R282 a_1781_295.n1 a_1781_295.n0 176.552
R283 a_1781_295.n0 a_1781_295.t3 161.201
R284 a_1723_413.t0 a_1723_413.t1 136.023
R285 a_319_21.t1 a_319_21.n1 462.451
R286 a_319_21.n0 a_319_21.t2 283.285
R287 a_319_21.n0 a_319_21.t3 190.099
R288 a_319_21.n1 a_319_21.t0 166.701
R289 a_319_21.n1 a_319_21.n0 76
R290 a_1815_47.t0 a_1815_47.t1 60
R291 D.n0 D.t0 373.281
R292 D.n0 D.t1 132.281
R293 D.n1 D.n0 76
R294 D.n1 D 23.129
R295 D D.n1 7.41
R296 a_193_369.t0 a_193_369.t1 64.64
R297 a_1887_47.t0 a_1887_47.t1 94.285
R298 a_1525_329.t0 a_1525_329.t1 49.25
R299 a_265_47.t0 a_265_47.t1 77.142
R300 a_1087_47.t0 a_1087_47.t1 60
R301 CLK.n0 CLK.t0 255.075
R302 CLK.n0 CLK.t1 218.64
R303 CLK.n1 CLK.n0 76
R304 CLK.n1 CLK 19.069
R305 CLK CLK.n1 2.909
C0 VPWR VGND 0.13fF
C1 VPWR Q 0.12fF
C2 SCE D 0.17fF
C3 VGND Q 0.14fF
C4 SCE VGND 0.16fF
C5 SCE CLK 0.10fF
C6 VPB VPWR 0.25fF
C7 SCD SCE 0.21fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__sdfstp_2.ext - technology: sky130A

.subckt sky130_fd_sc_hd__sdfstp_2 SCD CLK D SET_B SCE Q VPWR VGND VNB VPB
X0 VPWR.t5 a_1597_329.t5 a_2227_47.t1 VPB.t7 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1 VPWR.t2 a_2227_47.t2 Q.t1 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 Q.t3 a_2227_47.t3 VGND.t2 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 a_1597_329.t2 SET_B.t0 VPWR.t10 VPB.t14 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 VPWR.t12 SCD.t0 a_27_369.t1 VPB.t16 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X5 a_1081_413.t0 a_643_369.t2 a_997_413.t1 VPB.t11 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 a_809_369.t1 a_643_369.t3 VGND.t8 VNB.t9 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7 VGND.t4 a_1597_329.t6 a_2227_47.t0 VNB.t5 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 a_997_413.t2 a_809_369.t2 a_181_47.t3 VPB.t19 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9 VPWR.t11 SET_B.t1 a_1129_21.t0 VPB.t15 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10 a_1347_47.t1 a_997_413.t4 a_1129_21.t1 VNB.t7 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11 VPWR.t13 a_1129_21.t3 a_1081_413.t1 VPB.t17 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12 a_181_47.t5 SCE.t0 a_109_47.t0 VNB.t17 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13 a_1514_47.t0 a_997_413.t5 VGND.t7 VNB.t8 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X14 VPWR.t14 a_1781_295.t2 a_1723_413.t0 VPB.t18 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15 VGND.t9 SET_B.t2 a_1347_47.t0 VNB.t12 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16 a_27_369.t0 a_319_21.t2 a_181_47.t1 VPB.t8 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X17 VGND.t3 SCE.t1 a_319_21.t1 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18 a_1597_329.t3 a_809_369.t3 a_1514_47.t1 VNB.t19 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X19 a_1815_47.t1 a_643_369.t4 a_1597_329.t0 VNB.t10 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20 a_181_47.t0 D.t0 a_193_369.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X21 VGND.t10 SET_B.t3 a_1887_47.t1 VNB.t13 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22 a_1597_329.t1 a_643_369.t5 a_1525_329.t1 VPB.t12 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X23 a_265_47.t0 D.t1 a_181_47.t4 VNB.t15 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24 a_997_413.t0 a_643_369.t6 a_181_47.t2 VNB.t11 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X25 VGND.t1 a_2227_47.t4 Q.t2 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X26 Q.t0 a_2227_47.t5 VPWR.t1 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X27 a_1781_295.t1 a_1597_329.t7 VGND.t5 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X28 a_1887_47.t0 a_1781_295.t3 a_1815_47.t0 VNB.t14 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X29 a_1087_47.t1 a_809_369.t4 a_997_413.t3 VNB.t20 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X30 a_193_369.t1 SCE.t2 VPWR.t3 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X31 a_809_369.t0 a_643_369.t7 VPWR.t9 VPB.t13 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X32 a_1525_329.t0 a_997_413.t6 VPWR.t7 VPB.t9 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X33 a_1723_413.t1 a_809_369.t5 a_1597_329.t4 VPB.t20 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X34 VPWR.t4 SCE.t3 a_319_21.t0 VPB.t5 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X35 VPWR.t0 CLK.t0 a_643_369.t1 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X36 a_1129_21.t2 a_997_413.t7 VPWR.t8 VPB.t10 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X37 VGND.t6 a_319_21.t3 a_265_47.t1 VNB.t6 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X38 VGND.t11 a_1129_21.t4 a_1087_47.t0 VNB.t16 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X39 VGND.t0 CLK.t1 a_643_369.t0 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X40 a_1781_295.t0 a_1597_329.t8 VPWR.t6 VPB.t6 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X41 a_109_47.t1 SCD.t1 VGND.t12 VNB.t18 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
R0 a_1597_329.n6 a_1597_329.n5 381.354
R1 a_1597_329.n2 a_1597_329.t6 356.68
R2 a_1597_329.n5 a_1597_329.t2 355.821
R3 a_1597_329.n3 a_1597_329.n2 291.341
R4 a_1597_329.n1 a_1597_329.n0 269.852
R5 a_1597_329.n3 a_1597_329.t8 144.6
R6 a_1597_329.n2 a_1597_329.t5 133.352
R7 a_1597_329.n1 a_1597_329.t7 132.281
R8 a_1597_329.n4 a_1597_329.n1 111.574
R9 a_1597_329.n5 a_1597_329.n4 110.713
R10 a_1597_329.t1 a_1597_329.n6 104.362
R11 a_1597_329.n6 a_1597_329.t4 91.464
R12 a_1597_329.n0 a_1597_329.t0 84.285
R13 a_1597_329.n0 a_1597_329.t3 34.865
R14 a_1597_329.n4 a_1597_329.n3 32.133
R15 a_2227_47.t1 a_2227_47.n2 245.682
R16 a_2227_47.n0 a_2227_47.t2 212.079
R17 a_2227_47.n1 a_2227_47.t5 212.079
R18 a_2227_47.n2 a_2227_47.t0 159.132
R19 a_2227_47.n0 a_2227_47.t4 139.779
R20 a_2227_47.n1 a_2227_47.t3 139.779
R21 a_2227_47.n2 a_2227_47.n1 110.214
R22 a_2227_47.n1 a_2227_47.n0 67.918
R23 VPWR.n45 VPWR.t4 441.584
R24 VPWR.n7 VPWR.t6 370.56
R25 VPWR.n57 VPWR.n56 309.566
R26 VPWR.n12 VPWR.n11 306.463
R27 VPWR.n41 VPWR.n40 306.463
R28 VPWR.n23 VPWR.n22 292.5
R29 VPWR.n29 VPWR.n28 292.5
R30 VPWR.n1 VPWR.n0 172.237
R31 VPWR.n2 VPWR.t2 155.77
R32 VPWR.n28 VPWR.t8 138.369
R33 VPWR.n11 VPWR.t14 126.642
R34 VPWR.n28 VPWR.t13 91.464
R35 VPWR.n11 VPWR.t10 89.119
R36 VPWR.n22 VPWR.t7 87.945
R37 VPWR.n22 VPWR.t11 84.428
R38 VPWR.n0 VPWR.t5 58.484
R39 VPWR.n40 VPWR.t9 41.554
R40 VPWR.n40 VPWR.t0 41.554
R41 VPWR.n56 VPWR.t3 41.554
R42 VPWR.n56 VPWR.t12 41.554
R43 VPWR.n0 VPWR.t1 31.137
R44 VPWR.n4 VPWR.n3 4.65
R45 VPWR.n6 VPWR.n5 4.65
R46 VPWR.n8 VPWR.n7 4.65
R47 VPWR.n10 VPWR.n9 4.65
R48 VPWR.n13 VPWR.n12 4.65
R49 VPWR.n15 VPWR.n14 4.65
R50 VPWR.n17 VPWR.n16 4.65
R51 VPWR.n19 VPWR.n18 4.65
R52 VPWR.n21 VPWR.n20 4.65
R53 VPWR.n25 VPWR.n24 4.65
R54 VPWR.n27 VPWR.n26 4.65
R55 VPWR.n31 VPWR.n30 4.65
R56 VPWR.n33 VPWR.n32 4.65
R57 VPWR.n35 VPWR.n34 4.65
R58 VPWR.n37 VPWR.n36 4.65
R59 VPWR.n39 VPWR.n38 4.65
R60 VPWR.n42 VPWR.n41 4.65
R61 VPWR.n44 VPWR.n43 4.65
R62 VPWR.n47 VPWR.n46 4.65
R63 VPWR.n49 VPWR.n48 4.65
R64 VPWR.n51 VPWR.n50 4.65
R65 VPWR.n53 VPWR.n52 4.65
R66 VPWR.n55 VPWR.n54 4.65
R67 VPWR.n2 VPWR.n1 3.966
R68 VPWR.n58 VPWR.n57 3.932
R69 VPWR.n30 VPWR.n29 2.415
R70 VPWR.n24 VPWR.n23 1.788
R71 VPWR.n46 VPWR.n45 0.376
R72 VPWR.n4 VPWR.n2 0.214
R73 VPWR.n58 VPWR.n55 0.137
R74 VPWR VPWR.n58 0.123
R75 VPWR.n6 VPWR.n4 0.119
R76 VPWR.n8 VPWR.n6 0.119
R77 VPWR.n10 VPWR.n8 0.119
R78 VPWR.n13 VPWR.n10 0.119
R79 VPWR.n15 VPWR.n13 0.119
R80 VPWR.n17 VPWR.n15 0.119
R81 VPWR.n19 VPWR.n17 0.119
R82 VPWR.n21 VPWR.n19 0.119
R83 VPWR.n25 VPWR.n21 0.119
R84 VPWR.n27 VPWR.n25 0.119
R85 VPWR.n31 VPWR.n27 0.119
R86 VPWR.n33 VPWR.n31 0.119
R87 VPWR.n35 VPWR.n33 0.119
R88 VPWR.n37 VPWR.n35 0.119
R89 VPWR.n39 VPWR.n37 0.119
R90 VPWR.n42 VPWR.n39 0.119
R91 VPWR.n44 VPWR.n42 0.119
R92 VPWR.n47 VPWR.n44 0.119
R93 VPWR.n49 VPWR.n47 0.119
R94 VPWR.n51 VPWR.n49 0.119
R95 VPWR.n53 VPWR.n51 0.119
R96 VPWR.n55 VPWR.n53 0.119
R97 VPB.t6 VPB.t7 556.386
R98 VPB.t14 VPB.t6 556.386
R99 VPB.t13 VPB.t19 556.386
R100 VPB.t5 VPB.t1 556.386
R101 VPB.t8 VPB.t5 556.386
R102 VPB.t17 VPB.t10 378.816
R103 VPB.t12 VPB.t20 372.897
R104 VPB.t18 VPB.t14 361.059
R105 VPB.t15 VPB.t9 343.302
R106 VPB.t11 VPB.t17 301.869
R107 VPB.t10 VPB.t15 290.031
R108 VPB.t7 VPB.t2 281.152
R109 VPB.t2 VPB.t3 275.233
R110 VPB.t20 VPB.t18 260.436
R111 VPB.t19 VPB.t11 248.598
R112 VPB.t1 VPB.t13 248.598
R113 VPB.t0 VPB.t8 248.598
R114 VPB.t16 VPB.t4 248.598
R115 VPB.t9 VPB.t12 213.084
R116 VPB.t4 VPB.t0 213.084
R117 VPB VPB.t16 192.367
R118 Q.n2 Q.n1 292.5
R119 Q.n1 Q.n0 147.104
R120 Q Q.n5 95.021
R121 Q.n6 Q.n5 92.5
R122 Q.n1 Q.t0 35.46
R123 Q.n5 Q.t3 33.23
R124 Q.n1 Q.t1 26.595
R125 Q.n5 Q.t2 24.923
R126 Q.n4 Q 16.29
R127 Q.n0 Q 10.71
R128 Q.n6 Q 10.666
R129 Q.n3 Q.n2 6.4
R130 Q.n2 Q 4.848
R131 Q.n4 Q 3.49
R132 Q Q.n3 2.909
R133 Q Q.n6 2.521
R134 Q.n0 Q 2.439
R135 Q Q.n4 2.327
R136 Q.n3 Q 1.939
R137 VGND.n49 VGND.t6 157.996
R138 VGND.n57 VGND.t12 131.071
R139 VGND.n44 VGND.t3 131.071
R140 VGND.n30 VGND.t11 131.071
R141 VGND.n2 VGND.t1 112.461
R142 VGND.n8 VGND.n7 110.932
R143 VGND.n1 VGND.n0 108.12
R144 VGND.n40 VGND.n39 106.463
R145 VGND.n23 VGND.n22 92.5
R146 VGND.n7 VGND.t10 81.428
R147 VGND.n0 VGND.t4 54.285
R148 VGND.n22 VGND.t9 41.428
R149 VGND.n22 VGND.t7 39.151
R150 VGND.n7 VGND.t5 38.571
R151 VGND.n39 VGND.t8 38.571
R152 VGND.n39 VGND.t0 38.571
R153 VGND.n0 VGND.t2 25.934
R154 VGND.n58 VGND.n57 5.214
R155 VGND.n4 VGND.n3 4.65
R156 VGND.n6 VGND.n5 4.65
R157 VGND.n9 VGND.n8 4.65
R158 VGND.n11 VGND.n10 4.65
R159 VGND.n13 VGND.n12 4.65
R160 VGND.n15 VGND.n14 4.65
R161 VGND.n17 VGND.n16 4.65
R162 VGND.n19 VGND.n18 4.65
R163 VGND.n21 VGND.n20 4.65
R164 VGND.n25 VGND.n24 4.65
R165 VGND.n27 VGND.n26 4.65
R166 VGND.n29 VGND.n28 4.65
R167 VGND.n32 VGND.n31 4.65
R168 VGND.n34 VGND.n33 4.65
R169 VGND.n36 VGND.n35 4.65
R170 VGND.n38 VGND.n37 4.65
R171 VGND.n41 VGND.n40 4.65
R172 VGND.n43 VGND.n42 4.65
R173 VGND.n46 VGND.n45 4.65
R174 VGND.n48 VGND.n47 4.65
R175 VGND.n50 VGND.n49 4.65
R176 VGND.n52 VGND.n51 4.65
R177 VGND.n54 VGND.n53 4.65
R178 VGND.n56 VGND.n55 4.65
R179 VGND.n31 VGND.n30 4.189
R180 VGND.n2 VGND.n1 3.897
R181 VGND.n45 VGND.n44 2.8
R182 VGND.n24 VGND.n23 1.582
R183 VGND.n4 VGND.n2 0.224
R184 VGND.n6 VGND.n4 0.119
R185 VGND.n9 VGND.n6 0.119
R186 VGND.n11 VGND.n9 0.119
R187 VGND.n13 VGND.n11 0.119
R188 VGND.n15 VGND.n13 0.119
R189 VGND.n17 VGND.n15 0.119
R190 VGND.n19 VGND.n17 0.119
R191 VGND.n21 VGND.n19 0.119
R192 VGND.n25 VGND.n21 0.119
R193 VGND.n27 VGND.n25 0.119
R194 VGND.n29 VGND.n27 0.119
R195 VGND.n32 VGND.n29 0.119
R196 VGND.n34 VGND.n32 0.119
R197 VGND.n36 VGND.n34 0.119
R198 VGND.n38 VGND.n36 0.119
R199 VGND.n41 VGND.n38 0.119
R200 VGND.n43 VGND.n41 0.119
R201 VGND.n46 VGND.n43 0.119
R202 VGND.n48 VGND.n46 0.119
R203 VGND.n50 VGND.n48 0.119
R204 VGND.n52 VGND.n50 0.119
R205 VGND.n54 VGND.n52 0.119
R206 VGND.n56 VGND.n54 0.119
R207 VGND.n58 VGND.n56 0.119
R208 VGND VGND.n58 0.022
R209 VNB.t4 VNB.t5 6858.82
R210 VNB VNB.t18 6470.59
R211 VNB.t6 VNB.t3 6276.47
R212 VNB.t16 VNB.t7 6082.35
R213 VNB.t9 VNB.t11 6082.35
R214 VNB.t3 VNB.t0 6082.35
R215 VNB.t8 VNB.t19 4375.56
R216 VNB.t13 VNB.t4 3688.24
R217 VNB.t19 VNB.t10 3227.39
R218 VNB.t14 VNB.t13 3105.88
R219 VNB.t11 VNB.t20 2717.65
R220 VNB.t0 VNB.t9 2717.65
R221 VNB.t15 VNB.t6 2717.65
R222 VNB.t17 VNB.t15 2717.65
R223 VNB.t10 VNB.t14 2329.41
R224 VNB.t7 VNB.t12 2329.41
R225 VNB.t20 VNB.t16 2329.41
R226 VNB.t18 VNB.t17 2329.41
R227 VNB.t12 VNB.t8 2280.14
R228 VNB.t5 VNB.t2 2255.35
R229 VNB.t2 VNB.t1 2248.35
R230 SET_B.n0 SET_B.t2 360.179
R231 SET_B.n1 SET_B.t3 357.215
R232 SET_B.n0 SET_B.t1 166.576
R233 SET_B.n1 SET_B.t0 161.029
R234 SET_B.n2 SET_B.n1 137.809
R235 SET_B.n2 SET_B.n0 83
R236 SET_B SET_B.n2 3.4
R237 SCD.n0 SCD.t0 299.43
R238 SCD.n0 SCD.t1 206.244
R239 SCD.n1 SCD.n0 76
R240 SCD.n1 SCD 19.827
R241 SCD SCD.n1 14.305
R242 a_27_369.t0 a_27_369.t1 883.735
R243 a_643_369.n2 a_643_369.t6 393.633
R244 a_643_369.t1 a_643_369.n5 377.811
R245 a_643_369.n0 a_643_369.t5 343.241
R246 a_643_369.n0 a_643_369.t4 337.584
R247 a_643_369.n3 a_643_369.t7 267.297
R248 a_643_369.n4 a_643_369.t0 199.461
R249 a_643_369.n1 a_643_369.t2 147.521
R250 a_643_369.n3 a_643_369.n2 100.205
R251 a_643_369.n2 a_643_369.t3 91.58
R252 a_643_369.n4 a_643_369.n3 76
R253 a_643_369.n1 a_643_369.n0 49.157
R254 a_643_369.n5 a_643_369.n4 30.276
R255 a_643_369.n5 a_643_369.n1 5.776
R256 a_997_413.n4 a_997_413.n0 369.55
R257 a_997_413.n1 a_997_413.t7 312.131
R258 a_997_413.n2 a_997_413.t6 262.639
R259 a_997_413.n1 a_997_413.t4 238.224
R260 a_997_413.n2 a_997_413.t5 166.239
R261 a_997_413.n5 a_997_413.n4 141.906
R262 a_997_413.n3 a_997_413.n2 124.559
R263 a_997_413.n3 a_997_413.n1 76
R264 a_997_413.n0 a_997_413.t1 63.321
R265 a_997_413.n0 a_997_413.t2 63.321
R266 a_997_413.n4 a_997_413.n3 53.834
R267 a_997_413.n5 a_997_413.t3 38.571
R268 a_997_413.t0 a_997_413.n5 38.571
R269 a_1081_413.t0 a_1081_413.t1 168.857
R270 a_809_369.n2 a_809_369.t4 433.507
R271 a_809_369.n0 a_809_369.t3 385.062
R272 a_809_369.t0 a_809_369.n3 380.975
R273 a_809_369.n2 a_809_369.t2 321.333
R274 a_809_369.n1 a_809_369.t1 182.711
R275 a_809_369.n0 a_809_369.t5 148.348
R276 a_809_369.n1 a_809_369.n0 117.346
R277 a_809_369.n3 a_809_369.n2 38.615
R278 a_809_369.n3 a_809_369.n1 1.197
R279 a_181_47.n2 a_181_47.n1 481.592
R280 a_181_47.n0 a_181_47.t3 400.951
R281 a_181_47.n3 a_181_47.n2 321.187
R282 a_181_47.n0 a_181_47.t2 196.304
R283 a_181_47.n3 a_181_47.t1 41.554
R284 a_181_47.t0 a_181_47.n3 41.554
R285 a_181_47.n1 a_181_47.t4 38.571
R286 a_181_47.n1 a_181_47.t5 38.571
R287 a_181_47.n2 a_181_47.n0 13.323
R288 a_1129_21.n2 a_1129_21.n1 443.758
R289 a_1129_21.n0 a_1129_21.t1 249.309
R290 a_1129_21.n1 a_1129_21.n0 204.526
R291 a_1129_21.n1 a_1129_21.t3 139.821
R292 a_1129_21.n0 a_1129_21.t4 132.184
R293 a_1129_21.t0 a_1129_21.n2 84.428
R294 a_1129_21.n2 a_1129_21.t2 75.047
R295 a_1347_47.t0 a_1347_47.t1 60
R296 SCE.n0 SCE.t3 293.601
R297 SCE.n1 SCE.t2 292.153
R298 SCE.n1 SCE.t0 227.541
R299 SCE.n0 SCE.t1 202.561
R300 SCE.n2 SCE.n0 12.84
R301 SCE.n2 SCE.n1 8.415
R302 SCE SCE.n2 3.384
R303 a_109_47.t0 a_109_47.t1 60
R304 a_1514_47.t0 a_1514_47.t1 139.687
R305 a_1781_295.n0 a_1781_295.t2 453.613
R306 a_1781_295.t0 a_1781_295.n1 405.297
R307 a_1781_295.n1 a_1781_295.t1 209.699
R308 a_1781_295.n1 a_1781_295.n0 176.552
R309 a_1781_295.n0 a_1781_295.t3 161.201
R310 a_1723_413.t0 a_1723_413.t1 136.023
R311 a_319_21.t0 a_319_21.n1 462.451
R312 a_319_21.n0 a_319_21.t2 283.285
R313 a_319_21.n0 a_319_21.t3 190.099
R314 a_319_21.n1 a_319_21.t1 166.701
R315 a_319_21.n1 a_319_21.n0 76
R316 a_1815_47.t0 a_1815_47.t1 60
R317 D.n0 D.t0 373.281
R318 D.n0 D.t1 132.281
R319 D.n1 D.n0 76
R320 D.n1 D 23.129
R321 D D.n1 7.41
R322 a_193_369.t0 a_193_369.t1 64.64
R323 a_1887_47.t0 a_1887_47.t1 94.285
R324 a_1525_329.t0 a_1525_329.t1 49.25
R325 a_265_47.t0 a_265_47.t1 77.142
R326 a_1087_47.t0 a_1087_47.t1 60
R327 CLK.n0 CLK.t0 255.075
R328 CLK.n0 CLK.t1 218.64
R329 CLK.n1 CLK.n0 76
R330 CLK.n1 CLK 19.069
R331 CLK CLK.n1 2.909
C0 VPWR VGND 0.16fF
C1 VPWR Q 0.29fF
C2 SCE D 0.17fF
C3 VGND Q 0.25fF
C4 SCE VGND 0.16fF
C5 VPB VPWR 0.26fF
C6 SCE CLK 0.10fF
C7 SCD SCE 0.21fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__sdfstp_4.ext - technology: sky130A

.subckt sky130_fd_sc_hd__sdfstp_4 CLK D SCE SET_B SCD Q VPWR VGND VNB VPB
X0 VPWR.t12 a_2227_47.t2 Q.t3 VPB.t17 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 Q.t7 a_2227_47.t3 VGND.t10 VNB.t18 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 a_1597_329.t0 SET_B.t0 VPWR.t15 VPB.t20 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3 Q.t2 a_2227_47.t4 VPWR.t11 VPB.t16 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 VPWR.t7 SCD.t0 a_27_369.t0 VPB.t12 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X5 a_1081_413.t1 a_643_369.t2 a_997_413.t2 VPB.t9 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 a_809_369.t1 a_643_369.t3 VGND.t5 VNB.t11 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7 VGND.t11 a_1597_329.t5 a_2227_47.t0 VNB.t19 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 a_997_413.t0 a_809_369.t2 a_181_47.t0 VPB.t7 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9 VPWR.t16 SET_B.t1 a_1129_21.t0 VPB.t21 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10 a_1347_47.t1 a_997_413.t4 a_1129_21.t2 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11 VPWR.t0 a_1129_21.t3 a_1081_413.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12 a_181_47.t3 SCE.t0 a_109_47.t1 VNB.t10 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13 a_1514_47.t1 a_997_413.t5 VGND.t2 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X14 Q.t6 a_2227_47.t5 VGND.t9 VNB.t17 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X15 VPWR.t8 a_1781_295.t2 a_1723_413.t1 VPB.t13 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16 VGND.t8 a_2227_47.t6 Q.t5 VNB.t16 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X17 VGND.t13 SET_B.t2 a_1347_47.t0 VNB.t21 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18 a_27_369.t1 a_319_21.t2 a_181_47.t5 VPB.t22 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X19 VGND.t4 SCE.t1 a_319_21.t1 VNB.t6 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20 a_1597_329.t1 a_809_369.t3 a_1514_47.t0 VNB.t7 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X21 a_1815_47.t1 a_643_369.t4 a_1597_329.t3 VNB.t12 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22 a_181_47.t1 D.t0 a_193_369.t0 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X23 VPWR.t10 a_2227_47.t7 Q.t1 VPB.t15 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X24 VGND.t14 SET_B.t3 a_1887_47.t1 VNB.t22 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X25 VGND.t7 a_2227_47.t8 Q.t4 VNB.t15 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X26 a_1597_329.t4 a_643_369.t5 a_1525_329.t1 VPB.t10 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X27 a_265_47.t1 D.t1 a_181_47.t2 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X28 a_997_413.t3 a_643_369.t6 a_181_47.t4 VNB.t13 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X29 Q.t0 a_2227_47.t9 VPWR.t9 VPB.t14 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X30 a_1781_295.t1 a_1597_329.t6 VGND.t12 VNB.t20 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X31 a_1887_47.t0 a_1781_295.t3 a_1815_47.t0 VNB.t9 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X32 a_1087_47.t0 a_809_369.t4 a_997_413.t1 VNB.t8 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X33 a_193_369.t1 SCE.t2 VPWR.t4 VPB.t5 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X34 a_809_369.t0 a_643_369.t7 VPWR.t6 VPB.t11 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X35 a_1525_329.t0 a_997_413.t6 VPWR.t2 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X36 a_1723_413.t0 a_809_369.t5 a_1597_329.t2 VPB.t8 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X37 VPWR.t5 SCE.t3 a_319_21.t0 VPB.t6 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X38 VPWR.t13 a_1597_329.t7 a_2227_47.t1 VPB.t18 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X39 VPWR.t1 CLK.t0 a_643_369.t1 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X40 a_1129_21.t1 a_997_413.t7 VPWR.t3 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X41 VGND.t3 a_319_21.t3 a_265_47.t0 VNB.t5 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X42 VGND.t1 a_1129_21.t4 a_1087_47.t1 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X43 VGND.t0 CLK.t1 a_643_369.t0 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X44 a_1781_295.t0 a_1597_329.t8 VPWR.t14 VPB.t19 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X45 a_109_47.t0 SCD.t1 VGND.t6 VNB.t14 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
R0 a_2227_47.n0 a_2227_47.t2 212.079
R1 a_2227_47.n1 a_2227_47.t4 212.079
R2 a_2227_47.n2 a_2227_47.t7 212.079
R3 a_2227_47.n3 a_2227_47.t9 212.079
R4 a_2227_47.t1 a_2227_47.n4 207.93
R5 a_2227_47.n4 a_2227_47.t0 145.484
R6 a_2227_47.n0 a_2227_47.t8 139.779
R7 a_2227_47.n1 a_2227_47.t5 139.779
R8 a_2227_47.n2 a_2227_47.t6 139.779
R9 a_2227_47.n3 a_2227_47.t3 139.779
R10 a_2227_47.n4 a_2227_47.n3 110.214
R11 a_2227_47.n2 a_2227_47.n1 68.648
R12 a_2227_47.n1 a_2227_47.n0 61.345
R13 a_2227_47.n3 a_2227_47.n2 61.345
R14 Q Q.n7 298.706
R15 Q.n5 Q.n3 123.344
R16 Q.n1 Q.n0 92.5
R17 Q.n5 Q.n4 68.334
R18 Q.n7 Q.t1 26.595
R19 Q.n7 Q.t0 26.595
R20 Q.n3 Q.t3 26.595
R21 Q.n3 Q.t2 26.595
R22 Q.n0 Q.t5 24.923
R23 Q.n0 Q.t7 24.923
R24 Q.n4 Q.t4 24.923
R25 Q.n4 Q.t6 24.923
R26 Q.n6 Q 19.2
R27 Q.n6 Q.n2 13.084
R28 Q Q.n1 12.606
R29 Q.n8 Q 11.248
R30 Q Q.n5 10.429
R31 Q Q.n6 6.826
R32 Q.n2 Q 3.413
R33 Q.n8 Q 2.844
R34 Q.n6 Q 2.607
R35 Q.n2 Q 2.327
R36 Q Q.n8 1.939
R37 Q.n1 Q 0.581
R38 VPWR.n50 VPWR.t5 441.584
R39 VPWR.n12 VPWR.t14 370.56
R40 VPWR.n62 VPWR.n61 309.566
R41 VPWR.n17 VPWR.n16 306.463
R42 VPWR.n46 VPWR.n45 306.463
R43 VPWR.n28 VPWR.n27 292.5
R44 VPWR.n34 VPWR.n33 292.5
R45 VPWR.n2 VPWR.t12 149.562
R46 VPWR.n33 VPWR.t3 138.369
R47 VPWR.n1 VPWR.n0 132.865
R48 VPWR.n16 VPWR.t8 126.642
R49 VPWR.n6 VPWR.n5 117.036
R50 VPWR.n33 VPWR.t0 91.464
R51 VPWR.n16 VPWR.t15 89.119
R52 VPWR.n27 VPWR.t2 87.945
R53 VPWR.n27 VPWR.t16 84.428
R54 VPWR.n45 VPWR.t6 41.554
R55 VPWR.n45 VPWR.t1 41.554
R56 VPWR.n61 VPWR.t4 41.554
R57 VPWR.n61 VPWR.t7 41.554
R58 VPWR.n0 VPWR.t10 36.445
R59 VPWR.n5 VPWR.t9 32.505
R60 VPWR.n5 VPWR.t13 31.52
R61 VPWR.n0 VPWR.t11 26.595
R62 VPWR.n2 VPWR.n1 5.941
R63 VPWR.n4 VPWR.n3 4.65
R64 VPWR.n7 VPWR.n6 4.65
R65 VPWR.n9 VPWR.n8 4.65
R66 VPWR.n11 VPWR.n10 4.65
R67 VPWR.n13 VPWR.n12 4.65
R68 VPWR.n15 VPWR.n14 4.65
R69 VPWR.n18 VPWR.n17 4.65
R70 VPWR.n20 VPWR.n19 4.65
R71 VPWR.n22 VPWR.n21 4.65
R72 VPWR.n24 VPWR.n23 4.65
R73 VPWR.n26 VPWR.n25 4.65
R74 VPWR.n30 VPWR.n29 4.65
R75 VPWR.n32 VPWR.n31 4.65
R76 VPWR.n36 VPWR.n35 4.65
R77 VPWR.n38 VPWR.n37 4.65
R78 VPWR.n40 VPWR.n39 4.65
R79 VPWR.n42 VPWR.n41 4.65
R80 VPWR.n44 VPWR.n43 4.65
R81 VPWR.n47 VPWR.n46 4.65
R82 VPWR.n49 VPWR.n48 4.65
R83 VPWR.n52 VPWR.n51 4.65
R84 VPWR.n54 VPWR.n53 4.65
R85 VPWR.n56 VPWR.n55 4.65
R86 VPWR.n58 VPWR.n57 4.65
R87 VPWR.n60 VPWR.n59 4.65
R88 VPWR.n63 VPWR.n62 3.932
R89 VPWR.n35 VPWR.n34 2.415
R90 VPWR.n29 VPWR.n28 1.788
R91 VPWR.n51 VPWR.n50 0.376
R92 VPWR.n4 VPWR.n2 0.213
R93 VPWR.n63 VPWR.n60 0.137
R94 VPWR VPWR.n63 0.123
R95 VPWR.n7 VPWR.n4 0.119
R96 VPWR.n9 VPWR.n7 0.119
R97 VPWR.n11 VPWR.n9 0.119
R98 VPWR.n13 VPWR.n11 0.119
R99 VPWR.n15 VPWR.n13 0.119
R100 VPWR.n18 VPWR.n15 0.119
R101 VPWR.n20 VPWR.n18 0.119
R102 VPWR.n22 VPWR.n20 0.119
R103 VPWR.n24 VPWR.n22 0.119
R104 VPWR.n26 VPWR.n24 0.119
R105 VPWR.n30 VPWR.n26 0.119
R106 VPWR.n32 VPWR.n30 0.119
R107 VPWR.n36 VPWR.n32 0.119
R108 VPWR.n38 VPWR.n36 0.119
R109 VPWR.n40 VPWR.n38 0.119
R110 VPWR.n42 VPWR.n40 0.119
R111 VPWR.n44 VPWR.n42 0.119
R112 VPWR.n47 VPWR.n44 0.119
R113 VPWR.n49 VPWR.n47 0.119
R114 VPWR.n52 VPWR.n49 0.119
R115 VPWR.n54 VPWR.n52 0.119
R116 VPWR.n56 VPWR.n54 0.119
R117 VPWR.n58 VPWR.n56 0.119
R118 VPWR.n60 VPWR.n58 0.119
R119 VPB.t19 VPB.t18 556.386
R120 VPB.t20 VPB.t19 556.386
R121 VPB.t11 VPB.t7 556.386
R122 VPB.t6 VPB.t1 556.386
R123 VPB.t22 VPB.t6 556.386
R124 VPB.t0 VPB.t4 378.816
R125 VPB.t10 VPB.t8 372.897
R126 VPB.t13 VPB.t20 361.059
R127 VPB.t21 VPB.t3 343.302
R128 VPB.t9 VPB.t0 301.869
R129 VPB.t4 VPB.t21 290.031
R130 VPB.t18 VPB.t14 281.152
R131 VPB.t15 VPB.t16 278.193
R132 VPB.t8 VPB.t13 260.436
R133 VPB.t16 VPB.t17 248.598
R134 VPB.t14 VPB.t15 248.598
R135 VPB.t7 VPB.t9 248.598
R136 VPB.t1 VPB.t11 248.598
R137 VPB.t2 VPB.t22 248.598
R138 VPB.t12 VPB.t5 248.598
R139 VPB.t3 VPB.t10 213.084
R140 VPB.t5 VPB.t2 213.084
R141 VPB VPB.t12 192.367
R142 VGND.n54 VGND.t3 157.996
R143 VGND.n62 VGND.t6 131.071
R144 VGND.n49 VGND.t4 131.071
R145 VGND.n35 VGND.t1 131.071
R146 VGND.n13 VGND.n12 110.932
R147 VGND.n2 VGND.t7 107.255
R148 VGND.n45 VGND.n44 106.463
R149 VGND.n28 VGND.n27 92.5
R150 VGND.n12 VGND.t14 81.428
R151 VGND.n1 VGND.n0 74.084
R152 VGND.n6 VGND.n5 62.105
R153 VGND.n27 VGND.t13 41.428
R154 VGND.n27 VGND.t2 39.151
R155 VGND.n12 VGND.t12 38.571
R156 VGND.n44 VGND.t5 38.571
R157 VGND.n44 VGND.t0 38.571
R158 VGND.n0 VGND.t8 34.153
R159 VGND.n5 VGND.t10 30.461
R160 VGND.n5 VGND.t11 29.538
R161 VGND.n0 VGND.t9 24.923
R162 VGND.n2 VGND.n1 5.941
R163 VGND.n63 VGND.n62 5.214
R164 VGND.n4 VGND.n3 4.65
R165 VGND.n7 VGND.n6 4.65
R166 VGND.n9 VGND.n8 4.65
R167 VGND.n11 VGND.n10 4.65
R168 VGND.n14 VGND.n13 4.65
R169 VGND.n16 VGND.n15 4.65
R170 VGND.n18 VGND.n17 4.65
R171 VGND.n20 VGND.n19 4.65
R172 VGND.n22 VGND.n21 4.65
R173 VGND.n24 VGND.n23 4.65
R174 VGND.n26 VGND.n25 4.65
R175 VGND.n30 VGND.n29 4.65
R176 VGND.n32 VGND.n31 4.65
R177 VGND.n34 VGND.n33 4.65
R178 VGND.n37 VGND.n36 4.65
R179 VGND.n39 VGND.n38 4.65
R180 VGND.n41 VGND.n40 4.65
R181 VGND.n43 VGND.n42 4.65
R182 VGND.n46 VGND.n45 4.65
R183 VGND.n48 VGND.n47 4.65
R184 VGND.n51 VGND.n50 4.65
R185 VGND.n53 VGND.n52 4.65
R186 VGND.n55 VGND.n54 4.65
R187 VGND.n57 VGND.n56 4.65
R188 VGND.n59 VGND.n58 4.65
R189 VGND.n61 VGND.n60 4.65
R190 VGND.n36 VGND.n35 4.189
R191 VGND.n50 VGND.n49 2.8
R192 VGND.n29 VGND.n28 1.582
R193 VGND.n4 VGND.n2 0.212
R194 VGND.n7 VGND.n4 0.119
R195 VGND.n9 VGND.n7 0.119
R196 VGND.n11 VGND.n9 0.119
R197 VGND.n14 VGND.n11 0.119
R198 VGND.n16 VGND.n14 0.119
R199 VGND.n18 VGND.n16 0.119
R200 VGND.n20 VGND.n18 0.119
R201 VGND.n22 VGND.n20 0.119
R202 VGND.n24 VGND.n22 0.119
R203 VGND.n26 VGND.n24 0.119
R204 VGND.n30 VGND.n26 0.119
R205 VGND.n32 VGND.n30 0.119
R206 VGND.n34 VGND.n32 0.119
R207 VGND.n37 VGND.n34 0.119
R208 VGND.n39 VGND.n37 0.119
R209 VGND.n41 VGND.n39 0.119
R210 VGND.n43 VGND.n41 0.119
R211 VGND.n46 VGND.n43 0.119
R212 VGND.n48 VGND.n46 0.119
R213 VGND.n51 VGND.n48 0.119
R214 VGND.n53 VGND.n51 0.119
R215 VGND.n55 VGND.n53 0.119
R216 VGND.n57 VGND.n55 0.119
R217 VGND.n59 VGND.n57 0.119
R218 VGND.n61 VGND.n59 0.119
R219 VGND.n63 VGND.n61 0.119
R220 VGND VGND.n63 0.022
R221 VNB VNB.t14 6470.59
R222 VNB.t5 VNB.t6 6276.47
R223 VNB.t20 VNB.t19 6098.35
R224 VNB.t1 VNB.t2 6082.35
R225 VNB.t11 VNB.t13 6082.35
R226 VNB.t6 VNB.t0 6082.35
R227 VNB.t3 VNB.t7 4375.56
R228 VNB.t22 VNB.t20 3688.24
R229 VNB.t7 VNB.t12 3227.39
R230 VNB.t9 VNB.t22 3105.88
R231 VNB.t13 VNB.t8 2717.65
R232 VNB.t0 VNB.t11 2717.65
R233 VNB.t4 VNB.t5 2717.65
R234 VNB.t10 VNB.t4 2717.65
R235 VNB.t12 VNB.t9 2329.41
R236 VNB.t2 VNB.t21 2329.41
R237 VNB.t8 VNB.t1 2329.41
R238 VNB.t14 VNB.t10 2329.41
R239 VNB.t19 VNB.t18 2296.7
R240 VNB.t21 VNB.t3 2280.14
R241 VNB.t16 VNB.t17 2272.53
R242 VNB.t17 VNB.t15 2030.77
R243 VNB.t18 VNB.t16 2030.77
R244 SET_B.n0 SET_B.t2 360.179
R245 SET_B.n1 SET_B.t3 357.215
R246 SET_B.n0 SET_B.t1 166.576
R247 SET_B.n1 SET_B.t0 161.029
R248 SET_B.n2 SET_B.n1 137.809
R249 SET_B.n2 SET_B.n0 83
R250 SET_B SET_B.n2 3.4
R251 a_1597_329.n6 a_1597_329.n5 381.354
R252 a_1597_329.n5 a_1597_329.t0 355.821
R253 a_1597_329.n3 a_1597_329.n0 277.953
R254 a_1597_329.n2 a_1597_329.n1 269.852
R255 a_1597_329.n0 a_1597_329.t5 207.259
R256 a_1597_329.n0 a_1597_329.t7 202.439
R257 a_1597_329.n4 a_1597_329.t8 161.284
R258 a_1597_329.n2 a_1597_329.t6 132.281
R259 a_1597_329.n5 a_1597_329.n4 105.358
R260 a_1597_329.t4 a_1597_329.n6 104.362
R261 a_1597_329.n6 a_1597_329.t2 91.464
R262 a_1597_329.n1 a_1597_329.t3 84.285
R263 a_1597_329.n3 a_1597_329.n2 58.361
R264 a_1597_329.n4 a_1597_329.n3 50.671
R265 a_1597_329.n1 a_1597_329.t1 34.865
R266 SCD.n0 SCD.t0 299.43
R267 SCD.n0 SCD.t1 206.244
R268 SCD.n1 SCD.n0 76
R269 SCD SCD.n1 19.827
R270 SCD.n1 SCD 14.305
R271 a_27_369.t0 a_27_369.t1 883.735
R272 a_643_369.n2 a_643_369.t6 393.633
R273 a_643_369.t1 a_643_369.n5 377.811
R274 a_643_369.n0 a_643_369.t5 343.241
R275 a_643_369.n0 a_643_369.t4 337.584
R276 a_643_369.n3 a_643_369.t7 267.297
R277 a_643_369.n4 a_643_369.t0 199.461
R278 a_643_369.n1 a_643_369.t2 147.521
R279 a_643_369.n3 a_643_369.n2 100.205
R280 a_643_369.n2 a_643_369.t3 91.58
R281 a_643_369.n4 a_643_369.n3 76
R282 a_643_369.n1 a_643_369.n0 49.157
R283 a_643_369.n5 a_643_369.n4 30.276
R284 a_643_369.n5 a_643_369.n1 5.776
R285 a_997_413.n5 a_997_413.n4 369.55
R286 a_997_413.n0 a_997_413.t7 312.131
R287 a_997_413.n1 a_997_413.t6 262.639
R288 a_997_413.n0 a_997_413.t4 238.224
R289 a_997_413.n1 a_997_413.t5 166.239
R290 a_997_413.n4 a_997_413.n3 141.906
R291 a_997_413.n2 a_997_413.n1 124.559
R292 a_997_413.n2 a_997_413.n0 76
R293 a_997_413.n5 a_997_413.t2 63.321
R294 a_997_413.t0 a_997_413.n5 63.321
R295 a_997_413.n4 a_997_413.n2 53.834
R296 a_997_413.n3 a_997_413.t1 38.571
R297 a_997_413.n3 a_997_413.t3 38.571
R298 a_1081_413.t0 a_1081_413.t1 168.857
R299 a_809_369.n2 a_809_369.t4 433.507
R300 a_809_369.n0 a_809_369.t3 385.062
R301 a_809_369.t0 a_809_369.n3 380.975
R302 a_809_369.n2 a_809_369.t2 321.333
R303 a_809_369.n1 a_809_369.t1 182.711
R304 a_809_369.n0 a_809_369.t5 148.348
R305 a_809_369.n1 a_809_369.n0 117.346
R306 a_809_369.n3 a_809_369.n2 38.615
R307 a_809_369.n3 a_809_369.n1 1.197
R308 a_181_47.n2 a_181_47.n1 481.592
R309 a_181_47.n0 a_181_47.t0 400.951
R310 a_181_47.n3 a_181_47.n2 321.187
R311 a_181_47.n0 a_181_47.t4 196.304
R312 a_181_47.n3 a_181_47.t5 41.554
R313 a_181_47.t1 a_181_47.n3 41.554
R314 a_181_47.n1 a_181_47.t2 38.571
R315 a_181_47.n1 a_181_47.t3 38.571
R316 a_181_47.n2 a_181_47.n0 13.323
R317 a_1129_21.n2 a_1129_21.n1 443.758
R318 a_1129_21.n0 a_1129_21.t2 249.309
R319 a_1129_21.n1 a_1129_21.n0 204.526
R320 a_1129_21.n1 a_1129_21.t3 139.821
R321 a_1129_21.n0 a_1129_21.t4 132.184
R322 a_1129_21.t0 a_1129_21.n2 84.428
R323 a_1129_21.n2 a_1129_21.t1 75.047
R324 a_1347_47.t0 a_1347_47.t1 60
R325 SCE.n0 SCE.t3 293.601
R326 SCE.n1 SCE.t2 292.153
R327 SCE.n1 SCE.t0 227.541
R328 SCE.n0 SCE.t1 202.561
R329 SCE.n2 SCE.n0 12.84
R330 SCE.n2 SCE.n1 8.415
R331 SCE SCE.n2 3.384
R332 a_109_47.t0 a_109_47.t1 60
R333 a_1514_47.t0 a_1514_47.t1 139.687
R334 a_1781_295.n0 a_1781_295.t2 453.613
R335 a_1781_295.t0 a_1781_295.n1 405.297
R336 a_1781_295.n1 a_1781_295.t1 209.699
R337 a_1781_295.n1 a_1781_295.n0 176.552
R338 a_1781_295.n0 a_1781_295.t3 161.201
R339 a_1723_413.t0 a_1723_413.t1 136.023
R340 a_319_21.t0 a_319_21.n1 462.451
R341 a_319_21.n0 a_319_21.t2 283.285
R342 a_319_21.n0 a_319_21.t3 190.099
R343 a_319_21.n1 a_319_21.t1 166.701
R344 a_319_21.n1 a_319_21.n0 76
R345 a_1815_47.t0 a_1815_47.t1 60
R346 D.n0 D.t0 373.281
R347 D.n0 D.t1 132.281
R348 D.n1 D.n0 76
R349 D D.n1 23.129
R350 D.n1 D 7.41
R351 a_193_369.t0 a_193_369.t1 64.64
R352 a_1887_47.t0 a_1887_47.t1 94.285
R353 a_1525_329.t0 a_1525_329.t1 49.25
R354 a_265_47.t0 a_265_47.t1 77.142
R355 a_1087_47.t0 a_1087_47.t1 60
R356 CLK.n0 CLK.t0 255.075
R357 CLK.n0 CLK.t1 218.64
R358 CLK.n1 CLK.n0 76
R359 CLK.n1 CLK 19.069
R360 CLK CLK.n1 2.909
C0 VPWR VGND 0.19fF
C1 VPWR Q 0.66fF
C2 SCE D 0.17fF
C3 VGND Q 0.47fF
C4 SCE VGND 0.16fF
C5 VPB VPWR 0.28fF
C6 SCE CLK 0.10fF
C7 SCD SCE 0.21fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__sdfxbp_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__sdfxbp_1 VGND VPWR SCD Q_N D SCE CLK Q VNB VPB
X0 a_640_369.t0 a_299_47.t2 a_556_369.t2 VPB.t6 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1 VPWR.t1 SCE.t0 a_299_47.t1 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X2 a_556_369.t5 D.t0 a_465_369.t1 VPB.t17 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X3 a_1089_183.t1 a_930_413.t4 VPWR.t4 VPB.t7 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X4 a_1430_413.t0 a_193_47.t2 a_1346_413.t2 VPB.t15 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 Q.t1 a_1517_315.t2 VGND.t8 VNB.t14 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 Q_N.t1 a_1948_47.t2 VGND.t10 VNB.t16 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 VPWR.t3 CLK.t0 a_27_47.t0 VPB.t5 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X8 a_1346_413.t1 a_27_47.t2 a_1089_183.t0 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9 a_1089_183.t2 a_930_413.t5 VGND.t3 VNB.t7 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X10 a_657_47.t0 SCE.t1 a_556_369.t0 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11 VGND.t5 a_1346_413.t4 a_1517_315.t1 VNB.t11 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 a_930_413.t1 a_27_47.t3 a_556_369.t1 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X13 VPWR.t6 SCD.t0 a_640_369.t1 VPB.t9 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X14 a_193_47.t1 a_27_47.t4 VGND.t0 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15 a_483_47.t1 a_299_47.t3 VGND.t4 VNB.t10 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16 VGND.t9 a_1089_183.t4 a_1027_47.t1 VNB.t15 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17 a_930_413.t2 a_193_47.t3 a_556_369.t4 VPB.t16 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18 Q_N.t0 a_1948_47.t3 VPWR.t7 VPB.t10 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X19 VGND.t6 a_1517_315.t3 a_1475_47.t1 VNB.t13 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20 Q.t0 a_1517_315.t4 VPWR.t8 VPB.t11 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X21 a_1475_47.t0 a_27_47.t5 a_1346_413.t0 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X22 VPWR.t5 a_1346_413.t5 a_1517_315.t0 VPB.t8 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X23 a_193_47.t0 a_27_47.t6 VPWR.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X24 a_1023_413.t0 a_27_47.t7 a_930_413.t0 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X25 VGND.t7 a_1517_315.t5 a_1948_47.t1 VNB.t12 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X26 VPWR.t11 a_1517_315.t6 a_1430_413.t1 VPB.t14 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X27 a_1027_47.t0 a_193_47.t4 a_930_413.t3 VNB.t9 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X28 VGND.t1 SCE.t2 a_299_47.t0 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X29 VGND.t2 SCD.t1 a_657_47.t1 VNB.t5 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X30 VPWR.t9 a_1089_183.t5 a_1023_413.t1 VPB.t12 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X31 VPWR.t10 a_1517_315.t7 a_1948_47.t0 VPB.t13 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X32 a_465_369.t0 SCE.t3 VPWR.t2 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X33 VGND.t11 CLK.t1 a_27_47.t1 VNB.t17 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X34 a_556_369.t3 D.t1 a_483_47.t0 VNB.t6 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X35 a_1346_413.t3 a_193_47.t5 a_1089_183.t3 VNB.t8 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
R0 a_299_47.t1 a_299_47.n1 343.485
R1 a_299_47.n0 a_299_47.t2 340.853
R2 a_299_47.n0 a_299_47.t3 306.024
R3 a_299_47.n1 a_299_47.t0 239.196
R4 a_299_47.n1 a_299_47.n0 28.576
R5 a_556_369.n3 a_556_369.n2 411.84
R6 a_556_369.n2 a_556_369.t4 370.675
R7 a_556_369.n1 a_556_369.n0 207.322
R8 a_556_369.n1 a_556_369.t1 165.247
R9 a_556_369.n2 a_556_369.n1 70.776
R10 a_556_369.n0 a_556_369.t3 54.285
R11 a_556_369.t2 a_556_369.n3 41.554
R12 a_556_369.n3 a_556_369.t5 41.554
R13 a_556_369.n0 a_556_369.t0 40
R14 a_640_369.t0 a_640_369.t1 96.96
R15 VPB.t14 VPB.t8 624.454
R16 VPB.t9 VPB.t16 583.021
R17 VPB.t11 VPB.t13 556.386
R18 VPB.t0 VPB.t3 556.386
R19 VPB.t12 VPB.t7 390.654
R20 VPB.t15 VPB.t14 346.261
R21 VPB.t13 VPB.t10 287.071
R22 VPB.t1 VPB.t12 284.112
R23 VPB.t7 VPB.t2 281.152
R24 VPB.t16 VPB.t1 275.233
R25 VPB.t6 VPB.t9 275.233
R26 VPB.t4 VPB.t17 269.314
R27 VPB.t8 VPB.t11 248.598
R28 VPB.t2 VPB.t15 248.598
R29 VPB.t17 VPB.t6 248.598
R30 VPB.t3 VPB.t4 248.598
R31 VPB.t5 VPB.t0 248.598
R32 VPB VPB.t5 142.056
R33 SCE.n1 SCE.t2 321.771
R34 SCE.n2 SCE.t1 266.283
R35 SCE.n0 SCE.t3 240.999
R36 SCE.n2 SCE.n1 229.346
R37 SCE.n0 SCE.t0 174.833
R38 SCE SCE.n2 20.114
R39 SCE.n1 SCE.n0 8.763
R40 VPWR.n26 VPWR.t6 429.516
R41 VPWR.n6 VPWR.t11 425.042
R42 VPWR.n43 VPWR.n42 311.893
R43 VPWR.n36 VPWR.n35 307.627
R44 VPWR.n1 VPWR.n0 186.917
R45 VPWR.n17 VPWR.n16 174.594
R46 VPWR.n3 VPWR.n2 135.028
R47 VPWR.n16 VPWR.t9 113.978
R48 VPWR.n2 VPWR.t10 61.93
R49 VPWR.n35 VPWR.t2 41.554
R50 VPWR.n35 VPWR.t1 41.554
R51 VPWR.n42 VPWR.t0 41.554
R52 VPWR.n42 VPWR.t3 41.554
R53 VPWR.n16 VPWR.t4 35.46
R54 VPWR.n2 VPWR.t7 30.223
R55 VPWR.n0 VPWR.t8 26.595
R56 VPWR.n0 VPWR.t5 26.595
R57 VPWR.n18 VPWR.n17 16.564
R58 VPWR.n3 VPWR.n1 7.521
R59 VPWR.n27 VPWR.n26 6.4
R60 VPWR.n5 VPWR.n4 4.65
R61 VPWR.n7 VPWR.n6 4.65
R62 VPWR.n9 VPWR.n8 4.65
R63 VPWR.n11 VPWR.n10 4.65
R64 VPWR.n13 VPWR.n12 4.65
R65 VPWR.n15 VPWR.n14 4.65
R66 VPWR.n19 VPWR.n18 4.65
R67 VPWR.n21 VPWR.n20 4.65
R68 VPWR.n23 VPWR.n22 4.65
R69 VPWR.n25 VPWR.n24 4.65
R70 VPWR.n28 VPWR.n27 4.65
R71 VPWR.n30 VPWR.n29 4.65
R72 VPWR.n32 VPWR.n31 4.65
R73 VPWR.n34 VPWR.n33 4.65
R74 VPWR.n37 VPWR.n36 4.65
R75 VPWR.n39 VPWR.n38 4.65
R76 VPWR.n41 VPWR.n40 4.65
R77 VPWR.n44 VPWR.n43 3.932
R78 VPWR.n5 VPWR.n3 0.141
R79 VPWR.n44 VPWR.n41 0.137
R80 VPWR VPWR.n44 0.123
R81 VPWR.n7 VPWR.n5 0.119
R82 VPWR.n9 VPWR.n7 0.119
R83 VPWR.n11 VPWR.n9 0.119
R84 VPWR.n13 VPWR.n11 0.119
R85 VPWR.n15 VPWR.n13 0.119
R86 VPWR.n19 VPWR.n15 0.119
R87 VPWR.n21 VPWR.n19 0.119
R88 VPWR.n23 VPWR.n21 0.119
R89 VPWR.n25 VPWR.n23 0.119
R90 VPWR.n28 VPWR.n25 0.119
R91 VPWR.n30 VPWR.n28 0.119
R92 VPWR.n32 VPWR.n30 0.119
R93 VPWR.n34 VPWR.n32 0.119
R94 VPWR.n37 VPWR.n34 0.119
R95 VPWR.n39 VPWR.n37 0.119
R96 VPWR.n41 VPWR.n39 0.119
R97 D.n0 D.t1 321.868
R98 D.n0 D.t0 183.694
R99 D D.n0 85.503
R100 a_465_369.t0 a_465_369.t1 93.882
R101 a_930_413.n3 a_930_413.n2 400.546
R102 a_930_413.n0 a_930_413.t5 226.539
R103 a_930_413.n2 a_930_413.n1 207.742
R104 a_930_413.n0 a_930_413.t4 196.013
R105 a_930_413.n2 a_930_413.n0 92.738
R106 a_930_413.n3 a_930_413.t2 75.047
R107 a_930_413.t0 a_930_413.n3 72.702
R108 a_930_413.n1 a_930_413.t1 65
R109 a_930_413.n1 a_930_413.t3 45
R110 a_1089_183.n1 a_1089_183.t5 433.799
R111 a_1089_183.n3 a_1089_183.n2 381.512
R112 a_1089_183.n1 a_1089_183.t4 128.098
R113 a_1089_183.n2 a_1089_183.n0 125.628
R114 a_1089_183.n2 a_1089_183.n1 109.306
R115 a_1089_183.n3 a_1089_183.t0 89.119
R116 a_1089_183.n0 a_1089_183.t3 63.333
R117 a_1089_183.t1 a_1089_183.n3 37.523
R118 a_1089_183.n0 a_1089_183.t2 36.77
R119 a_193_47.t0 a_193_47.n3 300.537
R120 a_193_47.n0 a_193_47.t2 272.659
R121 a_193_47.n1 a_193_47.t3 269.802
R122 a_193_47.n1 a_193_47.t4 205.234
R123 a_193_47.n0 a_193_47.t5 195.261
R124 a_193_47.n3 a_193_47.t1 156.671
R125 a_193_47.n2 a_193_47.n0 14.334
R126 a_193_47.n3 a_193_47.n2 7.877
R127 a_193_47.n2 a_193_47.n1 4.65
R128 a_1346_413.n3 a_1346_413.n2 400.947
R129 a_1346_413.n0 a_1346_413.t5 212.079
R130 a_1346_413.n2 a_1346_413.n0 177.675
R131 a_1346_413.n2 a_1346_413.n1 151.491
R132 a_1346_413.n0 a_1346_413.t4 139.779
R133 a_1346_413.n1 a_1346_413.t3 73.333
R134 a_1346_413.n3 a_1346_413.t2 63.321
R135 a_1346_413.t1 a_1346_413.n3 63.321
R136 a_1346_413.n1 a_1346_413.t0 48.333
R137 a_1430_413.t0 a_1430_413.t1 204.035
R138 a_1517_315.n3 a_1517_315.t3 383.498
R139 a_1517_315.n0 a_1517_315.t7 256.987
R140 a_1517_315.n1 a_1517_315.t4 212.079
R141 a_1517_315.t0 a_1517_315.n4 178.49
R142 a_1517_315.n0 a_1517_315.t5 163.801
R143 a_1517_315.n1 a_1517_315.t2 139.779
R144 a_1517_315.n3 a_1517_315.t6 139.285
R145 a_1517_315.n1 a_1517_315.n0 129.263
R146 a_1517_315.n2 a_1517_315.t1 104.195
R147 a_1517_315.n4 a_1517_315.n3 102.569
R148 a_1517_315.n2 a_1517_315.n1 97.721
R149 a_1517_315.n4 a_1517_315.n2 19.236
R150 VGND.n25 VGND.t2 163.962
R151 VGND.n6 VGND.t6 146.638
R152 VGND.n2 VGND.n1 126.005
R153 VGND.n41 VGND.n40 107.239
R154 VGND.n17 VGND.n16 107.029
R155 VGND.n34 VGND.n33 106.463
R156 VGND.n16 VGND.t9 87.142
R157 VGND.n3 VGND.n0 68.028
R158 VGND.n16 VGND.t3 66.294
R159 VGND.n33 VGND.t1 61.428
R160 VGND.n0 VGND.t7 57.796
R161 VGND.n33 VGND.t4 41.428
R162 VGND.n40 VGND.t0 38.571
R163 VGND.n40 VGND.t11 38.571
R164 VGND.n1 VGND.t8 24.923
R165 VGND.n1 VGND.t5 24.923
R166 VGND.n0 VGND.t10 24.765
R167 VGND.n3 VGND.n2 7.521
R168 VGND.n5 VGND.n4 4.65
R169 VGND.n7 VGND.n6 4.65
R170 VGND.n9 VGND.n8 4.65
R171 VGND.n11 VGND.n10 4.65
R172 VGND.n13 VGND.n12 4.65
R173 VGND.n15 VGND.n14 4.65
R174 VGND.n18 VGND.n17 4.65
R175 VGND.n20 VGND.n19 4.65
R176 VGND.n22 VGND.n21 4.65
R177 VGND.n24 VGND.n23 4.65
R178 VGND.n26 VGND.n25 4.65
R179 VGND.n28 VGND.n27 4.65
R180 VGND.n30 VGND.n29 4.65
R181 VGND.n32 VGND.n31 4.65
R182 VGND.n35 VGND.n34 4.65
R183 VGND.n37 VGND.n36 4.65
R184 VGND.n39 VGND.n38 4.65
R185 VGND.n42 VGND.n41 3.932
R186 VGND.n5 VGND.n3 0.141
R187 VGND.n42 VGND.n39 0.137
R188 VGND VGND.n42 0.123
R189 VGND.n7 VGND.n5 0.119
R190 VGND.n9 VGND.n7 0.119
R191 VGND.n11 VGND.n9 0.119
R192 VGND.n13 VGND.n11 0.119
R193 VGND.n15 VGND.n13 0.119
R194 VGND.n18 VGND.n15 0.119
R195 VGND.n20 VGND.n18 0.119
R196 VGND.n22 VGND.n20 0.119
R197 VGND.n24 VGND.n22 0.119
R198 VGND.n26 VGND.n24 0.119
R199 VGND.n28 VGND.n26 0.119
R200 VGND.n30 VGND.n28 0.119
R201 VGND.n32 VGND.n30 0.119
R202 VGND.n35 VGND.n32 0.119
R203 VGND.n37 VGND.n35 0.119
R204 VGND.n39 VGND.n37 0.119
R205 Q.n0 Q.t0 412.546
R206 Q.n0 Q.t1 83.01
R207 Q Q.n0 5.417
R208 VNB.t5 VNB.t2 6715.84
R209 VNB.t0 VNB.t3 6082.35
R210 VNB.t13 VNB.t11 5321.88
R211 VNB.t14 VNB.t12 4545.05
R212 VNB VNB.t17 4270.59
R213 VNB.t15 VNB.t7 4003.85
R214 VNB.t2 VNB.t9 3406.45
R215 VNB.t8 VNB.t1 3332.35
R216 VNB.t3 VNB.t10 3300
R217 VNB.t6 VNB.t4 3105.88
R218 VNB.t1 VNB.t13 3073.53
R219 VNB.t9 VNB.t15 3062.58
R220 VNB.t17 VNB.t0 2717.65
R221 VNB.t10 VNB.t6 2523.53
R222 VNB.t4 VNB.t5 2458.82
R223 VNB.t7 VNB.t8 2363.68
R224 VNB.t12 VNB.t16 2345.05
R225 VNB.t11 VNB.t14 2030.77
R226 a_1948_47.t0 a_1948_47.n1 244.476
R227 a_1948_47.n0 a_1948_47.t3 239.038
R228 a_1948_47.n0 a_1948_47.t2 166.738
R229 a_1948_47.n1 a_1948_47.t1 166.489
R230 a_1948_47.n1 a_1948_47.n0 98.109
R231 Q_N Q_N.t0 233.568
R232 Q_N Q_N.t1 165.324
R233 CLK.n0 CLK.t0 292.947
R234 CLK.n0 CLK.t1 209.401
R235 CLK CLK.n0 78.067
R236 a_27_47.n0 a_27_47.t3 510.426
R237 a_27_47.n1 a_27_47.t5 448.258
R238 a_27_47.n3 a_27_47.t6 263.405
R239 a_27_47.n1 a_27_47.t2 254.388
R240 a_27_47.t0 a_27_47.n5 244.156
R241 a_27_47.n3 a_27_47.t4 228.059
R242 a_27_47.n4 a_27_47.t1 198.368
R243 a_27_47.n0 a_27_47.t7 137.901
R244 a_27_47.n2 a_27_47.n1 112.811
R245 a_27_47.n4 a_27_47.n3 76
R246 a_27_47.n5 a_27_47.n4 35.339
R247 a_27_47.n2 a_27_47.n0 10.451
R248 a_27_47.n5 a_27_47.n2 8.568
R249 a_657_47.t0 a_657_47.t1 65.714
R250 SCD.n0 SCD.t1 268.848
R251 SCD.n0 SCD.t0 236.714
R252 SCD SCD.n0 82.666
R253 a_483_47.t0 a_483_47.t1 68.571
R254 a_1027_47.t1 a_1027_47.t0 98.059
R255 a_1475_47.t1 a_1475_47.t0 93.059
R256 a_1023_413.t0 a_1023_413.t1 154.785
C0 VPB VPWR 0.22fF
C1 VPWR Q 0.15fF
C2 VPWR Q_N 0.11fF
C3 VGND Q 0.11fF
C4 VGND Q_N 0.11fF
C5 VPWR VGND 0.14fF
C6 SCE VGND 0.15fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__sdfxbp_2.ext - technology: sky130A

.subckt sky130_fd_sc_hd__sdfxbp_2 VGND VPWR SCD D Q_N SCE CLK Q VNB VPB
X0 VPWR.t8 a_1525_315.t2 Q.t1 VPB.t11 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_938_413.t2 a_27_47.t2 a_560_369.t4 VNB.t14 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X2 a_466_369.t1 SCE.t0 VPWR.t4 VPB.t7 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X3 Q.t3 a_1525_315.t3 VGND.t5 VNB.t9 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 VPWR.t3 SCD.t0 a_644_369.t0 VPB.t6 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X5 Q.t0 a_1525_315.t4 VPWR.t7 VPB.t10 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 VPWR.t2 SCE.t1 a_299_47.t0 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X7 VPWR.t5 a_1525_315.t5 a_1438_413.t1 VPB.t9 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 a_1354_413.t1 a_193_47.t2 a_1097_183.t0 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X9 VGND.t6 a_1525_315.t6 a_1483_47.t0 VNB.t8 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10 VPWR.t1 a_1097_183.t4 a_1031_413.t0 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11 VPWR.t9 CLK.t0 a_27_47.t1 VPB.t12 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X12 VPWR.t12 a_2049_47.t2 Q_N.t1 VPB.t17 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13 a_487_47.t0 a_299_47.t2 VGND.t12 VNB.t18 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14 Q_N.t0 a_2049_47.t3 VPWR.t13 VPB.t18 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 a_193_47.t1 a_27_47.t3 VGND.t8 VNB.t13 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16 a_1031_413.t1 a_27_47.t4 a_938_413.t3 VPB.t14 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17 VGND.t0 a_1354_413.t4 a_1525_315.t0 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X18 VGND.t7 a_1525_315.t7 a_2049_47.t1 VNB.t7 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19 a_1097_183.t2 a_938_413.t4 VPWR.t10 VPB.t13 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X20 a_1438_413.t0 a_193_47.t3 a_1354_413.t0 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21 VPWR.t0 a_1354_413.t5 a_1525_315.t1 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X22 a_1354_413.t2 a_27_47.t5 a_1097_183.t1 VPB.t15 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23 VGND.t9 a_2049_47.t4 Q_N.t3 VNB.t15 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X24 VGND.t2 SCE.t2 a_299_47.t1 VNB.t10 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X25 a_644_369.t1 a_299_47.t3 a_560_369.t5 VPB.t19 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X26 a_661_47.t1 SCE.t3 a_560_369.t3 VNB.t11 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X27 VGND.t3 SCD.t1 a_661_47.t0 VNB.t5 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X28 VGND.t11 a_1097_183.t5 a_1035_47.t1 VNB.t17 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X29 a_560_369.t1 D.t0 a_466_369.t0 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X30 VPWR.t6 a_1525_315.t8 a_2049_47.t0 VPB.t8 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X31 a_560_369.t0 D.t1 a_487_47.t1 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X32 a_1483_47.t1 a_27_47.t6 a_1354_413.t3 VNB.t12 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X33 Q_N.t2 a_2049_47.t5 VGND.t10 VNB.t16 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X34 a_193_47.t0 a_27_47.t7 VPWR.t11 VPB.t16 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X35 a_1035_47.t0 a_193_47.t4 a_938_413.t0 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X36 VGND.t4 a_1525_315.t9 Q.t2 VNB.t6 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X37 a_938_413.t1 a_193_47.t5 a_560_369.t2 VPB.t5 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X38 VGND.t1 CLK.t1 a_27_47.t0 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X39 a_1097_183.t3 a_938_413.t5 VGND.t13 VNB.t19 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
R0 a_1525_315.n4 a_1525_315.t6 383.498
R1 a_1525_315.n0 a_1525_315.t8 256.987
R2 a_1525_315.n1 a_1525_315.t2 212.079
R3 a_1525_315.n2 a_1525_315.t4 212.079
R4 a_1525_315.n0 a_1525_315.t7 163.801
R5 a_1525_315.n1 a_1525_315.t9 139.779
R6 a_1525_315.n2 a_1525_315.t3 139.779
R7 a_1525_315.n4 a_1525_315.t5 139.285
R8 a_1525_315.n1 a_1525_315.n0 130.724
R9 a_1525_315.t1 a_1525_315.n5 127.12
R10 a_1525_315.n3 a_1525_315.t0 103.537
R11 a_1525_315.n5 a_1525_315.n4 102.375
R12 a_1525_315.n3 a_1525_315.n2 100.642
R13 a_1525_315.n2 a_1525_315.n1 61.345
R14 a_1525_315.n5 a_1525_315.n3 20.012
R15 Q.n1 Q.n0 226.502
R16 Q Q.n2 95.021
R17 Q.n0 Q.t1 26.595
R18 Q.n0 Q.t0 26.595
R19 Q.n2 Q.t2 24.923
R20 Q.n2 Q.t3 24.923
R21 Q Q.n1 10.666
R22 VPWR.n35 VPWR.t3 429.516
R23 VPWR.n15 VPWR.t5 425.042
R24 VPWR.n52 VPWR.n51 311.893
R25 VPWR.n45 VPWR.n44 307.627
R26 VPWR.n5 VPWR.t8 280.058
R27 VPWR.n11 VPWR.n10 190.72
R28 VPWR.n24 VPWR.n23 174.594
R29 VPWR.n2 VPWR.t12 165.56
R30 VPWR.n1 VPWR.n0 131.24
R31 VPWR.n23 VPWR.t1 113.978
R32 VPWR.n0 VPWR.t6 61.93
R33 VPWR.n44 VPWR.t4 41.554
R34 VPWR.n44 VPWR.t2 41.554
R35 VPWR.n51 VPWR.t11 41.554
R36 VPWR.n51 VPWR.t9 41.554
R37 VPWR.n23 VPWR.t10 35.46
R38 VPWR.n0 VPWR.t13 30.223
R39 VPWR.n10 VPWR.t7 28.565
R40 VPWR.n10 VPWR.t0 28.565
R41 VPWR.n25 VPWR.n24 15.058
R42 VPWR.n36 VPWR.n35 4.894
R43 VPWR.n4 VPWR.n3 4.65
R44 VPWR.n7 VPWR.n6 4.65
R45 VPWR.n9 VPWR.n8 4.65
R46 VPWR.n12 VPWR.n11 4.65
R47 VPWR.n14 VPWR.n13 4.65
R48 VPWR.n16 VPWR.n15 4.65
R49 VPWR.n18 VPWR.n17 4.65
R50 VPWR.n20 VPWR.n19 4.65
R51 VPWR.n22 VPWR.n21 4.65
R52 VPWR.n26 VPWR.n25 4.65
R53 VPWR.n28 VPWR.n27 4.65
R54 VPWR.n30 VPWR.n29 4.65
R55 VPWR.n32 VPWR.n31 4.65
R56 VPWR.n34 VPWR.n33 4.65
R57 VPWR.n37 VPWR.n36 4.65
R58 VPWR.n39 VPWR.n38 4.65
R59 VPWR.n41 VPWR.n40 4.65
R60 VPWR.n43 VPWR.n42 4.65
R61 VPWR.n46 VPWR.n45 4.65
R62 VPWR.n48 VPWR.n47 4.65
R63 VPWR.n50 VPWR.n49 4.65
R64 VPWR.n53 VPWR.n52 3.941
R65 VPWR.n2 VPWR.n1 3.72
R66 VPWR.n6 VPWR.n5 3.011
R67 VPWR.n4 VPWR.n2 0.271
R68 VPWR.n53 VPWR.n50 0.137
R69 VPWR VPWR.n53 0.123
R70 VPWR.n7 VPWR.n4 0.119
R71 VPWR.n9 VPWR.n7 0.119
R72 VPWR.n12 VPWR.n9 0.119
R73 VPWR.n14 VPWR.n12 0.119
R74 VPWR.n16 VPWR.n14 0.119
R75 VPWR.n18 VPWR.n16 0.119
R76 VPWR.n20 VPWR.n18 0.119
R77 VPWR.n22 VPWR.n20 0.119
R78 VPWR.n26 VPWR.n22 0.119
R79 VPWR.n28 VPWR.n26 0.119
R80 VPWR.n30 VPWR.n28 0.119
R81 VPWR.n32 VPWR.n30 0.119
R82 VPWR.n34 VPWR.n32 0.119
R83 VPWR.n37 VPWR.n34 0.119
R84 VPWR.n39 VPWR.n37 0.119
R85 VPWR.n41 VPWR.n39 0.119
R86 VPWR.n43 VPWR.n41 0.119
R87 VPWR.n46 VPWR.n43 0.119
R88 VPWR.n48 VPWR.n46 0.119
R89 VPWR.n50 VPWR.n48 0.119
R90 VPB.t9 VPB.t0 633.333
R91 VPB.t6 VPB.t5 594.859
R92 VPB.t11 VPB.t8 562.305
R93 VPB.t16 VPB.t3 556.386
R94 VPB.t1 VPB.t13 390.654
R95 VPB.t2 VPB.t9 346.261
R96 VPB.t8 VPB.t18 287.071
R97 VPB.t14 VPB.t1 284.112
R98 VPB.t13 VPB.t15 281.152
R99 VPB.t7 VPB.t4 278.193
R100 VPB.t5 VPB.t14 275.233
R101 VPB.t19 VPB.t6 275.233
R102 VPB.t0 VPB.t10 260.436
R103 VPB.t18 VPB.t17 248.598
R104 VPB.t10 VPB.t11 248.598
R105 VPB.t15 VPB.t2 248.598
R106 VPB.t4 VPB.t19 248.598
R107 VPB.t3 VPB.t7 248.598
R108 VPB.t12 VPB.t16 248.598
R109 VPB VPB.t12 145.015
R110 a_27_47.n0 a_27_47.t2 510.426
R111 a_27_47.n1 a_27_47.t6 448.258
R112 a_27_47.n3 a_27_47.t7 263.171
R113 a_27_47.n1 a_27_47.t5 254.388
R114 a_27_47.t1 a_27_47.n5 243.779
R115 a_27_47.n3 a_27_47.t3 227.825
R116 a_27_47.n4 a_27_47.t0 198.368
R117 a_27_47.n0 a_27_47.t4 137.901
R118 a_27_47.n2 a_27_47.n1 112.819
R119 a_27_47.n4 a_27_47.n3 76
R120 a_27_47.n5 a_27_47.n4 35.339
R121 a_27_47.n2 a_27_47.n0 10.451
R122 a_27_47.n5 a_27_47.n2 8.604
R123 a_560_369.n3 a_560_369.n2 413.345
R124 a_560_369.n2 a_560_369.t2 373.036
R125 a_560_369.n1 a_560_369.n0 207.322
R126 a_560_369.n1 a_560_369.t4 163.742
R127 a_560_369.n2 a_560_369.n1 72.282
R128 a_560_369.n0 a_560_369.t0 54.285
R129 a_560_369.n3 a_560_369.t5 41.554
R130 a_560_369.t1 a_560_369.n3 41.554
R131 a_560_369.n0 a_560_369.t3 40
R132 a_938_413.n3 a_938_413.n2 400.546
R133 a_938_413.n0 a_938_413.t5 226.539
R134 a_938_413.n2 a_938_413.n1 207.742
R135 a_938_413.n0 a_938_413.t4 196.013
R136 a_938_413.n2 a_938_413.n0 92.738
R137 a_938_413.t1 a_938_413.n3 75.047
R138 a_938_413.n3 a_938_413.t3 72.702
R139 a_938_413.n1 a_938_413.t2 65
R140 a_938_413.n1 a_938_413.t0 45
R141 VNB.t5 VNB.t14 6845.25
R142 VNB.t13 VNB.t10 6211.76
R143 VNB.t8 VNB.t0 5418.94
R144 VNB.t6 VNB.t7 4593.41
R145 VNB VNB.t1 4270.59
R146 VNB.t17 VNB.t19 4003.85
R147 VNB.t14 VNB.t3 3406.45
R148 VNB.t2 VNB.t12 3332.35
R149 VNB.t10 VNB.t18 3300
R150 VNB.t4 VNB.t11 3105.88
R151 VNB.t12 VNB.t8 3073.53
R152 VNB.t3 VNB.t17 3062.58
R153 VNB.t1 VNB.t13 2717.65
R154 VNB.t18 VNB.t4 2523.53
R155 VNB.t11 VNB.t5 2458.82
R156 VNB.t19 VNB.t2 2363.68
R157 VNB.t7 VNB.t16 2345.05
R158 VNB.t0 VNB.t9 2127.47
R159 VNB.t16 VNB.t15 2030.77
R160 VNB.t9 VNB.t6 2030.77
R161 SCE.n1 SCE.t2 321.771
R162 SCE.n2 SCE.t3 266.283
R163 SCE.n0 SCE.t0 236.179
R164 SCE.n2 SCE.n1 177.27
R165 SCE.n0 SCE.t1 174.833
R166 SCE SCE.n2 20.114
R167 SCE.n1 SCE.n0 8.763
R168 a_466_369.t0 a_466_369.t1 98.5
R169 VGND.n33 VGND.t3 162.682
R170 VGND.n5 VGND.t4 148.486
R171 VGND.n14 VGND.t6 146.638
R172 VGND.n10 VGND.n9 128.205
R173 VGND.n2 VGND.t9 120.012
R174 VGND.n49 VGND.n48 107.239
R175 VGND.n25 VGND.n24 107.029
R176 VGND.n42 VGND.n41 106.463
R177 VGND.n24 VGND.t11 87.142
R178 VGND.n24 VGND.t13 66.294
R179 VGND.n1 VGND.n0 64.275
R180 VGND.n41 VGND.t2 61.428
R181 VGND.n0 VGND.t7 57.796
R182 VGND.n41 VGND.t12 41.428
R183 VGND.n48 VGND.t8 38.571
R184 VGND.n48 VGND.t1 38.571
R185 VGND.n9 VGND.t5 26.769
R186 VGND.n9 VGND.t0 26.769
R187 VGND.n0 VGND.t10 24.765
R188 VGND.n4 VGND.n3 4.65
R189 VGND.n6 VGND.n5 4.65
R190 VGND.n8 VGND.n7 4.65
R191 VGND.n11 VGND.n10 4.65
R192 VGND.n13 VGND.n12 4.65
R193 VGND.n15 VGND.n14 4.65
R194 VGND.n17 VGND.n16 4.65
R195 VGND.n19 VGND.n18 4.65
R196 VGND.n21 VGND.n20 4.65
R197 VGND.n23 VGND.n22 4.65
R198 VGND.n26 VGND.n25 4.65
R199 VGND.n28 VGND.n27 4.65
R200 VGND.n30 VGND.n29 4.65
R201 VGND.n32 VGND.n31 4.65
R202 VGND.n34 VGND.n33 4.65
R203 VGND.n36 VGND.n35 4.65
R204 VGND.n38 VGND.n37 4.65
R205 VGND.n40 VGND.n39 4.65
R206 VGND.n43 VGND.n42 4.65
R207 VGND.n45 VGND.n44 4.65
R208 VGND.n47 VGND.n46 4.65
R209 VGND.n50 VGND.n49 3.932
R210 VGND.n2 VGND.n1 3.72
R211 VGND.n4 VGND.n2 0.271
R212 VGND.n50 VGND.n47 0.137
R213 VGND VGND.n50 0.123
R214 VGND.n6 VGND.n4 0.119
R215 VGND.n8 VGND.n6 0.119
R216 VGND.n11 VGND.n8 0.119
R217 VGND.n13 VGND.n11 0.119
R218 VGND.n15 VGND.n13 0.119
R219 VGND.n17 VGND.n15 0.119
R220 VGND.n19 VGND.n17 0.119
R221 VGND.n21 VGND.n19 0.119
R222 VGND.n23 VGND.n21 0.119
R223 VGND.n26 VGND.n23 0.119
R224 VGND.n28 VGND.n26 0.119
R225 VGND.n30 VGND.n28 0.119
R226 VGND.n32 VGND.n30 0.119
R227 VGND.n34 VGND.n32 0.119
R228 VGND.n36 VGND.n34 0.119
R229 VGND.n38 VGND.n36 0.119
R230 VGND.n40 VGND.n38 0.119
R231 VGND.n43 VGND.n40 0.119
R232 VGND.n45 VGND.n43 0.119
R233 VGND.n47 VGND.n45 0.119
R234 SCD.n0 SCD.t1 268.848
R235 SCD.n0 SCD.t0 236.714
R236 SCD SCD.n0 82.4
R237 a_644_369.t0 a_644_369.t1 96.96
R238 a_299_47.t0 a_299_47.n1 343.828
R239 a_299_47.n0 a_299_47.t3 340.853
R240 a_299_47.n0 a_299_47.t2 306.024
R241 a_299_47.n1 a_299_47.t1 251.534
R242 a_299_47.n1 a_299_47.n0 29.469
R243 a_1438_413.t0 a_1438_413.t1 204.035
R244 a_193_47.t0 a_193_47.n3 278.596
R245 a_193_47.n0 a_193_47.t3 272.659
R246 a_193_47.n1 a_193_47.t5 268.251
R247 a_193_47.n1 a_193_47.t4 206.786
R248 a_193_47.n0 a_193_47.t2 195.261
R249 a_193_47.n3 a_193_47.t1 150.159
R250 a_193_47.n2 a_193_47.n0 13.802
R251 a_193_47.n3 a_193_47.n2 7.846
R252 a_193_47.n2 a_193_47.n1 4.65
R253 a_1097_183.n1 a_1097_183.t4 433.799
R254 a_1097_183.n3 a_1097_183.n2 381.512
R255 a_1097_183.n1 a_1097_183.t5 128.098
R256 a_1097_183.n2 a_1097_183.n0 125.628
R257 a_1097_183.n2 a_1097_183.n1 109.306
R258 a_1097_183.n3 a_1097_183.t1 89.119
R259 a_1097_183.n0 a_1097_183.t0 63.333
R260 a_1097_183.t2 a_1097_183.n3 37.523
R261 a_1097_183.n0 a_1097_183.t3 36.77
R262 a_1354_413.n3 a_1354_413.n2 400.947
R263 a_1354_413.n0 a_1354_413.t5 212.079
R264 a_1354_413.n2 a_1354_413.n0 178.257
R265 a_1354_413.n2 a_1354_413.n1 151.491
R266 a_1354_413.n0 a_1354_413.t4 139.779
R267 a_1354_413.n1 a_1354_413.t1 73.333
R268 a_1354_413.t0 a_1354_413.n3 63.321
R269 a_1354_413.n3 a_1354_413.t2 63.321
R270 a_1354_413.n1 a_1354_413.t3 48.333
R271 a_1483_47.t0 a_1483_47.t1 93.059
R272 a_1031_413.t0 a_1031_413.t1 154.785
R273 CLK.n0 CLK.t0 294.554
R274 CLK.n0 CLK.t1 209.401
R275 CLK CLK.n0 77.87
R276 a_2049_47.t0 a_2049_47.n2 240.007
R277 a_2049_47.n0 a_2049_47.t2 212.079
R278 a_2049_47.n1 a_2049_47.t3 212.079
R279 a_2049_47.n2 a_2049_47.t1 157.454
R280 a_2049_47.n0 a_2049_47.t4 139.779
R281 a_2049_47.n1 a_2049_47.t5 139.779
R282 a_2049_47.n2 a_2049_47.n1 112.075
R283 a_2049_47.n1 a_2049_47.n0 61.345
R284 Q_N Q_N.n1 169.677
R285 Q_N Q_N.n0 141.533
R286 Q_N.n1 Q_N.t1 26.595
R287 Q_N.n1 Q_N.t0 26.595
R288 Q_N.n0 Q_N.t3 24.923
R289 Q_N.n0 Q_N.t2 24.923
R290 a_487_47.t0 a_487_47.t1 68.571
R291 a_661_47.t0 a_661_47.t1 65.714
R292 a_1035_47.t1 a_1035_47.t0 98.059
R293 D.n0 D.t1 321.868
R294 D.n0 D.t0 183.694
R295 D D.n0 85.115
C0 VPWR VGND 0.19fF
C1 SCE VGND 0.15fF
C2 VPB VPWR 0.25fF
C3 VPWR Q 0.24fF
C4 VPWR Q_N 0.25fF
C5 VGND Q 0.17fF
C6 VGND Q_N 0.21fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__sdfxtp_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__sdfxtp_1 VPWR VGND Q CLK SCE D SCD VNB VPB
X0 a_640_369.t0 a_299_47.t2 a_556_369.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1 a_933_413.t0 a_193_47.t2 a_556_369.t5 VPB.t8 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 a_556_369.t3 D.t0 a_467_369.t1 VPB.t7 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X3 a_1030_47.t0 a_193_47.t3 a_933_413.t1 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X4 a_1092_183.t2 a_933_413.t4 VGND.t9 VNB.t15 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X5 VPWR.t0 a_1349_413.t4 a_1520_315.t1 VPB.t14 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 VPWR.t2 SCE.t0 a_299_47.t0 VPB.t5 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X7 Q.t1 a_1520_315.t2 VPWR.t4 VPB.t12 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 VPWR.t6 CLK.t0 a_27_47.t1 VPB.t11 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X9 a_467_369.t0 SCE.t1 VPWR.t3 VPB.t6 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X10 a_1026_413.t0 a_27_47.t2 a_933_413.t2 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11 a_657_47.t1 SCE.t2 a_556_369.t2 VNB.t7 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12 VPWR.t5 a_1520_315.t3 a_1433_413.t1 VPB.t13 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13 a_933_413.t3 a_27_47.t3 a_556_369.t1 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X14 Q.t0 a_1520_315.t4 VGND.t4 VNB.t10 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X15 VPWR.t8 a_1092_183.t4 a_1026_413.t1 VPB.t10 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16 VGND.t1 a_1092_183.t5 a_1030_47.t1 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17 VGND.t5 a_1520_315.t5 a_1478_47.t1 VNB.t11 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18 a_193_47.t1 a_27_47.t4 VGND.t2 VNB.t5 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19 a_483_47.t0 a_299_47.t3 VGND.t0 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20 a_1478_47.t0 a_27_47.t5 a_1349_413.t3 VNB.t6 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X21 VPWR.t7 SCD.t0 a_640_369.t1 VPB.t15 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X22 a_1433_413.t0 a_193_47.t4 a_1349_413.t0 VPB.t9 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23 VGND.t8 SCE.t3 a_299_47.t1 VNB.t14 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24 a_1092_183.t3 a_933_413.t5 VPWR.t9 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X25 a_1349_413.t2 a_27_47.t6 a_1092_183.t1 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X26 VGND.t6 a_1349_413.t5 a_1520_315.t0 VNB.t12 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X27 VGND.t3 SCD.t1 a_657_47.t0 VNB.t8 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X28 a_1349_413.t1 a_193_47.t5 a_1092_183.t0 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X29 a_193_47.t0 a_27_47.t7 VPWR.t1 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X30 VGND.t7 CLK.t1 a_27_47.t0 VNB.t13 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X31 a_556_369.t4 D.t1 a_483_47.t1 VNB.t9 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
R0 a_299_47.n0 a_299_47.t2 357.967
R1 a_299_47.t0 a_299_47.n1 343.322
R2 a_299_47.n0 a_299_47.t3 304.749
R3 a_299_47.n1 a_299_47.t1 252.518
R4 a_299_47.n1 a_299_47.n0 29.172
R5 a_556_369.n3 a_556_369.n2 412.969
R6 a_556_369.n2 a_556_369.t5 393.398
R7 a_556_369.n1 a_556_369.n0 208.452
R8 a_556_369.n1 a_556_369.t1 157.571
R9 a_556_369.n2 a_556_369.n1 70.776
R10 a_556_369.n0 a_556_369.t4 54.285
R11 a_556_369.t0 a_556_369.n3 41.554
R12 a_556_369.n3 a_556_369.t3 41.554
R13 a_556_369.n0 a_556_369.t2 40
R14 a_640_369.t0 a_640_369.t1 98.5
R15 VPB.t13 VPB.t14 624.454
R16 VPB.t15 VPB.t8 588.94
R17 VPB.t4 VPB.t5 556.386
R18 VPB.t10 VPB.t1 390.654
R19 VPB.t9 VPB.t13 346.261
R20 VPB.t2 VPB.t10 284.112
R21 VPB.t1 VPB.t3 281.152
R22 VPB.t0 VPB.t15 278.193
R23 VPB.t8 VPB.t2 275.233
R24 VPB.t14 VPB.t12 269.314
R25 VPB.t6 VPB.t7 263.395
R26 VPB.t5 VPB.t6 251.557
R27 VPB.t3 VPB.t9 248.598
R28 VPB.t7 VPB.t0 248.598
R29 VPB.t11 VPB.t4 248.598
R30 VPB VPB.t11 145.015
R31 a_193_47.t0 a_193_47.n3 283.442
R32 a_193_47.n0 a_193_47.t4 272.659
R33 a_193_47.n1 a_193_47.t2 271.388
R34 a_193_47.n1 a_193_47.t3 207.926
R35 a_193_47.n0 a_193_47.t5 195.261
R36 a_193_47.n3 a_193_47.t1 151.503
R37 a_193_47.n2 a_193_47.n0 13.211
R38 a_193_47.n3 a_193_47.n2 7.855
R39 a_193_47.n2 a_193_47.n1 4.65
R40 a_933_413.n3 a_933_413.n2 400.546
R41 a_933_413.n0 a_933_413.t4 226.539
R42 a_933_413.n2 a_933_413.n1 207.742
R43 a_933_413.n0 a_933_413.t5 196.013
R44 a_933_413.n2 a_933_413.n0 92.738
R45 a_933_413.t0 a_933_413.n3 75.047
R46 a_933_413.n3 a_933_413.t2 72.702
R47 a_933_413.n1 a_933_413.t3 65
R48 a_933_413.n1 a_933_413.t1 45
R49 D.n0 D.t1 321.868
R50 D.n0 D.t0 183.694
R51 D D.n0 83.757
R52 a_467_369.t0 a_467_369.t1 90.804
R53 a_1030_47.t1 a_1030_47.t0 98.059
R54 VNB.t8 VNB.t4 6809.77
R55 VNB.t5 VNB.t14 6211.76
R56 VNB.t11 VNB.t12 5321.88
R57 VNB VNB.t13 4270.59
R58 VNB.t3 VNB.t15 4003.85
R59 VNB.t4 VNB.t2 3406.45
R60 VNB.t1 VNB.t6 3332.35
R61 VNB.t14 VNB.t0 3170.59
R62 VNB.t9 VNB.t7 3105.88
R63 VNB.t6 VNB.t11 3073.53
R64 VNB.t2 VNB.t3 3062.58
R65 VNB.t13 VNB.t5 2717.65
R66 VNB.t0 VNB.t9 2523.53
R67 VNB.t7 VNB.t8 2458.82
R68 VNB.t15 VNB.t1 2363.68
R69 VNB.t12 VNB.t10 2200
R70 VGND.n20 VGND.t3 169.677
R71 VGND.n1 VGND.t5 146.638
R72 VGND.n2 VGND.n0 130.491
R73 VGND.n36 VGND.n35 107.239
R74 VGND.n12 VGND.n11 107.029
R75 VGND.n29 VGND.n28 105.856
R76 VGND.n11 VGND.t1 87.142
R77 VGND.n11 VGND.t9 66.294
R78 VGND.n28 VGND.t8 57.142
R79 VGND.n28 VGND.t0 40
R80 VGND.n35 VGND.t2 38.571
R81 VGND.n35 VGND.t7 38.571
R82 VGND.n0 VGND.t6 28.615
R83 VGND.n0 VGND.t4 27.692
R84 VGND.n4 VGND.n3 4.65
R85 VGND.n6 VGND.n5 4.65
R86 VGND.n8 VGND.n7 4.65
R87 VGND.n10 VGND.n9 4.65
R88 VGND.n13 VGND.n12 4.65
R89 VGND.n15 VGND.n14 4.65
R90 VGND.n17 VGND.n16 4.65
R91 VGND.n19 VGND.n18 4.65
R92 VGND.n21 VGND.n20 4.65
R93 VGND.n23 VGND.n22 4.65
R94 VGND.n25 VGND.n24 4.65
R95 VGND.n27 VGND.n26 4.65
R96 VGND.n30 VGND.n29 4.65
R97 VGND.n32 VGND.n31 4.65
R98 VGND.n34 VGND.n33 4.65
R99 VGND.n2 VGND.n1 4.048
R100 VGND.n37 VGND.n36 3.932
R101 VGND.n4 VGND.n2 0.194
R102 VGND.n37 VGND.n34 0.137
R103 VGND VGND.n37 0.123
R104 VGND.n6 VGND.n4 0.119
R105 VGND.n8 VGND.n6 0.119
R106 VGND.n10 VGND.n8 0.119
R107 VGND.n13 VGND.n10 0.119
R108 VGND.n15 VGND.n13 0.119
R109 VGND.n17 VGND.n15 0.119
R110 VGND.n19 VGND.n17 0.119
R111 VGND.n21 VGND.n19 0.119
R112 VGND.n23 VGND.n21 0.119
R113 VGND.n25 VGND.n23 0.119
R114 VGND.n27 VGND.n25 0.119
R115 VGND.n30 VGND.n27 0.119
R116 VGND.n32 VGND.n30 0.119
R117 VGND.n34 VGND.n32 0.119
R118 a_1092_183.n1 a_1092_183.t4 433.799
R119 a_1092_183.n3 a_1092_183.n2 381.512
R120 a_1092_183.n1 a_1092_183.t5 128.098
R121 a_1092_183.n2 a_1092_183.n0 125.628
R122 a_1092_183.n2 a_1092_183.n1 109.306
R123 a_1092_183.n3 a_1092_183.t1 89.119
R124 a_1092_183.n0 a_1092_183.t0 63.333
R125 a_1092_183.t3 a_1092_183.n3 37.523
R126 a_1092_183.n0 a_1092_183.t2 36.77
R127 a_1349_413.n3 a_1349_413.n2 400.947
R128 a_1349_413.n0 a_1349_413.t4 212.079
R129 a_1349_413.n2 a_1349_413.n0 173.92
R130 a_1349_413.n2 a_1349_413.n1 151.491
R131 a_1349_413.n0 a_1349_413.t5 139.779
R132 a_1349_413.n1 a_1349_413.t1 73.333
R133 a_1349_413.t0 a_1349_413.n3 63.321
R134 a_1349_413.n3 a_1349_413.t2 63.321
R135 a_1349_413.n1 a_1349_413.t3 48.333
R136 a_1520_315.t1 a_1520_315.n4 523.596
R137 a_1520_315.n3 a_1520_315.t5 383.498
R138 a_1520_315.n0 a_1520_315.t2 236.932
R139 a_1520_315.n0 a_1520_315.t4 164.632
R140 a_1520_315.n3 a_1520_315.t3 139.285
R141 a_1520_315.n1 a_1520_315.t0 104.842
R142 a_1520_315.n4 a_1520_315.n3 101.793
R143 a_1520_315.n1 a_1520_315.n0 96.557
R144 a_1520_315.n2 a_1520_315.n1 20.762
R145 a_1520_315.n4 a_1520_315.n2 1.939
R146 VPWR.n21 VPWR.t7 438.488
R147 VPWR.n1 VPWR.t5 425.042
R148 VPWR.n37 VPWR.n36 311.893
R149 VPWR.n30 VPWR.n29 307.627
R150 VPWR.n2 VPWR.n0 191.401
R151 VPWR.n10 VPWR.n9 174.594
R152 VPWR.n9 VPWR.t8 113.978
R153 VPWR.n29 VPWR.t3 43.093
R154 VPWR.n29 VPWR.t2 41.554
R155 VPWR.n36 VPWR.t1 41.554
R156 VPWR.n36 VPWR.t6 41.554
R157 VPWR.n9 VPWR.t9 35.46
R158 VPWR.n0 VPWR.t0 30.535
R159 VPWR.n0 VPWR.t4 29.55
R160 VPWR.n11 VPWR.n10 16.941
R161 VPWR.n4 VPWR.n3 4.65
R162 VPWR.n6 VPWR.n5 4.65
R163 VPWR.n8 VPWR.n7 4.65
R164 VPWR.n12 VPWR.n11 4.65
R165 VPWR.n14 VPWR.n13 4.65
R166 VPWR.n16 VPWR.n15 4.65
R167 VPWR.n18 VPWR.n17 4.65
R168 VPWR.n20 VPWR.n19 4.65
R169 VPWR.n22 VPWR.n21 4.65
R170 VPWR.n24 VPWR.n23 4.65
R171 VPWR.n26 VPWR.n25 4.65
R172 VPWR.n28 VPWR.n27 4.65
R173 VPWR.n31 VPWR.n30 4.65
R174 VPWR.n33 VPWR.n32 4.65
R175 VPWR.n35 VPWR.n34 4.65
R176 VPWR.n2 VPWR.n1 4.036
R177 VPWR.n38 VPWR.n37 3.941
R178 VPWR.n4 VPWR.n2 0.196
R179 VPWR.n38 VPWR.n35 0.137
R180 VPWR VPWR.n38 0.123
R181 VPWR.n6 VPWR.n4 0.119
R182 VPWR.n8 VPWR.n6 0.119
R183 VPWR.n12 VPWR.n8 0.119
R184 VPWR.n14 VPWR.n12 0.119
R185 VPWR.n16 VPWR.n14 0.119
R186 VPWR.n18 VPWR.n16 0.119
R187 VPWR.n20 VPWR.n18 0.119
R188 VPWR.n22 VPWR.n20 0.119
R189 VPWR.n24 VPWR.n22 0.119
R190 VPWR.n26 VPWR.n24 0.119
R191 VPWR.n28 VPWR.n26 0.119
R192 VPWR.n31 VPWR.n28 0.119
R193 VPWR.n33 VPWR.n31 0.119
R194 VPWR.n35 VPWR.n33 0.119
R195 SCE.n1 SCE.t3 319.83
R196 SCE.n2 SCE.t2 255.441
R197 SCE.n0 SCE.t1 244.212
R198 SCE.n2 SCE.n1 184.617
R199 SCE.n0 SCE.t0 175.54
R200 SCE SCE.n2 20.114
R201 SCE.n1 SCE.n0 9.329
R202 Q.n2 Q.n1 292.5
R203 Q.n3 Q.n2 146.523
R204 Q.n0 Q.t0 82.969
R205 Q.n1 Q.n0 64.987
R206 Q.n2 Q.t1 26.595
R207 Q.n3 Q 9.678
R208 Q.n1 Q 5.75
R209 Q.n0 Q 5.508
R210 Q Q.n3 2.881
R211 CLK.n0 CLK.t0 294.554
R212 CLK.n0 CLK.t1 209.401
R213 CLK CLK.n0 78.067
R214 a_27_47.n1 a_27_47.t3 501.814
R215 a_27_47.n0 a_27_47.t5 448.258
R216 a_27_47.n3 a_27_47.t7 263.171
R217 a_27_47.n0 a_27_47.t6 254.388
R218 a_27_47.t1 a_27_47.n5 243.779
R219 a_27_47.n3 a_27_47.t4 227.825
R220 a_27_47.n4 a_27_47.t0 198.368
R221 a_27_47.n1 a_27_47.t2 148.348
R222 a_27_47.n2 a_27_47.n0 112.772
R223 a_27_47.n2 a_27_47.n1 86.959
R224 a_27_47.n4 a_27_47.n3 76
R225 a_27_47.n5 a_27_47.n4 35.339
R226 a_27_47.n5 a_27_47.n2 8.622
R227 a_1026_413.t0 a_1026_413.t1 154.785
R228 a_657_47.t0 a_657_47.t1 65.714
R229 a_1433_413.t0 a_1433_413.t1 204.035
R230 a_1478_47.t1 a_1478_47.t0 93.059
R231 a_483_47.t0 a_483_47.t1 68.571
R232 SCD.n0 SCD.t1 255.149
R233 SCD.n0 SCD.t0 236.113
R234 SCD SCD.n0 82.956
C0 VGND Q 0.10fF
C1 VPWR VGND 0.10fF
C2 SCE VGND 0.15fF
C3 VPB VPWR 0.19fF
C4 VPWR Q 0.15fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__sdfxtp_2.ext - technology: sky130A

.subckt sky130_fd_sc_hd__sdfxtp_2 VGND VPWR SCD D SCE CLK Q VNB VPB
X0 VPWR.t5 SCD.t0 a_643_369.t1 VPB.t10 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1 Q.t1 a_1526_315.t2 VGND.t4 VNB.t8 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 a_939_413.t2 a_193_47.t2 a_559_369.t1 VPB.t8 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3 a_1355_413.t2 a_193_47.t3 a_1098_183.t1 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X4 VGND.t5 a_1526_315.t3 a_1484_47.t1 VNB.t7 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 VPWR.t10 SCE.t0 a_299_47.t1 VPB.t16 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X6 VPWR.t8 a_1355_413.t4 a_1526_315.t0 VPB.t14 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 VPWR.t1 a_1526_315.t4 Q.t3 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 VPWR.t4 CLK.t0 a_27_47.t1 VPB.t7 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X9 a_467_369.t1 SCE.t1 VPWR.t9 VPB.t15 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X10 VPWR.t2 a_1526_315.t5 a_1439_413.t1 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11 Q.t2 a_1526_315.t6 VPWR.t0 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 a_486_47.t0 a_299_47.t2 VGND.t0 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13 VPWR.t6 a_1098_183.t4 a_1032_413.t0 VPB.t12 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14 a_193_47.t1 a_27_47.t2 VGND.t8 VNB.t11 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15 a_1098_183.t2 a_939_413.t4 VGND.t7 VNB.t10 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X16 a_643_369.t0 a_299_47.t3 a_559_369.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X17 VGND.t9 a_1355_413.t5 a_1526_315.t1 VNB.t13 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X18 a_559_369.t2 D.t0 a_467_369.t0 VPB.t11 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X19 a_939_413.t3 a_27_47.t3 a_559_369.t3 VNB.t12 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X20 a_1032_413.t1 a_27_47.t4 a_939_413.t0 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21 VGND.t10 SCE.t2 a_299_47.t0 VNB.t14 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22 VGND.t6 a_1098_183.t5 a_1036_47.t0 VNB.t9 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23 a_1098_183.t3 a_939_413.t5 VPWR.t7 VPB.t13 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X24 a_1439_413.t0 a_193_47.t4 a_1355_413.t3 VPB.t9 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X25 a_660_47.t1 SCE.t3 a_559_369.t4 VNB.t15 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X26 VGND.t2 SCD.t1 a_660_47.t0 VNB.t5 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X27 a_1355_413.t0 a_27_47.t5 a_1098_183.t0 VPB.t5 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X28 a_1484_47.t0 a_27_47.t6 a_1355_413.t1 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X29 a_193_47.t0 a_27_47.t7 VPWR.t3 VPB.t6 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X30 a_559_369.t5 D.t1 a_486_47.t1 VNB.t16 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X31 a_1036_47.t1 a_193_47.t5 a_939_413.t1 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X32 VGND.t3 a_1526_315.t7 Q.t0 VNB.t6 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X33 VGND.t1 CLK.t1 a_27_47.t0 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
R0 SCD.n0 SCD.t1 268.848
R1 SCD.n0 SCD.t0 236.714
R2 SCD.n1 SCD.n0 76
R3 SCD.n1 SCD 6.53
R4  SCD.n1 2.351
R5 a_643_369.t0 a_643_369.t1 96.96
R6 VPWR.n25 VPWR.t5 429.516
R7 VPWR.n5 VPWR.t2 425.042
R8 VPWR.n42 VPWR.n41 311.893
R9 VPWR.n35 VPWR.n34 307.627
R10 VPWR.n1 VPWR.n0 191.982
R11 VPWR.n14 VPWR.n13 174.594
R12 VPWR.n2 VPWR.t1 170.567
R13 VPWR.n13 VPWR.t6 113.978
R14 VPWR.n34 VPWR.t9 43.093
R15 VPWR.n34 VPWR.t10 41.554
R16 VPWR.n41 VPWR.t3 41.554
R17 VPWR.n41 VPWR.t4 41.554
R18 VPWR.n13 VPWR.t7 35.46
R19 VPWR.n0 VPWR.t8 30.535
R20 VPWR.n0 VPWR.t0 29.55
R21 VPWR.n15 VPWR.n14 14.682
R22 VPWR.n26 VPWR.n25 5.27
R23 VPWR.n4 VPWR.n3 4.65
R24 VPWR.n6 VPWR.n5 4.65
R25 VPWR.n8 VPWR.n7 4.65
R26 VPWR.n10 VPWR.n9 4.65
R27 VPWR.n12 VPWR.n11 4.65
R28 VPWR.n16 VPWR.n15 4.65
R29 VPWR.n18 VPWR.n17 4.65
R30 VPWR.n20 VPWR.n19 4.65
R31 VPWR.n22 VPWR.n21 4.65
R32 VPWR.n24 VPWR.n23 4.65
R33 VPWR.n27 VPWR.n26 4.65
R34 VPWR.n29 VPWR.n28 4.65
R35 VPWR.n31 VPWR.n30 4.65
R36 VPWR.n33 VPWR.n32 4.65
R37 VPWR.n36 VPWR.n35 4.65
R38 VPWR.n38 VPWR.n37 4.65
R39 VPWR.n40 VPWR.n39 4.65
R40 VPWR.n43 VPWR.n42 3.941
R41 VPWR.n2 VPWR.n1 3.924
R42 VPWR.n4 VPWR.n2 0.233
R43 VPWR.n43 VPWR.n40 0.137
R44 VPWR VPWR.n43 0.123
R45 VPWR.n6 VPWR.n4 0.119
R46 VPWR.n8 VPWR.n6 0.119
R47 VPWR.n10 VPWR.n8 0.119
R48 VPWR.n12 VPWR.n10 0.119
R49 VPWR.n16 VPWR.n12 0.119
R50 VPWR.n18 VPWR.n16 0.119
R51 VPWR.n20 VPWR.n18 0.119
R52 VPWR.n22 VPWR.n20 0.119
R53 VPWR.n24 VPWR.n22 0.119
R54 VPWR.n27 VPWR.n24 0.119
R55 VPWR.n29 VPWR.n27 0.119
R56 VPWR.n31 VPWR.n29 0.119
R57 VPWR.n33 VPWR.n31 0.119
R58 VPWR.n36 VPWR.n33 0.119
R59 VPWR.n38 VPWR.n36 0.119
R60 VPWR.n40 VPWR.n38 0.119
R61 VPB.t3 VPB.t14 624.454
R62 VPB.t10 VPB.t8 600.778
R63 VPB.t6 VPB.t16 556.386
R64 VPB.t12 VPB.t13 390.654
R65 VPB.t9 VPB.t3 346.261
R66 VPB.t4 VPB.t12 284.112
R67 VPB.t13 VPB.t5 281.152
R68 VPB.t8 VPB.t4 275.233
R69 VPB.t0 VPB.t10 275.233
R70 VPB.t15 VPB.t11 272.274
R71 VPB.t14 VPB.t1 269.314
R72 VPB.t16 VPB.t15 251.557
R73 VPB.t1 VPB.t2 248.598
R74 VPB.t5 VPB.t9 248.598
R75 VPB.t11 VPB.t0 248.598
R76 VPB.t7 VPB.t6 248.598
R77 VPB VPB.t7 145.015
R78 a_1526_315.t0 a_1526_315.n5 523.596
R79 a_1526_315.n4 a_1526_315.t3 383.498
R80 a_1526_315.n0 a_1526_315.t4 212.079
R81 a_1526_315.n1 a_1526_315.t6 212.079
R82 a_1526_315.n0 a_1526_315.t7 139.779
R83 a_1526_315.n1 a_1526_315.t2 139.779
R84 a_1526_315.n4 a_1526_315.t5 139.285
R85 a_1526_315.n2 a_1526_315.t1 104.842
R86 a_1526_315.n5 a_1526_315.n4 101.793
R87 a_1526_315.n2 a_1526_315.n1 101.669
R88 a_1526_315.n1 a_1526_315.n0 61.345
R89 a_1526_315.n3 a_1526_315.n2 20.762
R90 a_1526_315.n5 a_1526_315.n3 1.939
R91 VGND.n26 VGND.t2 162.682
R92 VGND.n7 VGND.t5 146.638
R93 VGND.n2 VGND.n1 126.005
R94 VGND.n0 VGND.t3 117.624
R95 VGND.n42 VGND.n41 107.239
R96 VGND.n18 VGND.n17 107.029
R97 VGND.n35 VGND.n34 106.463
R98 VGND.n17 VGND.t6 87.142
R99 VGND.n17 VGND.t7 66.294
R100 VGND.n34 VGND.t10 61.428
R101 VGND.n34 VGND.t0 40
R102 VGND.n41 VGND.t8 38.571
R103 VGND.n41 VGND.t1 38.571
R104 VGND.n1 VGND.t9 28.615
R105 VGND.n1 VGND.t4 27.692
R106 VGND.n4 VGND.n3 4.65
R107 VGND.n6 VGND.n5 4.65
R108 VGND.n8 VGND.n7 4.65
R109 VGND.n10 VGND.n9 4.65
R110 VGND.n12 VGND.n11 4.65
R111 VGND.n14 VGND.n13 4.65
R112 VGND.n16 VGND.n15 4.65
R113 VGND.n19 VGND.n18 4.65
R114 VGND.n21 VGND.n20 4.65
R115 VGND.n23 VGND.n22 4.65
R116 VGND.n25 VGND.n24 4.65
R117 VGND.n27 VGND.n26 4.65
R118 VGND.n29 VGND.n28 4.65
R119 VGND.n31 VGND.n30 4.65
R120 VGND.n33 VGND.n32 4.65
R121 VGND.n36 VGND.n35 4.65
R122 VGND.n38 VGND.n37 4.65
R123 VGND.n40 VGND.n39 4.65
R124 VGND.n43 VGND.n42 3.932
R125 VGND.n3 VGND.n2 1.505
R126 VGND.n4 VGND.n0 0.861
R127 VGND.n43 VGND.n40 0.137
R128 VGND VGND.n43 0.123
R129 VGND.n6 VGND.n4 0.119
R130 VGND.n8 VGND.n6 0.119
R131 VGND.n10 VGND.n8 0.119
R132 VGND.n12 VGND.n10 0.119
R133 VGND.n14 VGND.n12 0.119
R134 VGND.n16 VGND.n14 0.119
R135 VGND.n19 VGND.n16 0.119
R136 VGND.n21 VGND.n19 0.119
R137 VGND.n23 VGND.n21 0.119
R138 VGND.n25 VGND.n23 0.119
R139 VGND.n27 VGND.n25 0.119
R140 VGND.n29 VGND.n27 0.119
R141 VGND.n31 VGND.n29 0.119
R142 VGND.n33 VGND.n31 0.119
R143 VGND.n36 VGND.n33 0.119
R144 VGND.n38 VGND.n36 0.119
R145 VGND.n40 VGND.n38 0.119
R146 Q.n3 Q.n2 292.5
R147 Q.n4 Q.n3 146.523
R148 Q Q.n0 93.613
R149 Q.n1 Q.n0 92.5
R150 Q.n2 Q.n1 59.366
R151 Q.n3 Q.t3 26.595
R152 Q.n3 Q.t2 26.595
R153 Q.n0 Q.t0 24.923
R154 Q.n0 Q.t1 24.923
R155 Q.n1 Q 11.501
R156 Q.n4 Q 9.678
R157 Q.n2 Q 5.75
R158 Q Q.n4 2.881
R159 VNB.t5 VNB.t12 6916.22
R160 VNB.t11 VNB.t14 6211.76
R161 VNB.t7 VNB.t13 5321.88
R162 VNB VNB.t1 4270.59
R163 VNB.t9 VNB.t10 4003.85
R164 VNB.t12 VNB.t4 3406.45
R165 VNB.t3 VNB.t2 3332.35
R166 VNB.t14 VNB.t0 3267.65
R167 VNB.t16 VNB.t15 3105.88
R168 VNB.t2 VNB.t7 3073.53
R169 VNB.t4 VNB.t9 3062.58
R170 VNB.t1 VNB.t11 2717.65
R171 VNB.t0 VNB.t16 2523.53
R172 VNB.t15 VNB.t5 2458.82
R173 VNB.t10 VNB.t3 2363.68
R174 VNB.t13 VNB.t8 2200
R175 VNB.t8 VNB.t6 2030.77
R176 a_193_47.t0 a_193_47.n3 278.596
R177 a_193_47.n0 a_193_47.t4 272.659
R178 a_193_47.n1 a_193_47.t2 268.057
R179 a_193_47.n1 a_193_47.t5 206.98
R180 a_193_47.n0 a_193_47.t3 195.261
R181 a_193_47.n3 a_193_47.t1 150.159
R182 a_193_47.n2 a_193_47.n0 14.375
R183 a_193_47.n3 a_193_47.n2 7.846
R184 a_193_47.n2 a_193_47.n1 4.65
R185 a_559_369.n3 a_559_369.n2 414.098
R186 a_559_369.n2 a_559_369.t1 395.981
R187 a_559_369.n1 a_559_369.n0 208.075
R188 a_559_369.n1 a_559_369.t3 163.742
R189 a_559_369.n2 a_559_369.n1 72.282
R190 a_559_369.n0 a_559_369.t5 54.285
R191 a_559_369.t0 a_559_369.n3 41.554
R192 a_559_369.n3 a_559_369.t2 41.554
R193 a_559_369.n0 a_559_369.t4 40
R194 a_939_413.n3 a_939_413.n2 400.546
R195 a_939_413.n0 a_939_413.t4 226.539
R196 a_939_413.n2 a_939_413.n1 207.742
R197 a_939_413.n0 a_939_413.t5 196.013
R198 a_939_413.n2 a_939_413.n0 92.738
R199 a_939_413.n3 a_939_413.t2 75.047
R200 a_939_413.t0 a_939_413.n3 72.702
R201 a_939_413.n1 a_939_413.t3 65
R202 a_939_413.n1 a_939_413.t1 45
R203 a_1098_183.n1 a_1098_183.t4 433.799
R204 a_1098_183.n3 a_1098_183.n2 381.512
R205 a_1098_183.n1 a_1098_183.t5 128.098
R206 a_1098_183.n2 a_1098_183.n0 125.628
R207 a_1098_183.n2 a_1098_183.n1 109.306
R208 a_1098_183.n3 a_1098_183.t0 89.119
R209 a_1098_183.n0 a_1098_183.t1 63.333
R210 a_1098_183.t3 a_1098_183.n3 37.523
R211 a_1098_183.n0 a_1098_183.t2 36.77
R212 a_1355_413.n3 a_1355_413.n2 400.947
R213 a_1355_413.n0 a_1355_413.t4 212.079
R214 a_1355_413.n2 a_1355_413.n0 173.92
R215 a_1355_413.n2 a_1355_413.n1 151.491
R216 a_1355_413.n0 a_1355_413.t5 139.779
R217 a_1355_413.n1 a_1355_413.t2 73.333
R218 a_1355_413.n3 a_1355_413.t3 63.321
R219 a_1355_413.t0 a_1355_413.n3 63.321
R220 a_1355_413.n1 a_1355_413.t1 48.333
R221 a_1484_47.t1 a_1484_47.t0 93.059
R222 SCE.n1 SCE.t2 321.304
R223 SCE.n2 SCE.t3 265.907
R224 SCE.n0 SCE.t1 237.785
R225 SCE.n2 SCE.n1 177.27
R226 SCE.n0 SCE.t0 174.833
R227 SCE SCE.n2 20.114
R228 SCE.n1 SCE.n0 8.763
R229 a_299_47.t1 a_299_47.n1 343.828
R230 a_299_47.n0 a_299_47.t3 340.555
R231 a_299_47.n0 a_299_47.t2 305.648
R232 a_299_47.n1 a_299_47.t0 251.534
R233 a_299_47.n1 a_299_47.n0 29.469
R234 CLK.n0 CLK.t0 294.554
R235 CLK.n0 CLK.t1 209.401
R236 CLK.n1 CLK.n0 76
R237  CLK.n1 10.422
R238 CLK.n1 CLK 2.011
R239 a_27_47.n0 a_27_47.t3 510.42
R240 a_27_47.n1 a_27_47.t6 448.258
R241 a_27_47.n3 a_27_47.t7 263.171
R242 a_27_47.n1 a_27_47.t5 254.388
R243 a_27_47.t1 a_27_47.n5 243.779
R244 a_27_47.n3 a_27_47.t2 227.825
R245 a_27_47.n4 a_27_47.t0 198.368
R246 a_27_47.n0 a_27_47.t4 137.905
R247 a_27_47.n2 a_27_47.n1 112.815
R248 a_27_47.n4 a_27_47.n3 76
R249 a_27_47.n5 a_27_47.n4 35.339
R250 a_27_47.n2 a_27_47.n0 10.445
R251 a_27_47.n5 a_27_47.n2 8.608
R252 a_467_369.t0 a_467_369.t1 95.421
R253 a_1439_413.t0 a_1439_413.t1 204.035
R254 a_486_47.t0 a_486_47.t1 68.571
R255 a_1032_413.t0 a_1032_413.t1 154.785
R256 D.n0 D.t1 321.868
R257 D.n0 D.t0 183.694
R258 D D.n0 83.757
R259 a_1036_47.t0 a_1036_47.t1 98.059
R260 a_660_47.t0 a_660_47.t1 65.714
C0 VPB VPWR 0.21fF
C1 VPWR Q 0.31fF
C2 VGND Q 0.21fF
C3 VPWR VGND 0.13fF
C4 SCE VGND 0.15fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__sdfxtp_4.ext - technology: sky130A

.subckt sky130_fd_sc_hd__sdfxtp_4 VGND VPWR SCD D SCE CLK Q VNB VPB
X0 Q.t3 a_1527_315.t2 VPWR.t8 VPB.t12 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_466_369.t1 SCE.t0 VPWR.t11 VPB.t15 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X2 VPWR.t7 a_1527_315.t3 Q.t2 VPB.t11 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 a_1356_413.t2 a_193_47.t2 a_1099_183.t3 VNB.t7 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X4 VPWR.t2 SCD.t0 a_644_369.t0 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X5 VPWR.t12 SCE.t1 a_299_47.t0 VPB.t16 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X6 Q.t1 a_1527_315.t4 VPWR.t6 VPB.t10 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 a_940_413.t2 a_193_47.t3 a_560_369.t2 VPB.t17 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 VPWR.t1 CLK.t0 a_27_47.t0 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X9 a_487_47.t1 a_299_47.t2 VGND.t11 VNB.t8 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10 VPWR.t9 a_1356_413.t4 a_1527_315.t0 VPB.t13 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 a_1099_183.t0 a_940_413.t4 VGND.t8 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X12 a_193_47.t0 a_27_47.t2 VGND.t2 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13 Q.t7 a_1527_315.t5 VGND.t6 VNB.t15 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14 VPWR.t4 a_1527_315.t6 a_1440_413.t1 VPB.t9 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15 VGND.t9 a_1356_413.t5 a_1527_315.t1 VNB.t16 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X16 a_940_413.t3 a_27_47.t3 a_560_369.t3 VNB.t9 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X17 VPWR.t10 a_1099_183.t4 a_1033_413.t0 VPB.t14 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18 VGND.t0 a_1099_183.t5 a_1037_47.t0 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19 VGND.t10 SCE.t2 a_299_47.t1 VNB.t18 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20 VGND.t7 a_1527_315.t7 a_1485_47.t1 VNB.t14 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21 Q.t6 a_1527_315.t8 VGND.t5 VNB.t13 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X22 a_644_369.t1 a_299_47.t3 a_560_369.t5 VPB.t7 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X23 a_661_47.t1 SCE.t3 a_560_369.t4 VNB.t17 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24 VGND.t1 SCD.t1 a_661_47.t0 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X25 VGND.t4 a_1527_315.t9 Q.t5 VNB.t12 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X26 a_560_369.t0 D.t0 a_466_369.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X27 a_1485_47.t0 a_27_47.t4 a_1356_413.t3 VNB.t10 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X28 a_560_369.t1 D.t1 a_487_47.t0 VNB.t5 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X29 VPWR.t5 a_1527_315.t10 Q.t0 VPB.t8 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X30 a_1033_413.t1 a_27_47.t5 a_940_413.t0 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X31 a_1037_47.t1 a_193_47.t4 a_940_413.t1 VNB.t6 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X32 a_193_47.t1 a_27_47.t6 VPWR.t3 VPB.t5 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X33 a_1099_183.t1 a_940_413.t5 VPWR.t0 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X34 a_1440_413.t0 a_193_47.t5 a_1356_413.t1 VPB.t18 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X35 VGND.t12 CLK.t1 a_27_47.t1 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X36 a_1356_413.t0 a_27_47.t7 a_1099_183.t2 VPB.t6 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X37 VGND.t3 a_1527_315.t11 Q.t4 VNB.t11 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
R0 a_1527_315.n12 a_1527_315.t7 383.498
R1 a_1527_315.n0 a_1527_315.t10 212.079
R2 a_1527_315.n2 a_1527_315.t2 212.079
R3 a_1527_315.n5 a_1527_315.t3 212.079
R4 a_1527_315.n8 a_1527_315.t4 212.079
R5 a_1527_315.t0 a_1527_315.n13 178.588
R6 a_1527_315.n0 a_1527_315.t11 139.779
R7 a_1527_315.n2 a_1527_315.t8 139.779
R8 a_1527_315.n5 a_1527_315.t9 139.779
R9 a_1527_315.n8 a_1527_315.t5 139.779
R10 a_1527_315.n12 a_1527_315.t6 139.285
R11 a_1527_315.n11 a_1527_315.t1 109.638
R12 a_1527_315.n13 a_1527_315.n12 103.927
R13 a_1527_315.n4 a_1527_315.n1 93.408
R14 a_1527_315.n10 a_1527_315.n9 76
R15 a_1527_315.n4 a_1527_315.n3 76
R16 a_1527_315.n7 a_1527_315.n6 76
R17 a_1527_315.n11 a_1527_315.n10 32.768
R18 a_1527_315.n1 a_1527_315.n0 27.751
R19 a_1527_315.n13 a_1527_315.n11 19.236
R20 a_1527_315.n7 a_1527_315.n4 17.408
R21 a_1527_315.n10 a_1527_315.n7 17.408
R22 a_1527_315.n3 a_1527_315.n2 16.066
R23 a_1527_315.n9 a_1527_315.n8 8.763
R24 a_1527_315.n6 a_1527_315.n5 2.921
R25 VPWR.n30 VPWR.t2 429.516
R26 VPWR.n10 VPWR.t4 425.042
R27 VPWR.n47 VPWR.n46 311.893
R28 VPWR.n40 VPWR.n39 307.627
R29 VPWR.n2 VPWR.t5 208.892
R30 VPWR.n6 VPWR.n5 190.72
R31 VPWR.n19 VPWR.n18 174.594
R32 VPWR.n1 VPWR.n0 173.841
R33 VPWR.n18 VPWR.t10 113.978
R34 VPWR.n39 VPWR.t11 41.554
R35 VPWR.n39 VPWR.t12 41.554
R36 VPWR.n46 VPWR.t3 41.554
R37 VPWR.n46 VPWR.t1 41.554
R38 VPWR.n18 VPWR.t0 35.46
R39 VPWR.n5 VPWR.t9 33.49
R40 VPWR.n5 VPWR.t6 30.535
R41 VPWR.n0 VPWR.t7 28.565
R42 VPWR.n0 VPWR.t8 26.595
R43 VPWR.n20 VPWR.n19 14.305
R44 VPWR.n31 VPWR.n30 4.894
R45 VPWR.n2 VPWR.n1 4.763
R46 VPWR.n4 VPWR.n3 4.65
R47 VPWR.n7 VPWR.n6 4.65
R48 VPWR.n9 VPWR.n8 4.65
R49 VPWR.n11 VPWR.n10 4.65
R50 VPWR.n13 VPWR.n12 4.65
R51 VPWR.n15 VPWR.n14 4.65
R52 VPWR.n17 VPWR.n16 4.65
R53 VPWR.n21 VPWR.n20 4.65
R54 VPWR.n23 VPWR.n22 4.65
R55 VPWR.n25 VPWR.n24 4.65
R56 VPWR.n27 VPWR.n26 4.65
R57 VPWR.n29 VPWR.n28 4.65
R58 VPWR.n32 VPWR.n31 4.65
R59 VPWR.n34 VPWR.n33 4.65
R60 VPWR.n36 VPWR.n35 4.65
R61 VPWR.n38 VPWR.n37 4.65
R62 VPWR.n41 VPWR.n40 4.65
R63 VPWR.n43 VPWR.n42 4.65
R64 VPWR.n45 VPWR.n44 4.65
R65 VPWR.n48 VPWR.n47 3.941
R66 VPWR.n4 VPWR.n2 0.262
R67 VPWR.n48 VPWR.n45 0.137
R68 VPWR VPWR.n48 0.123
R69 VPWR.n7 VPWR.n4 0.119
R70 VPWR.n9 VPWR.n7 0.119
R71 VPWR.n11 VPWR.n9 0.119
R72 VPWR.n13 VPWR.n11 0.119
R73 VPWR.n15 VPWR.n13 0.119
R74 VPWR.n17 VPWR.n15 0.119
R75 VPWR.n21 VPWR.n17 0.119
R76 VPWR.n23 VPWR.n21 0.119
R77 VPWR.n25 VPWR.n23 0.119
R78 VPWR.n27 VPWR.n25 0.119
R79 VPWR.n29 VPWR.n27 0.119
R80 VPWR.n32 VPWR.n29 0.119
R81 VPWR.n34 VPWR.n32 0.119
R82 VPWR.n36 VPWR.n34 0.119
R83 VPWR.n38 VPWR.n36 0.119
R84 VPWR.n41 VPWR.n38 0.119
R85 VPWR.n43 VPWR.n41 0.119
R86 VPWR.n45 VPWR.n43 0.119
R87 Q.n2 Q.n0 145.235
R88 Q.n2 Q.n1 106.083
R89 Q.n5 Q.n3 91.776
R90 Q.n5 Q.n4 52.624
R91 Q Q.n2 34.998
R92 Q.n0 Q.t2 26.595
R93 Q.n0 Q.t1 26.595
R94 Q.n1 Q.t0 26.595
R95 Q.n1 Q.t3 26.595
R96 Q Q.n5 26.465
R97 Q.n3 Q.t5 24.923
R98 Q.n3 Q.t7 24.923
R99 Q.n4 Q.t4 24.923
R100 Q.n4 Q.t6 24.923
R101 VPB.t9 VPB.t13 624.454
R102 VPB.t3 VPB.t17 600.778
R103 VPB.t5 VPB.t16 556.386
R104 VPB.t14 VPB.t1 390.654
R105 VPB.t18 VPB.t9 346.261
R106 VPB.t4 VPB.t14 284.112
R107 VPB.t13 VPB.t10 281.152
R108 VPB.t1 VPB.t6 281.152
R109 VPB.t15 VPB.t0 278.193
R110 VPB.t17 VPB.t4 275.233
R111 VPB.t7 VPB.t3 275.233
R112 VPB.t11 VPB.t12 254.517
R113 VPB.t12 VPB.t8 248.598
R114 VPB.t10 VPB.t11 248.598
R115 VPB.t6 VPB.t18 248.598
R116 VPB.t0 VPB.t7 248.598
R117 VPB.t16 VPB.t15 248.598
R118 VPB.t2 VPB.t5 248.598
R119 VPB VPB.t2 145.015
R120 SCE.n1 SCE.t2 321.771
R121 SCE.n2 SCE.t3 266.283
R122 SCE.n0 SCE.t0 236.179
R123 SCE.n2 SCE.n1 177.27
R124 SCE.n0 SCE.t1 174.833
R125 SCE SCE.n2 20.114
R126 SCE.n1 SCE.n0 8.763
R127 a_466_369.t0 a_466_369.t1 98.5
R128 a_193_47.t1 a_193_47.n3 278.596
R129 a_193_47.n0 a_193_47.t5 272.659
R130 a_193_47.n1 a_193_47.t3 268.251
R131 a_193_47.n1 a_193_47.t4 206.786
R132 a_193_47.n0 a_193_47.t2 195.261
R133 a_193_47.n3 a_193_47.t0 150.159
R134 a_193_47.n2 a_193_47.n0 14.749
R135 a_193_47.n3 a_193_47.n2 7.85
R136 a_193_47.n2 a_193_47.n1 4.65
R137 a_1099_183.n1 a_1099_183.t4 433.799
R138 a_1099_183.n3 a_1099_183.n2 381.512
R139 a_1099_183.n1 a_1099_183.t5 128.098
R140 a_1099_183.n2 a_1099_183.n0 125.628
R141 a_1099_183.n2 a_1099_183.n1 109.306
R142 a_1099_183.n3 a_1099_183.t2 89.119
R143 a_1099_183.n0 a_1099_183.t3 63.333
R144 a_1099_183.t1 a_1099_183.n3 37.523
R145 a_1099_183.n0 a_1099_183.t0 36.77
R146 a_1356_413.n3 a_1356_413.n2 400.947
R147 a_1356_413.n0 a_1356_413.t4 212.079
R148 a_1356_413.n2 a_1356_413.n0 173.92
R149 a_1356_413.n2 a_1356_413.n1 151.491
R150 a_1356_413.n0 a_1356_413.t5 139.779
R151 a_1356_413.n1 a_1356_413.t2 73.333
R152 a_1356_413.n3 a_1356_413.t1 63.321
R153 a_1356_413.t0 a_1356_413.n3 63.321
R154 a_1356_413.n1 a_1356_413.t3 48.333
R155 VNB.t4 VNB.t9 6916.22
R156 VNB.t3 VNB.t18 6211.76
R157 VNB.t14 VNB.t16 5321.88
R158 VNB VNB.t0 4270.59
R159 VNB.t2 VNB.t1 4003.85
R160 VNB.t9 VNB.t6 3406.45
R161 VNB.t7 VNB.t10 3332.35
R162 VNB.t18 VNB.t8 3300
R163 VNB.t5 VNB.t17 3105.88
R164 VNB.t10 VNB.t14 3073.53
R165 VNB.t6 VNB.t2 3062.58
R166 VNB.t0 VNB.t3 2717.65
R167 VNB.t8 VNB.t5 2523.53
R168 VNB.t17 VNB.t4 2458.82
R169 VNB.t1 VNB.t7 2363.68
R170 VNB.t16 VNB.t15 2296.7
R171 VNB.t12 VNB.t13 2079.12
R172 VNB.t13 VNB.t11 2030.77
R173 VNB.t15 VNB.t12 2030.77
R174 SCD.n0 SCD.t1 268.848
R175 SCD.n0 SCD.t0 236.714
R176 SCD SCD.n0 82.53
R177 a_644_369.t0 a_644_369.t1 96.96
R178 a_299_47.t0 a_299_47.n1 343.828
R179 a_299_47.n0 a_299_47.t3 340.853
R180 a_299_47.n0 a_299_47.t2 306.024
R181 a_299_47.n1 a_299_47.t1 251.534
R182 a_299_47.n1 a_299_47.n0 29.469
R183 a_560_369.n3 a_560_369.n2 414.098
R184 a_560_369.n2 a_560_369.t2 395.981
R185 a_560_369.n1 a_560_369.n0 208.075
R186 a_560_369.n1 a_560_369.t3 163.742
R187 a_560_369.n2 a_560_369.n1 72.282
R188 a_560_369.n0 a_560_369.t1 54.285
R189 a_560_369.n3 a_560_369.t5 41.554
R190 a_560_369.t0 a_560_369.n3 41.554
R191 a_560_369.n0 a_560_369.t4 40
R192 a_940_413.n3 a_940_413.n2 400.546
R193 a_940_413.n0 a_940_413.t4 226.539
R194 a_940_413.n2 a_940_413.n1 207.742
R195 a_940_413.n0 a_940_413.t5 196.013
R196 a_940_413.n2 a_940_413.n0 92.738
R197 a_940_413.n3 a_940_413.t2 75.047
R198 a_940_413.t0 a_940_413.n3 72.702
R199 a_940_413.n1 a_940_413.t3 65
R200 a_940_413.n1 a_940_413.t1 45
R201 CLK.n0 CLK.t0 294.554
R202 CLK.n0 CLK.t1 209.401
R203 CLK CLK.n0 78.067
R204 a_27_47.n0 a_27_47.t3 510.426
R205 a_27_47.n1 a_27_47.t4 448.258
R206 a_27_47.n3 a_27_47.t6 263.171
R207 a_27_47.n1 a_27_47.t7 254.388
R208 a_27_47.t0 a_27_47.n5 243.779
R209 a_27_47.n3 a_27_47.t2 227.825
R210 a_27_47.n4 a_27_47.t1 198.368
R211 a_27_47.n0 a_27_47.t5 137.901
R212 a_27_47.n2 a_27_47.n1 112.811
R213 a_27_47.n4 a_27_47.n3 76
R214 a_27_47.n5 a_27_47.n4 35.339
R215 a_27_47.n2 a_27_47.n0 10.451
R216 a_27_47.n5 a_27_47.n2 8.64
R217 VGND.n2 VGND.t3 199.014
R218 VGND.n30 VGND.t1 162.682
R219 VGND.n11 VGND.t7 146.638
R220 VGND.n6 VGND.n5 126.005
R221 VGND.n1 VGND.n0 115.841
R222 VGND.n46 VGND.n45 107.239
R223 VGND.n22 VGND.n21 107.029
R224 VGND.n39 VGND.n38 106.463
R225 VGND.n21 VGND.t0 87.142
R226 VGND.n21 VGND.t8 66.294
R227 VGND.n38 VGND.t10 61.428
R228 VGND.n38 VGND.t11 41.428
R229 VGND.n45 VGND.t2 38.571
R230 VGND.n45 VGND.t12 38.571
R231 VGND.n5 VGND.t9 31.384
R232 VGND.n5 VGND.t6 28.615
R233 VGND.n0 VGND.t4 26.769
R234 VGND.n0 VGND.t5 24.923
R235 VGND.n2 VGND.n1 4.763
R236 VGND.n4 VGND.n3 4.65
R237 VGND.n8 VGND.n7 4.65
R238 VGND.n10 VGND.n9 4.65
R239 VGND.n12 VGND.n11 4.65
R240 VGND.n14 VGND.n13 4.65
R241 VGND.n16 VGND.n15 4.65
R242 VGND.n18 VGND.n17 4.65
R243 VGND.n20 VGND.n19 4.65
R244 VGND.n23 VGND.n22 4.65
R245 VGND.n25 VGND.n24 4.65
R246 VGND.n27 VGND.n26 4.65
R247 VGND.n29 VGND.n28 4.65
R248 VGND.n31 VGND.n30 4.65
R249 VGND.n33 VGND.n32 4.65
R250 VGND.n35 VGND.n34 4.65
R251 VGND.n37 VGND.n36 4.65
R252 VGND.n40 VGND.n39 4.65
R253 VGND.n42 VGND.n41 4.65
R254 VGND.n44 VGND.n43 4.65
R255 VGND.n47 VGND.n46 3.932
R256 VGND.n7 VGND.n6 3.011
R257 VGND.n4 VGND.n2 0.262
R258 VGND.n47 VGND.n44 0.137
R259 VGND VGND.n47 0.123
R260 VGND.n8 VGND.n4 0.119
R261 VGND.n10 VGND.n8 0.119
R262 VGND.n12 VGND.n10 0.119
R263 VGND.n14 VGND.n12 0.119
R264 VGND.n16 VGND.n14 0.119
R265 VGND.n18 VGND.n16 0.119
R266 VGND.n20 VGND.n18 0.119
R267 VGND.n23 VGND.n20 0.119
R268 VGND.n25 VGND.n23 0.119
R269 VGND.n27 VGND.n25 0.119
R270 VGND.n29 VGND.n27 0.119
R271 VGND.n31 VGND.n29 0.119
R272 VGND.n33 VGND.n31 0.119
R273 VGND.n35 VGND.n33 0.119
R274 VGND.n37 VGND.n35 0.119
R275 VGND.n40 VGND.n37 0.119
R276 VGND.n42 VGND.n40 0.119
R277 VGND.n44 VGND.n42 0.119
R278 a_487_47.t0 a_487_47.t1 68.571
R279 a_1440_413.t0 a_1440_413.t1 204.035
R280 a_1033_413.t0 a_1033_413.t1 154.785
R281 a_1037_47.t0 a_1037_47.t1 98.059
R282 a_1485_47.t1 a_1485_47.t0 93.059
R283 a_661_47.t0 a_661_47.t1 65.714
R284 D.n0 D.t1 321.868
R285 D.n0 D.t0 183.694
R286 D D.n0 82.206
C0 VGND Q 0.39fF
C1 VPWR VGND 0.13fF
C2 SCE VGND 0.15fF
C3 VPB VPWR 0.22fF
C4 VPWR Q 0.52fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__sdlclkp_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__sdlclkp_1 SCE CLK GCLK GATE VGND VPWR VNB VPB
X0 a_1094_47.t0 a_464_315.t2 a_1012_47.t0 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1 a_464_315.t0 a_286_413.t4 VPWR.t2 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 a_464_315.t1 a_286_413.t5 VGND.t1 VNB.t9 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 VPWR.t3 CLK.t0 a_1012_47.t2 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X4 a_1012_47.t1 a_464_315.t3 VPWR.t1 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X5 a_109_369.t0 SCE.t0 VPWR.t5 VPB.t5 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X6 VPWR.t0 a_464_315.t4 a_382_413.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7 a_382_413.t1 a_256_147.t2 a_286_413.t1 VPB.t6 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 a_286_413.t2 a_256_243.t2 a_27_47.t4 VPB.t10 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9 a_27_47.t1 GATE.t0 VGND.t5 VNB.t6 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10 a_256_147.t0 CLK.t1 VPWR.t4 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X11 VGND.t4 a_256_147.t3 a_256_243.t1 VNB.t5 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12 GCLK.t0 a_1012_47.t3 VPWR.t7 VPB.t8 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13 a_27_47.t2 GATE.t1 a_109_369.t1 VPB.t9 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X14 a_256_147.t1 CLK.t2 VGND.t3 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15 GCLK.t1 a_1012_47.t4 VGND.t6 VNB.t7 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X16 VPWR.t6 a_256_147.t4 a_256_243.t0 VPB.t7 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X17 a_286_413.t0 a_256_147.t5 a_27_47.t3 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X18 VGND.t2 CLK.t3 a_1094_47.t1 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19 a_394_47.t1 a_256_243.t3 a_286_413.t3 VNB.t10 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X20 VGND.t0 a_464_315.t5 a_394_47.t0 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21 VGND.t7 SCE.t1 a_27_47.t0 VNB.t8 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
R0 a_464_315.n1 a_464_315.t5 392.561
R1 a_464_315.n0 a_464_315.t2 321.771
R2 a_464_315.n4 a_464_315.n3 309.954
R3 a_464_315.n2 a_464_315.t1 227.805
R4 a_464_315.n3 a_464_315.n0 226.83
R5 a_464_315.n0 a_464_315.t3 183.597
R6 a_464_315.n4 a_464_315.t0 175.531
R7 a_464_315.n1 a_464_315.t4 148.348
R8 a_464_315.n2 a_464_315.n1 115.585
R9 a_464_315.n5 a_464_315.n4 15.153
R10 a_464_315.n3 a_464_315.n2 5.527
R11 a_1012_47.n2 a_1012_47.n1 332.537
R12 a_1012_47.n1 a_1012_47.t0 242.189
R13 a_1012_47.n0 a_1012_47.t3 241.534
R14 a_1012_47.n0 a_1012_47.t4 169.234
R15 a_1012_47.n1 a_1012_47.n0 76
R16 a_1012_47.n2 a_1012_47.t2 41.554
R17 a_1012_47.t1 a_1012_47.n2 41.554
R18 a_1094_47.t0 a_1094_47.t1 117.142
R19 VNB VNB.t8 6470.59
R20 VNB.t3 VNB.t1 6082.35
R21 VNB.t9 VNB.t5 5321.88
R22 VNB.t10 VNB.t0 3947.06
R23 VNB.t1 VNB.t2 3623.53
R24 VNB.t4 VNB.t10 3397.06
R25 VNB.t6 VNB.t4 3105.88
R26 VNB.t0 VNB.t9 2811.39
R27 VNB.t5 VNB.t3 2717.65
R28 VNB.t8 VNB.t6 2717.65
R29 VNB.t2 VNB.t7 2255.35
R30 a_286_413.n3 a_286_413.n2 387.22
R31 a_286_413.n1 a_286_413.t4 232.471
R32 a_286_413.n2 a_286_413.n0 162.792
R33 a_286_413.n1 a_286_413.t5 160.171
R34 a_286_413.n2 a_286_413.n1 93.347
R35 a_286_413.t1 a_286_413.n3 77.392
R36 a_286_413.n3 a_286_413.t2 77.392
R37 a_286_413.n0 a_286_413.t3 63.333
R38 a_286_413.n0 a_286_413.t0 61.666
R39 VPWR.n8 VPWR.n7 438.28
R40 VPWR.n2 VPWR.t1 425.096
R41 VPWR.n1 VPWR.n0 309.368
R42 VPWR.n16 VPWR.n15 292.5
R43 VPWR.n29 VPWR.t5 233.522
R44 VPWR.n15 VPWR.t0 136.023
R45 VPWR.n15 VPWR.t2 78.565
R46 VPWR.n7 VPWR.t4 61.562
R47 VPWR.n7 VPWR.t6 61.562
R48 VPWR.n0 VPWR.t3 50.789
R49 VPWR.n0 VPWR.t7 39.3
R50 VPWR.n4 VPWR.n3 4.65
R51 VPWR.n6 VPWR.n5 4.65
R52 VPWR.n10 VPWR.n9 4.65
R53 VPWR.n12 VPWR.n11 4.65
R54 VPWR.n14 VPWR.n13 4.65
R55 VPWR.n18 VPWR.n17 4.65
R56 VPWR.n20 VPWR.n19 4.65
R57 VPWR.n22 VPWR.n21 4.65
R58 VPWR.n24 VPWR.n23 4.65
R59 VPWR.n26 VPWR.n25 4.65
R60 VPWR.n28 VPWR.n27 4.65
R61 VPWR.n30 VPWR.n29 4.65
R62 VPWR.n17 VPWR.n16 3.506
R63 VPWR.n9 VPWR.n8 1.396
R64 VPWR.n3 VPWR.n2 0.814
R65 VPWR.n4 VPWR.n1 0.76
R66 VPWR.n6 VPWR.n4 0.119
R67 VPWR.n10 VPWR.n6 0.119
R68 VPWR.n12 VPWR.n10 0.119
R69 VPWR.n14 VPWR.n12 0.119
R70 VPWR.n18 VPWR.n14 0.119
R71 VPWR.n20 VPWR.n18 0.119
R72 VPWR.n22 VPWR.n20 0.119
R73 VPWR.n24 VPWR.n22 0.119
R74 VPWR.n26 VPWR.n24 0.119
R75 VPWR.n28 VPWR.n26 0.119
R76 VPWR.n30 VPWR.n28 0.119
R77 VPWR VPWR.n30 0.022
R78 VPB.t4 VPB.t1 562.305
R79 VPB.t2 VPB.t7 550.467
R80 VPB.t0 VPB.t2 402.492
R81 VPB.t6 VPB.t0 349.221
R82 VPB.t7 VPB.t4 325.545
R83 VPB.t9 VPB.t10 310.747
R84 VPB.t10 VPB.t6 284.112
R85 VPB.t3 VPB.t8 281.152
R86 VPB.t1 VPB.t3 248.598
R87 VPB.t5 VPB.t9 213.084
R88 VPB VPB.t5 192.367
R89 VGND.n9 VGND.n8 111.421
R90 VGND.n1 VGND.n0 106.463
R91 VGND.n20 VGND.n19 106.463
R92 VGND.n3 VGND.n2 96.655
R93 VGND.n8 VGND.t0 65.714
R94 VGND.n2 VGND.t6 41.648
R95 VGND.n8 VGND.t1 41.296
R96 VGND.n2 VGND.t2 38.571
R97 VGND.n0 VGND.t3 38.571
R98 VGND.n0 VGND.t4 38.571
R99 VGND.n19 VGND.t5 38.571
R100 VGND.n19 VGND.t7 38.571
R101 VGND.n5 VGND.n4 4.65
R102 VGND.n7 VGND.n6 4.65
R103 VGND.n10 VGND.n9 4.65
R104 VGND.n12 VGND.n11 4.65
R105 VGND.n14 VGND.n13 4.65
R106 VGND.n16 VGND.n15 4.65
R107 VGND.n18 VGND.n17 4.65
R108 VGND.n3 VGND.n1 4.099
R109 VGND.n21 VGND.n20 3.932
R110 VGND.n21 VGND.n18 0.137
R111 VGND.n5 VGND.n3 0.137
R112 VGND VGND.n21 0.123
R113 VGND.n7 VGND.n5 0.119
R114 VGND.n10 VGND.n7 0.119
R115 VGND.n12 VGND.n10 0.119
R116 VGND.n14 VGND.n12 0.119
R117 VGND.n16 VGND.n14 0.119
R118 VGND.n18 VGND.n16 0.119
R119 CLK.n0 CLK.t0 333.497
R120 CLK.n1 CLK.t1 182.814
R121 CLK.n0 CLK.t3 169.617
R122 CLK.n1 CLK.t2 149.791
R123 CLK.n3 CLK.n0 118.322
R124 CLK.n2 CLK.n1 76
R125 CLK CLK.n3 9.309
R126 CLK.n2 CLK 1.651
R127 CLK.n3 CLK.n2 1.032
R128 SCE.n0 SCE.t0 287.994
R129 SCE.n0 SCE.t1 194.808
R130 SCE.n1 SCE.n0 76
R131 SCE.n1 SCE 14.305
R132 SCE SCE.n1 2.76
R133 a_109_369.t0 a_109_369.t1 64.64
R134 a_382_413.t0 a_382_413.t1 206.38
R135 a_256_147.t0 a_256_147.n3 445.769
R136 a_256_147.n0 a_256_147.t2 230.255
R137 a_256_147.n0 a_256_147.t5 219.994
R138 a_256_147.n1 a_256_147.t3 215.731
R139 a_256_147.n1 a_256_147.t4 183.597
R140 a_256_147.n2 a_256_147.t1 173.203
R141 a_256_147.n2 a_256_147.n1 81.647
R142 a_256_147.n3 a_256_147.n2 14.268
R143 a_256_147.n3 a_256_147.n0 11.67
R144 a_256_243.n0 a_256_243.t2 552.941
R145 a_256_243.n2 a_256_243.n1 356.031
R146 a_256_243.n1 a_256_243.t1 146.004
R147 a_256_243.n2 a_256_243.t0 127.045
R148 a_256_243.n0 a_256_243.t3 121.631
R149 a_256_243.n1 a_256_243.n0 17.604
R150 a_27_47.n2 a_27_47.n1 407.566
R151 a_27_47.n1 a_27_47.t0 163.186
R152 a_27_47.n1 a_27_47.n0 144.603
R153 a_27_47.n2 a_27_47.t4 89.119
R154 a_27_47.n0 a_27_47.t3 65
R155 a_27_47.t2 a_27_47.n2 62.588
R156 a_27_47.n0 a_27_47.t1 29.534
R157 GATE.n0 GATE.t1 295.166
R158 GATE.n0 GATE.t0 201.98
R159 GATE GATE.n0 87.165
R160 GCLK.n0 GCLK.t0 207.566
R161 GCLK GCLK.t1 157.339
R162 GCLK.n0 GCLK 8.185
R163 GCLK GCLK.n0 6.859
R164 a_394_47.t0 a_394_47.t1 138.059
C0 SCE GATE 0.11fF
C1 VPB VPWR 0.15fF
C2 VPWR VGND 0.10fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__sdlclkp_2.ext - technology: sky130A

.subckt sky130_fd_sc_hd__sdlclkp_2 SCE CLK GCLK GATE VGND VPWR VNB VPB
X0 GCLK.t1 a_1020_47.t3 VPWR.t2 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_109_369.t1 SCE.t0 VPWR.t7 VPB.t10 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X2 a_465_315.t0 a_287_413.t4 VPWR.t8 VPB.t11 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 a_257_147.t0 CLK.t0 VPWR.t4 VPB.t7 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X4 a_1102_47.t1 a_465_315.t2 a_1020_47.t1 VNB.t8 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 VGND.t5 a_1020_47.t4 GCLK.t3 VNB.t6 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 a_287_413.t2 a_257_147.t2 a_27_47.t4 VNB.t11 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X7 VGND.t8 a_257_147.t3 a_257_243.t1 VNB.t10 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 VPWR.t5 a_465_315.t3 a_383_413.t0 VPB.t8 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9 VGND.t3 CLK.t1 a_1102_47.t0 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10 a_27_47.t2 GATE.t0 VGND.t1 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11 VPWR.t0 CLK.t2 a_1020_47.t0 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X12 GCLK.t2 a_1020_47.t5 VGND.t4 VNB.t5 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 a_287_413.t3 a_257_243.t2 a_27_47.t3 VPB.t6 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14 a_383_413.t1 a_257_147.t4 a_287_413.t1 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15 a_257_147.t1 CLK.t3 VGND.t2 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16 a_27_47.t0 GATE.t1 a_109_369.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X17 VPWR.t3 a_257_147.t5 a_257_243.t0 VPB.t5 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X18 a_1020_47.t2 a_465_315.t4 VPWR.t6 VPB.t9 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X19 a_395_47.t0 a_257_243.t3 a_287_413.t0 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X20 VGND.t6 a_465_315.t5 a_395_47.t1 VNB.t7 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21 VPWR.t1 a_1020_47.t6 GCLK.t0 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X22 VGND.t0 SCE.t1 a_27_47.t1 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23 a_465_315.t1 a_287_413.t5 VGND.t7 VNB.t9 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
R0 a_1020_47.n3 a_1020_47.n2 332.537
R1 a_1020_47.n2 a_1020_47.t1 245.002
R2 a_1020_47.n0 a_1020_47.t6 212.079
R3 a_1020_47.n1 a_1020_47.t3 212.079
R4 a_1020_47.n0 a_1020_47.t4 139.779
R5 a_1020_47.n1 a_1020_47.t5 139.779
R6 a_1020_47.n2 a_1020_47.n1 84.033
R7 a_1020_47.n1 a_1020_47.n0 61.345
R8 a_1020_47.t0 a_1020_47.n3 41.554
R9 a_1020_47.n3 a_1020_47.t2 41.554
R10 VPWR.n11 VPWR.n10 438.28
R11 VPWR.n5 VPWR.t6 425.096
R12 VPWR.n1 VPWR.n0 306.463
R13 VPWR.n19 VPWR.n18 292.5
R14 VPWR.n32 VPWR.t7 233.522
R15 VPWR.n2 VPWR.t1 155.222
R16 VPWR.n18 VPWR.t5 136.023
R17 VPWR.n18 VPWR.t8 78.565
R18 VPWR.n10 VPWR.t4 61.562
R19 VPWR.n10 VPWR.t3 61.562
R20 VPWR.n0 VPWR.t0 50.789
R21 VPWR.n0 VPWR.t2 39.3
R22 VPWR.n4 VPWR.n3 4.65
R23 VPWR.n7 VPWR.n6 4.65
R24 VPWR.n9 VPWR.n8 4.65
R25 VPWR.n13 VPWR.n12 4.65
R26 VPWR.n15 VPWR.n14 4.65
R27 VPWR.n17 VPWR.n16 4.65
R28 VPWR.n21 VPWR.n20 4.65
R29 VPWR.n23 VPWR.n22 4.65
R30 VPWR.n25 VPWR.n24 4.65
R31 VPWR.n27 VPWR.n26 4.65
R32 VPWR.n29 VPWR.n28 4.65
R33 VPWR.n31 VPWR.n30 4.65
R34 VPWR.n33 VPWR.n32 4.65
R35 VPWR.n2 VPWR.n1 3.788
R36 VPWR.n20 VPWR.n19 3.419
R37 VPWR.n6 VPWR.n5 1.745
R38 VPWR.n4 VPWR.n2 0.24
R39 VPWR.n12 VPWR.n11 0.232
R40 VPWR.n7 VPWR.n4 0.119
R41 VPWR.n9 VPWR.n7 0.119
R42 VPWR.n13 VPWR.n9 0.119
R43 VPWR.n15 VPWR.n13 0.119
R44 VPWR.n17 VPWR.n15 0.119
R45 VPWR.n21 VPWR.n17 0.119
R46 VPWR.n23 VPWR.n21 0.119
R47 VPWR.n25 VPWR.n23 0.119
R48 VPWR.n27 VPWR.n25 0.119
R49 VPWR.n29 VPWR.n27 0.119
R50 VPWR.n31 VPWR.n29 0.119
R51 VPWR.n33 VPWR.n31 0.119
R52 VPWR VPWR.n33 0.02
R53 GCLK.n1 GCLK.n0 143.021
R54 GCLK GCLK.n2 92.737
R55 GCLK.n3 GCLK 36.279
R56 GCLK.n3 GCLK 27.3
R57 GCLK.n0 GCLK.t0 26.595
R58 GCLK.n0 GCLK.t1 26.595
R59 GCLK.n2 GCLK.t3 24.923
R60 GCLK.n2 GCLK.t2 24.923
R61 GCLK GCLK.n3 17.23
R62 GCLK GCLK.n1 8.573
R63 GCLK.n1 GCLK 7.186
R64 VPB.t11 VPB.t5 577.102
R65 VPB.t7 VPB.t9 556.386
R66 VPB.t8 VPB.t11 402.492
R67 VPB.t4 VPB.t8 349.221
R68 VPB.t5 VPB.t7 325.545
R69 VPB.t0 VPB.t6 313.707
R70 VPB.t6 VPB.t4 284.112
R71 VPB.t1 VPB.t3 281.152
R72 VPB.t3 VPB.t2 248.598
R73 VPB.t9 VPB.t1 248.598
R74 VPB.t10 VPB.t0 213.084
R75 VPB VPB.t10 189.408
R76 SCE.n0 SCE.t0 287.994
R77 SCE.n0 SCE.t1 194.808
R78 SCE.n1 SCE.n0 76
R79 SCE.n1 SCE 14.305
R80 SCE SCE.n1 2.76
R81 a_109_369.t0 a_109_369.t1 64.64
R82 a_287_413.n3 a_287_413.n2 387.22
R83 a_287_413.n1 a_287_413.t4 232.471
R84 a_287_413.n2 a_287_413.n0 162.792
R85 a_287_413.n1 a_287_413.t5 160.171
R86 a_287_413.n2 a_287_413.n1 93.347
R87 a_287_413.t1 a_287_413.n3 77.392
R88 a_287_413.n3 a_287_413.t3 77.392
R89 a_287_413.n0 a_287_413.t0 63.333
R90 a_287_413.n0 a_287_413.t2 61.666
R91 a_465_315.t0 a_465_315.n3 471.119
R92 a_465_315.n1 a_465_315.t5 392.561
R93 a_465_315.n0 a_465_315.t2 321.771
R94 a_465_315.n3 a_465_315.n0 229.466
R95 a_465_315.n2 a_465_315.t1 227.805
R96 a_465_315.n0 a_465_315.t4 183.597
R97 a_465_315.n1 a_465_315.t3 148.348
R98 a_465_315.n2 a_465_315.n1 115.585
R99 a_465_315.n3 a_465_315.n2 5.527
R100 CLK.n0 CLK.t2 333.497
R101 CLK.n1 CLK.t0 182.814
R102 CLK.n0 CLK.t1 169.617
R103 CLK.n1 CLK.t3 146.17
R104 CLK.n3 CLK.n0 120.18
R105 CLK.n2 CLK.n1 76
R106 CLK CLK.n3 9.309
R107 CLK.n2 CLK 1.651
R108 CLK.n3 CLK.n2 1.032
R109 a_257_147.t0 a_257_147.n3 449.16
R110 a_257_147.n0 a_257_147.t4 230.255
R111 a_257_147.n0 a_257_147.t2 219.994
R112 a_257_147.n1 a_257_147.t3 215.731
R113 a_257_147.n1 a_257_147.t5 183.597
R114 a_257_147.n2 a_257_147.t1 175.94
R115 a_257_147.n2 a_257_147.n1 82.776
R116 a_257_147.n3 a_257_147.n2 17.063
R117 a_257_147.n3 a_257_147.n0 11.661
R118 a_1102_47.t0 a_1102_47.t1 60
R119 VNB VNB.t1 6438.23
R120 VNB.t3 VNB.t8 6244.12
R121 VNB.t9 VNB.t10 5321.88
R122 VNB.t0 VNB.t7 3947.06
R123 VNB.t4 VNB.t5 3623.53
R124 VNB.t11 VNB.t0 3397.06
R125 VNB.t2 VNB.t11 3138.24
R126 VNB.t7 VNB.t9 2859.74
R127 VNB.t10 VNB.t3 2717.65
R128 VNB.t1 VNB.t2 2717.65
R129 VNB.t8 VNB.t4 2329.41
R130 VNB.t5 VNB.t6 2030.77
R131 VGND.n2 VGND.t5 112.025
R132 VGND.n17 VGND.n16 111.421
R133 VGND.n10 VGND.n9 106.463
R134 VGND.n28 VGND.n27 106.463
R135 VGND.n1 VGND.n0 92.5
R136 VGND.n0 VGND.t3 78.571
R137 VGND.n16 VGND.t6 65.714
R138 VGND.n0 VGND.t4 58.791
R139 VGND.n16 VGND.t7 43.648
R140 VGND.n9 VGND.t2 38.571
R141 VGND.n9 VGND.t8 38.571
R142 VGND.n27 VGND.t1 38.571
R143 VGND.n27 VGND.t0 38.571
R144 VGND.n2 VGND.n1 5.474
R145 VGND.n4 VGND.n3 4.65
R146 VGND.n6 VGND.n5 4.65
R147 VGND.n8 VGND.n7 4.65
R148 VGND.n11 VGND.n10 4.65
R149 VGND.n13 VGND.n12 4.65
R150 VGND.n15 VGND.n14 4.65
R151 VGND.n18 VGND.n17 4.65
R152 VGND.n20 VGND.n19 4.65
R153 VGND.n22 VGND.n21 4.65
R154 VGND.n24 VGND.n23 4.65
R155 VGND.n26 VGND.n25 4.65
R156 VGND.n29 VGND.n28 3.932
R157 VGND.n4 VGND.n2 0.223
R158 VGND.n29 VGND.n26 0.137
R159 VGND VGND.n29 0.121
R160 VGND.n6 VGND.n4 0.119
R161 VGND.n8 VGND.n6 0.119
R162 VGND.n11 VGND.n8 0.119
R163 VGND.n13 VGND.n11 0.119
R164 VGND.n15 VGND.n13 0.119
R165 VGND.n18 VGND.n15 0.119
R166 VGND.n20 VGND.n18 0.119
R167 VGND.n22 VGND.n20 0.119
R168 VGND.n24 VGND.n22 0.119
R169 VGND.n26 VGND.n24 0.119
R170 a_27_47.n2 a_27_47.n1 412.029
R171 a_27_47.n1 a_27_47.t1 163.563
R172 a_27_47.n1 a_27_47.n0 143.658
R173 a_27_47.n2 a_27_47.t3 89.119
R174 a_27_47.n0 a_27_47.t4 66.666
R175 a_27_47.t0 a_27_47.n2 64.933
R176 a_27_47.n0 a_27_47.t2 28.317
R177 a_257_243.n0 a_257_243.t2 552.941
R178 a_257_243.t0 a_257_243.n1 492.58
R179 a_257_243.n1 a_257_243.t1 145.151
R180 a_257_243.n0 a_257_243.t3 121.631
R181 a_257_243.n1 a_257_243.n0 16.843
R182 a_383_413.t0 a_383_413.t1 206.38
R183 GATE.n0 GATE.t1 294.772
R184 GATE.n0 GATE.t0 201.586
R185 GATE GATE.n0 86.729
R186 a_395_47.t1 a_395_47.t0 138.059
C0 VPWR GCLK 0.27fF
C1 SCE GATE 0.11fF
C2 VPB VPWR 0.16fF
C3 VGND GCLK 0.20fF
C4 VPWR VGND 0.11fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__sdlclkp_4.ext - technology: sky130A

.subckt sky130_fd_sc_hd__sdlclkp_4 SCE CLK GCLK GATE VGND VPWR VNB VPB
X0 a_257_147.t0 CLK.t0 VPWR.t1 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1 a_109_369.t0 SCE.t0 VPWR.t8 VPB.t12 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X2 a_465_315.t0 a_287_413.t4 VPWR.t9 VPB.t13 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 VPWR.t2 a_1045_47.t3 GCLK.t3 VPB.t5 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 a_287_413.t0 a_257_147.t2 a_27_47.t2 VNB.t10 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X5 VPWR.t10 a_257_147.t3 a_257_243.t0 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X6 GCLK.t2 a_1045_47.t4 VPWR.t3 VPB.t7 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 VGND.t8 a_257_147.t4 a_257_243.t1 VNB.t9 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 VGND.t3 a_1045_47.t5 GCLK.t7 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 VPWR.t6 a_465_315.t2 a_383_413.t0 VPB.t10 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10 VPWR.t4 a_1045_47.t6 GCLK.t1 VPB.t8 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 a_1127_47.t0 a_465_315.t3 a_1045_47.t1 VNB.t6 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 a_27_47.t1 GATE.t0 VGND.t7 VNB.t8 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13 GCLK.t0 a_1045_47.t7 VPWR.t5 VPB.t9 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14 a_287_413.t2 a_257_243.t2 a_27_47.t4 VPB.t6 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15 a_383_413.t1 a_257_147.t5 a_287_413.t1 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16 VGND.t9 CLK.t1 a_1127_47.t1 VNB.t12 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X17 a_257_147.t1 CLK.t2 VGND.t10 VNB.t11 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18 GCLK.t6 a_1045_47.t8 VGND.t2 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X19 GCLK.t5 a_1045_47.t9 VGND.t1 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X20 a_27_47.t3 GATE.t1 a_109_369.t1 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X21 VPWR.t0 CLK.t3 a_1045_47.t2 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X22 a_1045_47.t0 a_465_315.t4 VPWR.t7 VPB.t11 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X23 a_395_47.t1 a_257_243.t3 a_287_413.t3 VNB.t13 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X24 VGND.t0 a_1045_47.t10 GCLK.t4 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X25 VGND.t5 a_465_315.t5 a_395_47.t0 VNB.t5 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X26 VGND.t6 SCE.t1 a_27_47.t0 VNB.t7 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X27 a_465_315.t1 a_287_413.t5 VGND.t4 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
R0 CLK.n0 CLK.t3 241.534
R1 CLK.n2 CLK.t0 181.093
R2 CLK.n0 CLK.t1 169.234
R3 CLK.n1 CLK.t2 145.671
R4 CLK.n3 CLK.n0 91.49
R5 CLK.n3 CLK.n2 9.3
R6 CLK.n2 CLK.n1 5.635
R7 CLK CLK.n4 1.551
R8 CLK.n4 CLK.n3 0.775
R9 VPWR.n10 VPWR.t7 556.339
R10 VPWR.n16 VPWR.n15 438.28
R11 VPWR.n6 VPWR.n5 306.463
R12 VPWR.n24 VPWR.n23 292.5
R13 VPWR.n37 VPWR.t8 233.522
R14 VPWR.n1 VPWR.n0 169.933
R15 VPWR.n2 VPWR.t2 161.526
R16 VPWR.n23 VPWR.t6 136.023
R17 VPWR.n23 VPWR.t9 78.565
R18 VPWR.n15 VPWR.t1 61.562
R19 VPWR.n15 VPWR.t10 61.562
R20 VPWR.n5 VPWR.t0 32.505
R21 VPWR.n5 VPWR.t5 31.52
R22 VPWR.n0 VPWR.t3 26.595
R23 VPWR.n0 VPWR.t4 26.595
R24 VPWR.n4 VPWR.n3 4.65
R25 VPWR.n7 VPWR.n6 4.65
R26 VPWR.n9 VPWR.n8 4.65
R27 VPWR.n12 VPWR.n11 4.65
R28 VPWR.n14 VPWR.n13 4.65
R29 VPWR.n18 VPWR.n17 4.65
R30 VPWR.n20 VPWR.n19 4.65
R31 VPWR.n22 VPWR.n21 4.65
R32 VPWR.n26 VPWR.n25 4.65
R33 VPWR.n28 VPWR.n27 4.65
R34 VPWR.n30 VPWR.n29 4.65
R35 VPWR.n32 VPWR.n31 4.65
R36 VPWR.n34 VPWR.n33 4.65
R37 VPWR.n36 VPWR.n35 4.65
R38 VPWR.n38 VPWR.n37 4.65
R39 VPWR.n2 VPWR.n1 3.911
R40 VPWR.n25 VPWR.n24 3.419
R41 VPWR.n11 VPWR.n10 1.396
R42 VPWR.n17 VPWR.n16 1.047
R43 VPWR.n4 VPWR.n2 0.23
R44 VPWR.n7 VPWR.n4 0.119
R45 VPWR.n9 VPWR.n7 0.119
R46 VPWR.n12 VPWR.n9 0.119
R47 VPWR.n14 VPWR.n12 0.119
R48 VPWR.n18 VPWR.n14 0.119
R49 VPWR.n20 VPWR.n18 0.119
R50 VPWR.n22 VPWR.n20 0.119
R51 VPWR.n26 VPWR.n22 0.119
R52 VPWR.n28 VPWR.n26 0.119
R53 VPWR.n30 VPWR.n28 0.119
R54 VPWR.n32 VPWR.n30 0.119
R55 VPWR.n34 VPWR.n32 0.119
R56 VPWR.n36 VPWR.n34 0.119
R57 VPWR.n38 VPWR.n36 0.119
R58 VPWR VPWR.n38 0.02
R59 a_257_147.t0 a_257_147.n3 445.769
R60 a_257_147.n0 a_257_147.t5 230.255
R61 a_257_147.n0 a_257_147.t2 219.994
R62 a_257_147.n1 a_257_147.t4 215.731
R63 a_257_147.n1 a_257_147.t3 183.597
R64 a_257_147.n2 a_257_147.t1 173.203
R65 a_257_147.n2 a_257_147.n1 81.647
R66 a_257_147.n3 a_257_147.n2 14.268
R67 a_257_147.n3 a_257_147.n0 11.679
R68 VPB.t4 VPB.t11 568.224
R69 VPB.t13 VPB.t1 556.386
R70 VPB.t10 VPB.t13 402.492
R71 VPB.t0 VPB.t10 349.221
R72 VPB.t1 VPB.t4 325.545
R73 VPB.t2 VPB.t6 313.707
R74 VPB.t6 VPB.t0 284.112
R75 VPB.t3 VPB.t9 281.152
R76 VPB.t7 VPB.t5 248.598
R77 VPB.t8 VPB.t7 248.598
R78 VPB.t9 VPB.t8 248.598
R79 VPB.t11 VPB.t3 248.598
R80 VPB.t12 VPB.t2 213.084
R81 VPB VPB.t12 189.408
R82 SCE.n0 SCE.t0 288.201
R83 SCE.n0 SCE.t1 195.015
R84 SCE.n1 SCE.n0 76
R85 SCE.n1 SCE 14.03
R86 SCE SCE.n1 2.707
R87 a_109_369.t0 a_109_369.t1 64.64
R88 a_287_413.n3 a_287_413.n2 387.22
R89 a_287_413.n1 a_287_413.t4 232.471
R90 a_287_413.n2 a_287_413.n0 162.792
R91 a_287_413.n1 a_287_413.t5 160.171
R92 a_287_413.n2 a_287_413.n1 93.347
R93 a_287_413.t1 a_287_413.n3 77.392
R94 a_287_413.n3 a_287_413.t2 77.392
R95 a_287_413.n0 a_287_413.t3 63.333
R96 a_287_413.n0 a_287_413.t0 61.666
R97 a_465_315.t0 a_465_315.n3 471.119
R98 a_465_315.n1 a_465_315.t5 392.561
R99 a_465_315.n3 a_465_315.n0 239.237
R100 a_465_315.n0 a_465_315.t4 233.007
R101 a_465_315.n2 a_465_315.t1 227.805
R102 a_465_315.n0 a_465_315.t3 160.707
R103 a_465_315.n1 a_465_315.t2 148.348
R104 a_465_315.n2 a_465_315.n1 115.585
R105 a_465_315.n3 a_465_315.n2 5.527
R106 a_1045_47.n6 a_1045_47.n5 322.579
R107 a_1045_47.n0 a_1045_47.t3 221.719
R108 a_1045_47.n1 a_1045_47.t4 221.719
R109 a_1045_47.n2 a_1045_47.t6 221.719
R110 a_1045_47.n3 a_1045_47.t7 221.719
R111 a_1045_47.n5 a_1045_47.t1 214.177
R112 a_1045_47.n0 a_1045_47.t10 149.419
R113 a_1045_47.n1 a_1045_47.t9 149.419
R114 a_1045_47.n2 a_1045_47.t5 149.419
R115 a_1045_47.n3 a_1045_47.t8 149.419
R116 a_1045_47.n5 a_1045_47.n4 76
R117 a_1045_47.n1 a_1045_47.n0 74.977
R118 a_1045_47.n2 a_1045_47.n1 74.977
R119 a_1045_47.n4 a_1045_47.n2 58.911
R120 a_1045_47.n6 a_1045_47.t2 26.595
R121 a_1045_47.t0 a_1045_47.n6 26.595
R122 a_1045_47.n4 a_1045_47.n3 16.066
R123 GCLK.n5 GCLK.n4 143.336
R124 GCLK.n1 GCLK.n0 142.77
R125 GCLK GCLK.n7 107.22
R126 GCLK GCLK.n2 95.828
R127 GCLK.n3 GCLK 54.964
R128 GCLK.n3 GCLK 46.772
R129 GCLK.n0 GCLK.t1 26.595
R130 GCLK.n0 GCLK.t0 26.595
R131 GCLK.n4 GCLK.t3 26.595
R132 GCLK.n4 GCLK.t2 26.595
R133 GCLK.n2 GCLK.t7 24.923
R134 GCLK.n2 GCLK.t6 24.923
R135 GCLK.n7 GCLK.t4 24.923
R136 GCLK.n7 GCLK.t5 24.923
R137 GCLK.n6 GCLK 14.276
R138 GCLK.n6 GCLK.n3 14.03
R139 GCLK.n6 GCLK 11.093
R140 GCLK GCLK.n1 9.243
R141 GCLK.n1 GCLK 7.748
R142 GCLK GCLK.n5 7.733
R143 GCLK.n5 GCLK 6.482
R144 GCLK GCLK.n6 3.413
R145 GCLK.n3 GCLK 2.215
R146 a_27_47.n2 a_27_47.n1 412.029
R147 a_27_47.n1 a_27_47.t0 163.563
R148 a_27_47.n1 a_27_47.n0 143.658
R149 a_27_47.n2 a_27_47.t4 89.119
R150 a_27_47.n0 a_27_47.t2 66.666
R151 a_27_47.t3 a_27_47.n2 64.933
R152 a_27_47.n0 a_27_47.t1 28.317
R153 VNB VNB.t7 6438.23
R154 VNB.t11 VNB.t6 6292.47
R155 VNB.t4 VNB.t9 5321.88
R156 VNB.t13 VNB.t5 3947.06
R157 VNB.t10 VNB.t13 3397.06
R158 VNB.t8 VNB.t10 3138.24
R159 VNB.t5 VNB.t4 2859.74
R160 VNB.t9 VNB.t11 2717.65
R161 VNB.t7 VNB.t8 2717.65
R162 VNB.t12 VNB.t2 2586.81
R163 VNB.t1 VNB.t0 2030.77
R164 VNB.t3 VNB.t1 2030.77
R165 VNB.t2 VNB.t3 2030.77
R166 VNB.t6 VNB.t12 1740.66
R167 a_257_243.n0 a_257_243.t2 552.941
R168 a_257_243.t0 a_257_243.n1 488.627
R169 a_257_243.n1 a_257_243.t1 146.004
R170 a_257_243.n0 a_257_243.t3 121.631
R171 a_257_243.n1 a_257_243.n0 17.613
R172 VGND.n1 VGND.n0 111.956
R173 VGND.n23 VGND.n22 111.421
R174 VGND.n16 VGND.n15 106.463
R175 VGND.n34 VGND.n33 106.463
R176 VGND.n2 VGND.t0 103.713
R177 VGND.n6 VGND.n5 92.5
R178 VGND.n22 VGND.t5 65.714
R179 VGND.n22 VGND.t4 43.648
R180 VGND.n5 VGND.t2 39.692
R181 VGND.n15 VGND.t10 38.571
R182 VGND.n15 VGND.t8 38.571
R183 VGND.n33 VGND.t7 38.571
R184 VGND.n33 VGND.t6 38.571
R185 VGND.n5 VGND.t9 31.384
R186 VGND.n0 VGND.t1 24.923
R187 VGND.n0 VGND.t3 24.923
R188 VGND.n4 VGND.n3 4.65
R189 VGND.n8 VGND.n7 4.65
R190 VGND.n10 VGND.n9 4.65
R191 VGND.n12 VGND.n11 4.65
R192 VGND.n14 VGND.n13 4.65
R193 VGND.n17 VGND.n16 4.65
R194 VGND.n19 VGND.n18 4.65
R195 VGND.n21 VGND.n20 4.65
R196 VGND.n24 VGND.n23 4.65
R197 VGND.n26 VGND.n25 4.65
R198 VGND.n28 VGND.n27 4.65
R199 VGND.n30 VGND.n29 4.65
R200 VGND.n32 VGND.n31 4.65
R201 VGND.n35 VGND.n34 3.932
R202 VGND.n2 VGND.n1 3.911
R203 VGND.n7 VGND.n6 1.086
R204 VGND.n4 VGND.n2 0.23
R205 VGND.n35 VGND.n32 0.137
R206 VGND VGND.n35 0.121
R207 VGND.n8 VGND.n4 0.119
R208 VGND.n10 VGND.n8 0.119
R209 VGND.n12 VGND.n10 0.119
R210 VGND.n14 VGND.n12 0.119
R211 VGND.n17 VGND.n14 0.119
R212 VGND.n19 VGND.n17 0.119
R213 VGND.n21 VGND.n19 0.119
R214 VGND.n24 VGND.n21 0.119
R215 VGND.n26 VGND.n24 0.119
R216 VGND.n28 VGND.n26 0.119
R217 VGND.n30 VGND.n28 0.119
R218 VGND.n32 VGND.n30 0.119
R219 a_383_413.t0 a_383_413.t1 206.38
R220 a_1127_47.t0 a_1127_47.t1 38.769
R221 GATE.n0 GATE.t1 294.772
R222 GATE.n0 GATE.t0 201.586
R223 GATE GATE.n0 86.729
R224 a_395_47.t0 a_395_47.t1 138.059
C0 VGND GCLK 0.42fF
C1 VPWR VGND 0.11fF
C2 VPWR GCLK 0.55fF
C3 SCE GATE 0.11fF
C4 VPB VPWR 0.18fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__sedfxbp_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__sedfxbp_1 VPWR VGND CLK Q_N SCD DE D Q SCE VNB VPB
X0 a_2177_47.t0 a_27_47.t2 a_2051_413.t1 VNB.t6 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X1 a_381_369.t1 D.t0 a_299_47.t4 VPB.t21 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X2 a_1537_413.t1 a_27_47.t3 a_1446_413.t0 VPB.t6 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3 VPWR.t10 DE.t0 a_423_343.t1 VPB.t11 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X4 VPWR.t5 CLK.t0 a_27_47.t1 VPB.t7 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X5 VPWR.t6 SCE.t0 a_885_21.t1 VPB.t13 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X6 Q.t0 a_2051_413.t4 VGND.t3 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 VGND.t2 SCE.t1 a_885_21.t0 VNB.t13 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 Q_N.t0 a_791_264.t2 VGND.t11 VNB.t17 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 VPWR.t0 a_1610_159.t2 a_1537_413.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10 a_1610_159.t1 a_1446_413.t4 VPWR.t8 VPB.t10 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X11 a_1561_47.t1 a_193_47.t2 a_1446_413.t2 VNB.t20 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X12 VGND.t9 DE.t1 a_423_343.t0 VNB.t11 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13 a_1974_47.t0 a_1610_159.t3 VGND.t0 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14 a_915_47.t0 a_885_21.t2 a_1231_369.t0 VPB.t8 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X15 a_193_47.t0 a_27_47.t4 VGND.t5 VNB.t5 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16 a_2051_413.t2 a_193_47.t3 a_1974_47.t1 VNB.t21 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X17 a_729_47.t0 a_423_343.t2 VGND.t10 VNB.t10 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18 Q_N.t1 a_791_264.t3 VPWR.t12 VPB.t16 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X19 a_729_369.t0 DE.t2 VPWR.t9 VPB.t12 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X20 Q.t1 a_2051_413.t5 VPWR.t2 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X21 a_299_47.t2 a_791_264.t4 a_729_47.t1 VNB.t18 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22 a_1446_413.t1 a_27_47.t5 a_915_47.t4 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X23 a_2135_413.t0 a_193_47.t4 a_2051_413.t3 VPB.t19 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24 a_193_47.t1 a_27_47.t6 VPWR.t4 VPB.t5 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X25 a_1231_369.t1 SCD.t0 VPWR.t7 VPB.t15 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X26 a_915_47.t2 SCE.t2 a_1226_119.t0 VNB.t14 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X27 VPWR.t3 a_2051_413.t6 a_791_264.t1 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X28 a_2051_413.t0 a_27_47.t7 a_1960_413.t1 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X29 a_299_47.t3 a_791_264.t5 a_729_369.t1 VPB.t17 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X30 a_381_47.t1 D.t1 a_299_47.t5 VNB.t15 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X31 VPWR.t13 a_791_264.t6 a_2135_413.t1 VPB.t18 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X32 VGND.t1 a_1610_159.t4 a_1561_47.t0 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X33 VPWR.t11 a_423_343.t3 a_381_369.t0 VPB.t9 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X34 a_915_47.t3 SCE.t3 a_299_47.t1 VPB.t14 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X35 a_1960_413.t0 a_1610_159.t5 VPWR.t1 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X36 VGND.t4 a_2051_413.t7 a_791_264.t0 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X37 a_1226_119.t1 SCD.t1 VGND.t6 VNB.t16 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X38 VGND.t12 a_791_264.t7 a_2177_47.t1 VNB.t19 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X39 a_1446_413.t3 a_193_47.t5 a_915_47.t5 VPB.t20 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X40 a_915_47.t1 a_885_21.t3 a_299_47.t0 VNB.t8 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X41 VGND.t13 CLK.t1 a_27_47.t0 VNB.t7 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X42 VGND.t8 DE.t3 a_381_47.t0 VNB.t12 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X43 a_1610_159.t0 a_1446_413.t5 VGND.t7 VNB.t9 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
R0 a_27_47.n1 a_27_47.t2 443.438
R1 a_27_47.n0 a_27_47.t5 269.985
R2 a_27_47.n3 a_27_47.t6 263.405
R3 a_27_47.n1 a_27_47.t7 254.388
R4 a_27_47.t1 a_27_47.n5 244.156
R5 a_27_47.n3 a_27_47.t4 228.059
R6 a_27_47.n4 a_27_47.t0 195.871
R7 a_27_47.n0 a_27_47.t3 142.49
R8 a_27_47.n2 a_27_47.n1 113.844
R9 a_27_47.n4 a_27_47.n3 76
R10 a_27_47.n5 a_27_47.n4 35.339
R11 a_27_47.n5 a_27_47.n2 10.69
R12 a_27_47.n2 a_27_47.n0 2.9
R13 a_2051_413.n5 a_2051_413.n4 349.52
R14 a_2051_413.n0 a_2051_413.t5 212.079
R15 a_2051_413.n4 a_2051_413.n3 193.388
R16 a_2051_413.n1 a_2051_413.t7 176.733
R17 a_2051_413.n4 a_2051_413.n2 176.238
R18 a_2051_413.n2 a_2051_413.t6 163.879
R19 a_2051_413.n0 a_2051_413.t4 139.779
R20 a_2051_413.n3 a_2051_413.t1 76.666
R21 a_2051_413.n1 a_2051_413.n0 70.839
R22 a_2051_413.n5 a_2051_413.t3 63.321
R23 a_2051_413.t0 a_2051_413.n5 63.321
R24 a_2051_413.n3 a_2051_413.t2 50
R25 a_2051_413.n2 a_2051_413.n1 33.74
R26 a_2177_47.t1 a_2177_47.t0 93.059
R27 VNB.t8 VNB.t13 8836.4
R28 VNB.t12 VNB.t11 6082.35
R29 VNB.t5 VNB.t15 6082.35
R30 VNB.t17 VNB.t2 5874.73
R31 VNB.t9 VNB.t0 5346.86
R32 VNB VNB.t7 4270.59
R33 VNB.t14 VNB.t4 4015.64
R34 VNB.t21 VNB.t6 3429.41
R35 VNB.t20 VNB.t1 3429.41
R36 VNB.t10 VNB.t18 3300
R37 VNB.t0 VNB.t21 3138.24
R38 VNB.t1 VNB.t9 3130.33
R39 VNB.t6 VNB.t19 3073.53
R40 VNB.t4 VNB.t20 2847.06
R41 VNB.t11 VNB.t10 2847.06
R42 VNB.t13 VNB.t16 2717.65
R43 VNB.t18 VNB.t8 2717.65
R44 VNB.t7 VNB.t5 2717.65
R45 VNB.t2 VNB.t3 2345.05
R46 VNB.t16 VNB.t14 2329.41
R47 VNB.t15 VNB.t12 2329.41
R48 VNB.t19 VNB.t17 2303.7
R49 D.n0 D.t1 216.76
R50 D.n0 D.t0 215.106
R51 D D.n0 34.479
R52 a_299_47.n1 a_299_47.t4 321.627
R53 a_299_47.n3 a_299_47.n2 233.623
R54 a_299_47.n1 a_299_47.t5 139.932
R55 a_299_47.t1 a_299_47.n3 53.867
R56 a_299_47.n3 a_299_47.t3 41.554
R57 a_299_47.n0 a_299_47.t0 37.55
R58 a_299_47.n0 a_299_47.t2 36.873
R59 a_299_47.n2 a_299_47.n1 8.177
R60 a_299_47.n2 a_299_47.n0 8.115
R61 a_381_369.t0 a_381_369.t1 64.64
R62 VPB.t16 VPB.t2 787.227
R63 VPB.t14 VPB.t13 622.849
R64 VPB.t10 VPB.t1 556.386
R65 VPB.t9 VPB.t11 556.386
R66 VPB.t5 VPB.t21 556.386
R67 VPB.t0 VPB.t10 390.654
R68 VPB.t8 VPB.t20 383.22
R69 VPB.t13 VPB.t15 351.016
R70 VPB.t19 VPB.t18 337.383
R71 VPB.t15 VPB.t8 309.152
R72 VPB.t6 VPB.t0 304.828
R73 VPB.t12 VPB.t17 301.869
R74 VPB.t2 VPB.t3 287.071
R75 VPB.t18 VPB.t16 287.071
R76 VPB.t17 VPB.t14 272.274
R77 VPB.t1 VPB.t4 269.314
R78 VPB.t11 VPB.t12 260.436
R79 VPB.t20 VPB.t6 256.559
R80 VPB.t4 VPB.t19 248.598
R81 VPB.t7 VPB.t5 248.598
R82 VPB.t21 VPB.t9 213.084
R83 VPB VPB.t7 142.056
R84 a_1446_413.n3 a_1446_413.n2 388.236
R85 a_1446_413.n0 a_1446_413.t5 230.482
R86 a_1446_413.n0 a_1446_413.t4 196.013
R87 a_1446_413.n2 a_1446_413.n1 183.768
R88 a_1446_413.n2 a_1446_413.n0 95.938
R89 a_1446_413.t0 a_1446_413.n3 72.702
R90 a_1446_413.n3 a_1446_413.t3 70.357
R91 a_1446_413.n1 a_1446_413.t2 51.666
R92 a_1446_413.n1 a_1446_413.t1 45
R93 a_1537_413.t0 a_1537_413.t1 171.202
R94 DE.n0 DE.t2 319.725
R95 DE.n2 DE.n1 238.689
R96 DE.n0 DE.t0 178.339
R97 DE.n1 DE.n0 147.813
R98 DE.n2 DE.t3 130.384
R99 DE.n1 DE.t1 130.14
R100 DE DE.n2 82.892
R101 a_423_343.n1 a_423_343.t3 299.566
R102 a_423_343.n0 a_423_343.t2 258.036
R103 a_423_343.t1 a_423_343.n1 230.699
R104 a_423_343.n0 a_423_343.t0 151.679
R105 a_423_343.n1 a_423_343.n0 11.133
R106 VPWR.n12 VPWR.t1 375.462
R107 VPWR.n54 VPWR.n53 311.893
R108 VPWR.n30 VPWR.n29 306.598
R109 VPWR.n45 VPWR.t11 228.681
R110 VPWR.n41 VPWR.n40 176.72
R111 VPWR.n17 VPWR.n16 171.436
R112 VPWR.n1 VPWR.n0 143.182
R113 VPWR.n3 VPWR.n2 132.968
R114 VPWR.n16 VPWR.t0 106.098
R115 VPWR.n2 VPWR.t13 95.255
R116 VPWR.n0 VPWR.t3 61.912
R117 VPWR.n29 VPWR.t7 61.562
R118 VPWR.n29 VPWR.t6 60.023
R119 VPWR.n40 VPWR.t9 44.632
R120 VPWR.n40 VPWR.t10 44.632
R121 VPWR.n16 VPWR.t8 43.34
R122 VPWR.n53 VPWR.t4 41.554
R123 VPWR.n53 VPWR.t5 41.554
R124 VPWR.n0 VPWR.t2 30.241
R125 VPWR.n2 VPWR.t12 26.498
R126 VPWR.n4 VPWR.n3 13.176
R127 VPWR.n5 VPWR.n4 4.65
R128 VPWR.n7 VPWR.n6 4.65
R129 VPWR.n9 VPWR.n8 4.65
R130 VPWR.n11 VPWR.n10 4.65
R131 VPWR.n13 VPWR.n12 4.65
R132 VPWR.n15 VPWR.n14 4.65
R133 VPWR.n18 VPWR.n17 4.65
R134 VPWR.n20 VPWR.n19 4.65
R135 VPWR.n22 VPWR.n21 4.65
R136 VPWR.n24 VPWR.n23 4.65
R137 VPWR.n26 VPWR.n25 4.65
R138 VPWR.n28 VPWR.n27 4.65
R139 VPWR.n31 VPWR.n30 4.65
R140 VPWR.n33 VPWR.n32 4.65
R141 VPWR.n35 VPWR.n34 4.65
R142 VPWR.n37 VPWR.n36 4.65
R143 VPWR.n39 VPWR.n38 4.65
R144 VPWR.n42 VPWR.n41 4.65
R145 VPWR.n44 VPWR.n43 4.65
R146 VPWR.n46 VPWR.n45 4.65
R147 VPWR.n48 VPWR.n47 4.65
R148 VPWR.n50 VPWR.n49 4.65
R149 VPWR.n52 VPWR.n51 4.65
R150 VPWR.n55 VPWR.n54 3.932
R151 VPWR.n5 VPWR.n1 0.139
R152 VPWR.n55 VPWR.n52 0.137
R153 VPWR VPWR.n55 0.123
R154 VPWR.n7 VPWR.n5 0.119
R155 VPWR.n9 VPWR.n7 0.119
R156 VPWR.n11 VPWR.n9 0.119
R157 VPWR.n13 VPWR.n11 0.119
R158 VPWR.n15 VPWR.n13 0.119
R159 VPWR.n18 VPWR.n15 0.119
R160 VPWR.n20 VPWR.n18 0.119
R161 VPWR.n22 VPWR.n20 0.119
R162 VPWR.n24 VPWR.n22 0.119
R163 VPWR.n26 VPWR.n24 0.119
R164 VPWR.n28 VPWR.n26 0.119
R165 VPWR.n31 VPWR.n28 0.119
R166 VPWR.n33 VPWR.n31 0.119
R167 VPWR.n35 VPWR.n33 0.119
R168 VPWR.n37 VPWR.n35 0.119
R169 VPWR.n39 VPWR.n37 0.119
R170 VPWR.n42 VPWR.n39 0.119
R171 VPWR.n44 VPWR.n42 0.119
R172 VPWR.n46 VPWR.n44 0.119
R173 VPWR.n48 VPWR.n46 0.119
R174 VPWR.n50 VPWR.n48 0.119
R175 VPWR.n52 VPWR.n50 0.119
R176 CLK.n0 CLK.t0 292.947
R177 CLK.n0 CLK.t1 209.401
R178 CLK CLK.n0 78.067
R179 SCE.t1 SCE.t2 604.106
R180 SCE.n1 SCE.t3 352.394
R181 SCE.n0 SCE.t0 189.586
R182 SCE.n0 SCE.t1 142.029
R183 SCE SCE.n1 77.631
R184 SCE.n1 SCE.n0 74.085
R185 a_885_21.n0 a_885_21.t3 495.544
R186 a_885_21.n1 a_885_21.t2 351.552
R187 a_885_21.t1 a_885_21.n1 226.125
R188 a_885_21.n0 a_885_21.t0 131.071
R189 a_885_21.n1 a_885_21.n0 74.939
R190 VGND.n12 VGND.t0 152.016
R191 VGND.n47 VGND.t8 145.81
R192 VGND.n31 VGND.n30 130.388
R193 VGND.n43 VGND.n42 109.76
R194 VGND.n56 VGND.n55 107.239
R195 VGND.n18 VGND.n17 106.11
R196 VGND.n3 VGND.n0 74.893
R197 VGND.n17 VGND.t7 74.865
R198 VGND.n2 VGND.n1 70.639
R199 VGND.n1 VGND.t12 57.782
R200 VGND.n0 VGND.t4 57.781
R201 VGND.n42 VGND.t10 41.428
R202 VGND.n42 VGND.t9 41.428
R203 VGND.n17 VGND.t1 40
R204 VGND.n30 VGND.t6 38.571
R205 VGND.n30 VGND.t2 38.571
R206 VGND.n55 VGND.t5 38.571
R207 VGND.n55 VGND.t13 38.571
R208 VGND.n0 VGND.t3 24.78
R209 VGND.n1 VGND.t11 24.778
R210 VGND.n3 VGND.n2 10.535
R211 VGND.n5 VGND.n4 4.65
R212 VGND.n7 VGND.n6 4.65
R213 VGND.n9 VGND.n8 4.65
R214 VGND.n11 VGND.n10 4.65
R215 VGND.n14 VGND.n13 4.65
R216 VGND.n16 VGND.n15 4.65
R217 VGND.n19 VGND.n18 4.65
R218 VGND.n21 VGND.n20 4.65
R219 VGND.n23 VGND.n22 4.65
R220 VGND.n25 VGND.n24 4.65
R221 VGND.n27 VGND.n26 4.65
R222 VGND.n29 VGND.n28 4.65
R223 VGND.n33 VGND.n32 4.65
R224 VGND.n35 VGND.n34 4.65
R225 VGND.n37 VGND.n36 4.65
R226 VGND.n39 VGND.n38 4.65
R227 VGND.n41 VGND.n40 4.65
R228 VGND.n44 VGND.n43 4.65
R229 VGND.n46 VGND.n45 4.65
R230 VGND.n48 VGND.n47 4.65
R231 VGND.n50 VGND.n49 4.65
R232 VGND.n52 VGND.n51 4.65
R233 VGND.n54 VGND.n53 4.65
R234 VGND.n57 VGND.n56 3.932
R235 VGND.n13 VGND.n12 2.635
R236 VGND.n32 VGND.n31 0.752
R237 VGND.n5 VGND.n3 0.138
R238 VGND.n57 VGND.n54 0.137
R239 VGND VGND.n57 0.123
R240 VGND.n7 VGND.n5 0.119
R241 VGND.n9 VGND.n7 0.119
R242 VGND.n11 VGND.n9 0.119
R243 VGND.n14 VGND.n11 0.119
R244 VGND.n16 VGND.n14 0.119
R245 VGND.n19 VGND.n16 0.119
R246 VGND.n21 VGND.n19 0.119
R247 VGND.n23 VGND.n21 0.119
R248 VGND.n25 VGND.n23 0.119
R249 VGND.n27 VGND.n25 0.119
R250 VGND.n29 VGND.n27 0.119
R251 VGND.n33 VGND.n29 0.119
R252 VGND.n35 VGND.n33 0.119
R253 VGND.n37 VGND.n35 0.119
R254 VGND.n39 VGND.n37 0.119
R255 VGND.n41 VGND.n39 0.119
R256 VGND.n44 VGND.n41 0.119
R257 VGND.n46 VGND.n44 0.119
R258 VGND.n48 VGND.n46 0.119
R259 VGND.n50 VGND.n48 0.119
R260 VGND.n52 VGND.n50 0.119
R261 VGND.n54 VGND.n52 0.119
R262 Q Q.t1 153.46
R263 Q Q.t0 100.27
R264 a_791_264.n0 a_791_264.t6 368.968
R265 a_791_264.n3 a_791_264.t4 310.621
R266 a_791_264.t1 a_791_264.n5 248.537
R267 a_791_264.n1 a_791_264.t3 245.819
R268 a_791_264.n5 a_791_264.n2 232.442
R269 a_791_264.n3 a_791_264.t5 194.941
R270 a_791_264.n0 a_791_264.t7 189.586
R271 a_791_264.n2 a_791_264.t2 152.633
R272 a_791_264.n4 a_791_264.t0 148.576
R273 a_791_264.n4 a_791_264.n3 136.275
R274 a_791_264.n1 a_791_264.n0 96.4
R275 a_791_264.n2 a_791_264.n1 29.962
R276 a_791_264.n5 a_791_264.n4 7.717
R277 Q_N Q_N.t1 148.433
R278 Q_N Q_N.t0 102.677
R279 a_1610_159.n1 a_1610_159.t2 406.399
R280 a_1610_159.n0 a_1610_159.t5 318.12
R281 a_1610_159.t1 a_1610_159.n3 262.563
R282 a_1610_159.n0 a_1610_159.t3 194.476
R283 a_1610_159.n1 a_1610_159.t4 130.052
R284 a_1610_159.n2 a_1610_159.n1 100.533
R285 a_1610_159.n2 a_1610_159.t0 93.987
R286 a_1610_159.n3 a_1610_159.n0 92.484
R287 a_1610_159.n3 a_1610_159.n2 9.323
R288 a_193_47.n1 a_193_47.t2 389.542
R289 a_193_47.n1 a_193_47.t5 273.571
R290 a_193_47.t1 a_193_47.n3 249.337
R291 a_193_47.n0 a_193_47.t4 232.651
R292 a_193_47.n0 a_193_47.t3 222.372
R293 a_193_47.n3 a_193_47.t0 207.871
R294 a_193_47.n2 a_193_47.n1 93.104
R295 a_193_47.n3 a_193_47.n2 9.98
R296 a_193_47.n2 a_193_47.n0 7.6
R297 a_1561_47.t0 a_1561_47.t1 111.393
R298 a_1974_47.n0 a_1974_47.t1 70
R299 a_1974_47.n0 a_1974_47.t0 26.393
R300 a_1974_47.n1 a_1974_47.n0 14.4
R301 a_1231_369.t0 a_1231_369.t1 101.578
R302 a_915_47.n0 a_915_47.t3 305.928
R303 a_915_47.n5 a_915_47.n4 221.84
R304 a_915_47.n5 a_915_47.t5 117.17
R305 a_915_47.n2 a_915_47.n1 97.479
R306 a_915_47.n4 a_915_47.n3 92.5
R307 a_915_47.n1 a_915_47.t4 75.384
R308 a_915_47.t0 a_915_47.n5 61.587
R309 a_915_47.n0 a_915_47.t1 46.679
R310 a_915_47.n3 a_915_47.t2 32.197
R311 a_915_47.n4 a_915_47.n2 9.521
R312 a_915_47.n2 a_915_47.n0 7.415
R313 a_729_47.t0 a_729_47.t1 102.857
R314 a_729_369.t0 a_729_369.t1 110.812
R315 a_2135_413.t0 a_2135_413.t1 197
R316 SCD.n0 SCD.t1 206.188
R317 SCD.n0 SCD.t0 183.694
R318 SCD SCD.n0 87.674
R319 a_1226_119.t0 a_1226_119.t1 60
R320 a_1960_413.t0 a_1960_413.t1 143.059
R321 a_381_47.t0 a_381_47.t1 60
C0 VGND Q 0.17fF
C1 VPWR VGND 0.15fF
C2 VPB VGND 0.10fF
C3 VPWR Q_N 0.16fF
C4 D DE 0.13fF
C5 VGND Q_N 0.17fF
C6 VPWR Q 0.21fF
C7 VPB VPWR 0.30fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__sedfxbp_2.ext - technology: sky130A

.subckt sky130_fd_sc_hd__sedfxbp_2 VPWR VGND CLK Q_N SCD DE D Q SCE VNB VPB
X0 a_2177_47.t1 a_27_47.t2 a_2051_413.t1 VNB.t11 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X1 VGND.t7 a_791_264.t2 Q_N.t1 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 a_381_369.t0 D.t0 a_299_47.t1 VPB.t5 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X3 a_1537_413.t1 a_27_47.t3 a_1446_413.t1 VPB.t8 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 VGND.t2 a_2051_413.t4 a_791_264.t0 VNB.t8 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 VPWR.t5 DE.t0 a_423_343.t0 VPB.t18 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X6 VPWR.t14 CLK.t0 a_27_47.t0 VPB.t19 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X7 VPWR.t13 SCE.t0 a_885_21.t0 VPB.t16 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X8 VGND.t10 SCE.t1 a_885_21.t1 VNB.t14 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9 VGND.t4 a_2051_413.t5 Q.t3 VNB.t7 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 Q_N.t0 a_791_264.t3 VGND.t6 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 VPWR.t0 a_1610_159.t2 a_1537_413.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12 a_1610_159.t0 a_1446_413.t4 VPWR.t11 VPB.t21 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X13 a_1561_47.t0 a_193_47.t2 a_1446_413.t2 VNB.t22 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X14 VGND.t14 DE.t1 a_423_343.t1 VNB.t20 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15 a_1974_47.t1 a_1610_159.t3 VGND.t0 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16 VPWR.t9 a_791_264.t4 Q_N.t3 VPB.t12 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17 VPWR.t4 a_2051_413.t6 Q.t1 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X18 a_915_47.t5 a_885_21.t2 a_1231_369.t1 VPB.t14 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X19 a_193_47.t1 a_27_47.t4 VGND.t5 VNB.t10 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20 a_2051_413.t2 a_193_47.t3 a_1974_47.t0 VNB.t23 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X21 a_729_47.t1 a_423_343.t2 VGND.t12 VNB.t17 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22 Q.t0 a_2051_413.t7 VPWR.t3 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X23 Q_N.t2 a_791_264.t5 VPWR.t8 VPB.t11 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X24 a_729_369.t0 DE.t2 VPWR.t6 VPB.t15 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X25 VPWR.t2 a_2051_413.t8 a_791_264.t1 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X26 a_299_47.t2 a_791_264.t6 a_729_47.t0 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X27 a_1446_413.t0 a_27_47.t5 a_915_47.t0 VNB.t9 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X28 a_2135_413.t1 a_193_47.t4 a_2051_413.t3 VPB.t22 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X29 a_193_47.t0 a_27_47.t6 VPWR.t7 VPB.t7 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X30 a_1231_369.t0 SCD.t0 VPWR.t12 VPB.t13 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X31 a_915_47.t2 SCE.t2 a_1226_119.t0 VNB.t15 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X32 a_2051_413.t0 a_27_47.t7 a_1960_413.t0 VPB.t6 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X33 a_299_47.t3 a_791_264.t7 a_729_369.t1 VPB.t10 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X34 a_381_47.t0 D.t1 a_299_47.t0 VNB.t19 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X35 VPWR.t10 a_791_264.t8 a_2135_413.t0 VPB.t9 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X36 VGND.t1 a_1610_159.t4 a_1561_47.t1 VNB.t5 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X37 VPWR.t15 a_423_343.t3 a_381_369.t1 VPB.t20 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X38 a_915_47.t3 SCE.t3 a_299_47.t5 VPB.t17 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X39 a_1960_413.t1 a_1610_159.t5 VPWR.t1 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X40 a_1226_119.t1 SCD.t1 VGND.t9 VNB.t12 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X41 VGND.t8 a_791_264.t9 a_2177_47.t0 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X42 a_1446_413.t3 a_193_47.t5 a_915_47.t1 VPB.t23 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X43 a_915_47.t4 a_885_21.t3 a_299_47.t4 VNB.t13 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X44 VGND.t11 CLK.t1 a_27_47.t1 VNB.t16 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X45 VGND.t13 DE.t3 a_381_47.t1 VNB.t18 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X46 a_1610_159.t1 a_1446_413.t5 VGND.t15 VNB.t21 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X47 Q.t2 a_2051_413.t9 VGND.t3 VNB.t6 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
R0 a_27_47.n1 a_27_47.t2 443.438
R1 a_27_47.n0 a_27_47.t5 269.985
R2 a_27_47.n3 a_27_47.t6 263.405
R3 a_27_47.n1 a_27_47.t7 254.388
R4 a_27_47.t0 a_27_47.n5 244.156
R5 a_27_47.n3 a_27_47.t4 228.059
R6 a_27_47.n4 a_27_47.t1 195.871
R7 a_27_47.n0 a_27_47.t3 142.49
R8 a_27_47.n2 a_27_47.n1 113.844
R9 a_27_47.n4 a_27_47.n3 76
R10 a_27_47.n5 a_27_47.n4 35.339
R11 a_27_47.n5 a_27_47.n2 10.69
R12 a_27_47.n2 a_27_47.n0 2.9
R13 a_2051_413.n6 a_2051_413.n5 349.52
R14 a_2051_413.n0 a_2051_413.t6 212.079
R15 a_2051_413.n1 a_2051_413.t7 212.079
R16 a_2051_413.n5 a_2051_413.n4 193.388
R17 a_2051_413.n2 a_2051_413.t4 176.733
R18 a_2051_413.n5 a_2051_413.n3 176.613
R19 a_2051_413.n3 a_2051_413.t8 163.879
R20 a_2051_413.n0 a_2051_413.t5 139.779
R21 a_2051_413.n1 a_2051_413.t9 139.779
R22 a_2051_413.n4 a_2051_413.t1 76.666
R23 a_2051_413.n2 a_2051_413.n1 70.839
R24 a_2051_413.n6 a_2051_413.t3 63.321
R25 a_2051_413.t0 a_2051_413.n6 63.321
R26 a_2051_413.n1 a_2051_413.n0 61.345
R27 a_2051_413.n4 a_2051_413.t2 50
R28 a_2051_413.n3 a_2051_413.n2 33.74
R29 a_2177_47.t0 a_2177_47.t1 93.059
R30 VNB.t13 VNB.t14 8836.4
R31 VNB.t18 VNB.t20 6082.35
R32 VNB.t10 VNB.t19 6082.35
R33 VNB.t1 VNB.t8 5874.73
R34 VNB.t21 VNB.t4 5346.86
R35 VNB VNB.t16 4270.59
R36 VNB.t15 VNB.t9 4015.64
R37 VNB.t23 VNB.t11 3429.41
R38 VNB.t22 VNB.t5 3429.41
R39 VNB.t17 VNB.t3 3300
R40 VNB.t4 VNB.t23 3138.24
R41 VNB.t5 VNB.t21 3130.33
R42 VNB.t11 VNB.t0 3073.53
R43 VNB.t9 VNB.t22 2847.06
R44 VNB.t20 VNB.t17 2847.06
R45 VNB.t14 VNB.t12 2717.65
R46 VNB.t3 VNB.t13 2717.65
R47 VNB.t16 VNB.t10 2717.65
R48 VNB.t8 VNB.t6 2345.05
R49 VNB.t12 VNB.t15 2329.41
R50 VNB.t19 VNB.t18 2329.41
R51 VNB.t0 VNB.t2 2303.7
R52 VNB.t6 VNB.t7 2030.77
R53 VNB.t2 VNB.t1 2030.77
R54 a_791_264.n0 a_791_264.t8 368.968
R55 a_791_264.n5 a_791_264.t6 310.621
R56 a_791_264.t1 a_791_264.n7 248.537
R57 a_791_264.n3 a_791_264.t4 245.819
R58 a_791_264.n1 a_791_264.t5 245.819
R59 a_791_264.n7 a_791_264.n4 232.442
R60 a_791_264.n5 a_791_264.t7 194.941
R61 a_791_264.n0 a_791_264.t9 189.586
R62 a_791_264.n2 a_791_264.t3 152.633
R63 a_791_264.n4 a_791_264.t2 152.633
R64 a_791_264.n6 a_791_264.t0 148.576
R65 a_791_264.n6 a_791_264.n5 136.65
R66 a_791_264.n1 a_791_264.n0 96.4
R67 a_791_264.n3 a_791_264.n2 79.464
R68 a_791_264.n4 a_791_264.n3 29.962
R69 a_791_264.n2 a_791_264.n1 29.962
R70 a_791_264.n7 a_791_264.n6 7.717
R71 Q_N Q_N.n0 122.94
R72 Q_N Q_N.n1 63.278
R73 Q_N.n0 Q_N.t3 26.595
R74 Q_N.n0 Q_N.t2 26.595
R75 Q_N.n1 Q_N.t1 24.923
R76 Q_N.n1 Q_N.t0 24.923
R77 VGND.n22 VGND.t0 152.016
R78 VGND.n57 VGND.t13 145.81
R79 VGND.n41 VGND.n40 130.388
R80 VGND.n53 VGND.n52 109.76
R81 VGND.n5 VGND.t7 109.721
R82 VGND.n2 VGND.t4 109.607
R83 VGND.n66 VGND.n65 107.239
R84 VGND.n28 VGND.n27 106.11
R85 VGND.n27 VGND.t15 74.865
R86 VGND.n1 VGND.n0 72.154
R87 VGND.n11 VGND.n10 70.639
R88 VGND.n10 VGND.t8 57.782
R89 VGND.n0 VGND.t2 57.779
R90 VGND.n52 VGND.t12 41.428
R91 VGND.n52 VGND.t14 41.428
R92 VGND.n27 VGND.t1 40
R93 VGND.n40 VGND.t9 38.571
R94 VGND.n40 VGND.t10 38.571
R95 VGND.n65 VGND.t5 38.571
R96 VGND.n65 VGND.t11 38.571
R97 VGND.n0 VGND.t3 24.782
R98 VGND.n10 VGND.t6 24.778
R99 VGND.n6 VGND.n5 6.4
R100 VGND.n12 VGND.n11 6.4
R101 VGND.n4 VGND.n3 4.65
R102 VGND.n7 VGND.n6 4.65
R103 VGND.n9 VGND.n8 4.65
R104 VGND.n13 VGND.n12 4.65
R105 VGND.n15 VGND.n14 4.65
R106 VGND.n17 VGND.n16 4.65
R107 VGND.n19 VGND.n18 4.65
R108 VGND.n21 VGND.n20 4.65
R109 VGND.n24 VGND.n23 4.65
R110 VGND.n26 VGND.n25 4.65
R111 VGND.n29 VGND.n28 4.65
R112 VGND.n31 VGND.n30 4.65
R113 VGND.n33 VGND.n32 4.65
R114 VGND.n35 VGND.n34 4.65
R115 VGND.n37 VGND.n36 4.65
R116 VGND.n39 VGND.n38 4.65
R117 VGND.n43 VGND.n42 4.65
R118 VGND.n45 VGND.n44 4.65
R119 VGND.n47 VGND.n46 4.65
R120 VGND.n49 VGND.n48 4.65
R121 VGND.n51 VGND.n50 4.65
R122 VGND.n54 VGND.n53 4.65
R123 VGND.n56 VGND.n55 4.65
R124 VGND.n58 VGND.n57 4.65
R125 VGND.n60 VGND.n59 4.65
R126 VGND.n62 VGND.n61 4.65
R127 VGND.n64 VGND.n63 4.65
R128 VGND.n67 VGND.n66 3.932
R129 VGND.n2 VGND.n1 3.804
R130 VGND.n23 VGND.n22 2.635
R131 VGND.n42 VGND.n41 0.752
R132 VGND.n4 VGND.n2 0.216
R133 VGND.n67 VGND.n64 0.137
R134 VGND VGND.n67 0.123
R135 VGND.n7 VGND.n4 0.119
R136 VGND.n9 VGND.n7 0.119
R137 VGND.n13 VGND.n9 0.119
R138 VGND.n15 VGND.n13 0.119
R139 VGND.n17 VGND.n15 0.119
R140 VGND.n19 VGND.n17 0.119
R141 VGND.n21 VGND.n19 0.119
R142 VGND.n24 VGND.n21 0.119
R143 VGND.n26 VGND.n24 0.119
R144 VGND.n29 VGND.n26 0.119
R145 VGND.n31 VGND.n29 0.119
R146 VGND.n33 VGND.n31 0.119
R147 VGND.n35 VGND.n33 0.119
R148 VGND.n37 VGND.n35 0.119
R149 VGND.n39 VGND.n37 0.119
R150 VGND.n43 VGND.n39 0.119
R151 VGND.n45 VGND.n43 0.119
R152 VGND.n47 VGND.n45 0.119
R153 VGND.n49 VGND.n47 0.119
R154 VGND.n51 VGND.n49 0.119
R155 VGND.n54 VGND.n51 0.119
R156 VGND.n56 VGND.n54 0.119
R157 VGND.n58 VGND.n56 0.119
R158 VGND.n60 VGND.n58 0.119
R159 VGND.n62 VGND.n60 0.119
R160 VGND.n64 VGND.n62 0.119
R161 D.n0 D.t1 216.76
R162 D.n0 D.t0 215.106
R163 D D.n0 34.479
R164 a_299_47.t1 a_299_47.n3 321.627
R165 a_299_47.n2 a_299_47.n0 233.622
R166 a_299_47.n3 a_299_47.t0 139.932
R167 a_299_47.n0 a_299_47.t5 53.867
R168 a_299_47.n0 a_299_47.t3 41.554
R169 a_299_47.n1 a_299_47.t4 37.55
R170 a_299_47.n1 a_299_47.t2 36.873
R171 a_299_47.n3 a_299_47.n2 8.177
R172 a_299_47.n2 a_299_47.n1 8.115
R173 a_381_369.t0 a_381_369.t1 64.64
R174 VPB.t12 VPB.t2 787.227
R175 VPB.t17 VPB.t16 622.849
R176 VPB.t21 VPB.t1 556.386
R177 VPB.t20 VPB.t18 556.386
R178 VPB.t7 VPB.t5 556.386
R179 VPB.t0 VPB.t21 390.654
R180 VPB.t14 VPB.t23 383.22
R181 VPB.t16 VPB.t13 351.016
R182 VPB.t22 VPB.t9 337.383
R183 VPB.t13 VPB.t14 309.152
R184 VPB.t8 VPB.t0 304.828
R185 VPB.t15 VPB.t10 301.869
R186 VPB.t2 VPB.t3 287.071
R187 VPB.t9 VPB.t11 287.071
R188 VPB.t10 VPB.t17 272.274
R189 VPB.t1 VPB.t6 269.314
R190 VPB.t18 VPB.t15 260.436
R191 VPB.t23 VPB.t8 256.559
R192 VPB.t3 VPB.t4 248.598
R193 VPB.t11 VPB.t12 248.598
R194 VPB.t6 VPB.t22 248.598
R195 VPB.t19 VPB.t7 248.598
R196 VPB.t5 VPB.t20 213.084
R197 VPB VPB.t19 142.056
R198 a_1446_413.n3 a_1446_413.n2 388.236
R199 a_1446_413.n0 a_1446_413.t5 230.482
R200 a_1446_413.n0 a_1446_413.t4 196.013
R201 a_1446_413.n2 a_1446_413.n1 183.768
R202 a_1446_413.n2 a_1446_413.n0 95.938
R203 a_1446_413.t1 a_1446_413.n3 72.702
R204 a_1446_413.n3 a_1446_413.t3 70.357
R205 a_1446_413.n1 a_1446_413.t2 51.666
R206 a_1446_413.n1 a_1446_413.t0 45
R207 a_1537_413.t0 a_1537_413.t1 171.202
R208 DE.n0 DE.t2 319.725
R209 DE.n2 DE.n1 238.689
R210 DE.n0 DE.t0 178.339
R211 DE.n1 DE.n0 147.813
R212 DE.n2 DE.t3 130.384
R213 DE.n1 DE.t1 130.14
R214 DE DE.n2 82.892
R215 a_423_343.n1 a_423_343.t3 299.566
R216 a_423_343.n0 a_423_343.t2 258.036
R217 a_423_343.t0 a_423_343.n1 230.699
R218 a_423_343.n0 a_423_343.t1 151.679
R219 a_423_343.n1 a_423_343.n0 11.133
R220 VPWR.n22 VPWR.t1 375.462
R221 VPWR.n64 VPWR.n63 311.893
R222 VPWR.n40 VPWR.n39 306.598
R223 VPWR.n55 VPWR.t15 228.681
R224 VPWR.n51 VPWR.n50 176.72
R225 VPWR.n27 VPWR.n26 171.436
R226 VPWR.n2 VPWR.t4 158.694
R227 VPWR.n7 VPWR.t9 154.252
R228 VPWR.n1 VPWR.n0 140.629
R229 VPWR.n13 VPWR.n12 132.968
R230 VPWR.n26 VPWR.t0 106.098
R231 VPWR.n12 VPWR.t10 95.255
R232 VPWR.n0 VPWR.t2 61.911
R233 VPWR.n39 VPWR.t12 61.562
R234 VPWR.n39 VPWR.t13 60.023
R235 VPWR.n50 VPWR.t6 44.632
R236 VPWR.n50 VPWR.t5 44.632
R237 VPWR.n26 VPWR.t11 43.34
R238 VPWR.n63 VPWR.t7 41.554
R239 VPWR.n63 VPWR.t14 41.554
R240 VPWR.n0 VPWR.t3 30.242
R241 VPWR.n12 VPWR.t8 26.498
R242 VPWR.n14 VPWR.n13 13.176
R243 VPWR.n4 VPWR.n3 4.65
R244 VPWR.n6 VPWR.n5 4.65
R245 VPWR.n9 VPWR.n8 4.65
R246 VPWR.n11 VPWR.n10 4.65
R247 VPWR.n15 VPWR.n14 4.65
R248 VPWR.n17 VPWR.n16 4.65
R249 VPWR.n19 VPWR.n18 4.65
R250 VPWR.n21 VPWR.n20 4.65
R251 VPWR.n23 VPWR.n22 4.65
R252 VPWR.n25 VPWR.n24 4.65
R253 VPWR.n28 VPWR.n27 4.65
R254 VPWR.n30 VPWR.n29 4.65
R255 VPWR.n32 VPWR.n31 4.65
R256 VPWR.n34 VPWR.n33 4.65
R257 VPWR.n36 VPWR.n35 4.65
R258 VPWR.n38 VPWR.n37 4.65
R259 VPWR.n41 VPWR.n40 4.65
R260 VPWR.n43 VPWR.n42 4.65
R261 VPWR.n45 VPWR.n44 4.65
R262 VPWR.n47 VPWR.n46 4.65
R263 VPWR.n49 VPWR.n48 4.65
R264 VPWR.n52 VPWR.n51 4.65
R265 VPWR.n54 VPWR.n53 4.65
R266 VPWR.n56 VPWR.n55 4.65
R267 VPWR.n58 VPWR.n57 4.65
R268 VPWR.n60 VPWR.n59 4.65
R269 VPWR.n62 VPWR.n61 4.65
R270 VPWR.n65 VPWR.n64 3.932
R271 VPWR.n2 VPWR.n1 3.804
R272 VPWR.n8 VPWR.n7 0.752
R273 VPWR.n4 VPWR.n2 0.216
R274 VPWR.n65 VPWR.n62 0.137
R275 VPWR VPWR.n65 0.123
R276 VPWR.n6 VPWR.n4 0.119
R277 VPWR.n9 VPWR.n6 0.119
R278 VPWR.n11 VPWR.n9 0.119
R279 VPWR.n15 VPWR.n11 0.119
R280 VPWR.n17 VPWR.n15 0.119
R281 VPWR.n19 VPWR.n17 0.119
R282 VPWR.n21 VPWR.n19 0.119
R283 VPWR.n23 VPWR.n21 0.119
R284 VPWR.n25 VPWR.n23 0.119
R285 VPWR.n28 VPWR.n25 0.119
R286 VPWR.n30 VPWR.n28 0.119
R287 VPWR.n32 VPWR.n30 0.119
R288 VPWR.n34 VPWR.n32 0.119
R289 VPWR.n36 VPWR.n34 0.119
R290 VPWR.n38 VPWR.n36 0.119
R291 VPWR.n41 VPWR.n38 0.119
R292 VPWR.n43 VPWR.n41 0.119
R293 VPWR.n45 VPWR.n43 0.119
R294 VPWR.n47 VPWR.n45 0.119
R295 VPWR.n49 VPWR.n47 0.119
R296 VPWR.n52 VPWR.n49 0.119
R297 VPWR.n54 VPWR.n52 0.119
R298 VPWR.n56 VPWR.n54 0.119
R299 VPWR.n58 VPWR.n56 0.119
R300 VPWR.n60 VPWR.n58 0.119
R301 VPWR.n62 VPWR.n60 0.119
R302 CLK.n0 CLK.t0 292.947
R303 CLK.n0 CLK.t1 209.401
R304 CLK CLK.n0 78.067
R305 SCE.t1 SCE.t2 604.106
R306 SCE.n1 SCE.t3 352.394
R307 SCE.n0 SCE.t0 189.586
R308 SCE.n0 SCE.t1 142.029
R309 SCE SCE.n1 77.631
R310 SCE.n1 SCE.n0 74.085
R311 a_885_21.n0 a_885_21.t3 495.544
R312 a_885_21.n1 a_885_21.t2 351.552
R313 a_885_21.t0 a_885_21.n1 226.125
R314 a_885_21.n0 a_885_21.t1 131.071
R315 a_885_21.n1 a_885_21.n0 74.939
R316 Q Q.n0 124.895
R317 Q Q.n1 63.679
R318 Q.n0 Q.t1 26.595
R319 Q.n0 Q.t0 26.595
R320 Q.n1 Q.t3 24.923
R321 Q.n1 Q.t2 24.923
R322 a_1610_159.n1 a_1610_159.t2 406.399
R323 a_1610_159.n0 a_1610_159.t5 318.12
R324 a_1610_159.t0 a_1610_159.n3 262.563
R325 a_1610_159.n0 a_1610_159.t3 194.476
R326 a_1610_159.n1 a_1610_159.t4 130.052
R327 a_1610_159.n2 a_1610_159.n1 100.533
R328 a_1610_159.n2 a_1610_159.t1 93.987
R329 a_1610_159.n3 a_1610_159.n0 92.484
R330 a_1610_159.n3 a_1610_159.n2 9.323
R331 a_193_47.n1 a_193_47.t2 389.542
R332 a_193_47.n1 a_193_47.t5 273.571
R333 a_193_47.t0 a_193_47.n3 249.337
R334 a_193_47.n0 a_193_47.t4 232.651
R335 a_193_47.n0 a_193_47.t3 222.372
R336 a_193_47.n3 a_193_47.t1 207.871
R337 a_193_47.n2 a_193_47.n1 93.104
R338 a_193_47.n3 a_193_47.n2 9.98
R339 a_193_47.n2 a_193_47.n0 7.6
R340 a_1561_47.t1 a_1561_47.t0 111.393
R341 a_1974_47.n0 a_1974_47.t0 70
R342 a_1974_47.n0 a_1974_47.t1 26.393
R343 a_1974_47.n1 a_1974_47.n0 14.4
R344 a_1231_369.t0 a_1231_369.t1 101.578
R345 a_915_47.t3 a_915_47.n5 305.929
R346 a_915_47.n2 a_915_47.n0 221.84
R347 a_915_47.n0 a_915_47.t1 117.17
R348 a_915_47.n4 a_915_47.n3 97.479
R349 a_915_47.n2 a_915_47.n1 92.5
R350 a_915_47.n3 a_915_47.t0 75.384
R351 a_915_47.n0 a_915_47.t5 61.587
R352 a_915_47.n5 a_915_47.t4 46.68
R353 a_915_47.n1 a_915_47.t2 32.197
R354 a_915_47.n4 a_915_47.n2 9.521
R355 a_915_47.n5 a_915_47.n4 7.415
R356 a_729_47.t0 a_729_47.t1 102.857
R357 a_729_369.t0 a_729_369.t1 110.812
R358 a_2135_413.t0 a_2135_413.t1 197
R359 SCD.n0 SCD.t1 206.188
R360 SCD.n0 SCD.t0 183.694
R361 SCD SCD.n0 87.674
R362 a_1226_119.t0 a_1226_119.t1 60
R363 a_1960_413.t0 a_1960_413.t1 143.059
R364 a_381_47.t0 a_381_47.t1 60
C0 D DE 0.13fF
C1 VPWR Q 0.36fF
C2 VGND Q_N 0.28fF
C3 VPB VPWR 0.33fF
C4 VGND Q 0.27fF
C5 VPWR VGND 0.19fF
C6 VPB VGND 0.11fF
C7 VPWR Q_N 0.33fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__sedfxtp_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__sedfxtp_1 VPWR VGND CLK SCD DE D Q SCE VNB VPB
X0 a_2177_47.t1 a_27_47.t2 a_2051_413.t3 VNB.t14 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X1 a_381_369.t1 D.t0 a_299_47.t3 VPB.t14 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X2 a_1537_413.t1 a_27_47.t3 a_1446_413.t3 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3 VPWR.t4 DE.t0 a_423_343.t1 VPB.t5 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X4 VPWR.t6 CLK.t0 a_27_47.t1 VPB.t7 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X5 VPWR.t7 SCE.t0 a_885_21.t1 VPB.t8 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X6 VGND.t6 SCE.t1 a_885_21.t0 VNB.t9 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7 VPWR.t0 a_1610_159.t2 a_1537_413.t0 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 a_1610_159.t1 a_1446_413.t4 VPWR.t2 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X9 a_1561_47.t0 a_193_47.t2 a_1446_413.t0 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X10 VGND.t9 a_2051_413.t4 a_791_264.t0 VNB.t16 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11 VGND.t3 DE.t1 a_423_343.t0 VNB.t7 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12 a_1974_47.t1 a_1610_159.t3 VGND.t11 VNB.t17 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13 a_915_47.t0 a_885_21.t2 a_1231_369.t0 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X14 a_193_47.t0 a_27_47.t4 VGND.t8 VNB.t13 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15 a_2051_413.t0 a_193_47.t3 a_1974_47.t0 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X16 a_729_47.t0 a_423_343.t2 VGND.t4 VNB.t20 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17 a_729_369.t0 DE.t2 VPWR.t3 VPB.t6 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X18 Q.t0 a_2051_413.t5 VGND.t10 VNB.t15 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X19 a_299_47.t0 a_791_264.t2 a_729_47.t1 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20 a_1446_413.t2 a_27_47.t5 a_915_47.t5 VNB.t12 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X21 a_2135_413.t0 a_193_47.t4 a_2051_413.t1 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22 a_193_47.t1 a_27_47.t6 VPWR.t9 VPB.t11 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X23 a_1231_369.t1 SCD.t0 VPWR.t8 VPB.t10 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X24 a_915_47.t3 SCE.t2 a_1226_119.t0 VNB.t8 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X25 a_2051_413.t2 a_27_47.t7 a_1960_413.t0 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X26 a_299_47.t1 a_791_264.t3 a_729_369.t1 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X27 a_381_47.t1 D.t1 a_299_47.t4 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X28 VPWR.t1 a_791_264.t4 a_2135_413.t1 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X29 VGND.t12 a_1610_159.t4 a_1561_47.t1 VNB.t18 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X30 Q.t1 a_2051_413.t6 VPWR.t10 VPB.t13 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X31 VPWR.t5 a_423_343.t3 a_381_369.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X32 a_915_47.t4 SCE.t3 a_299_47.t2 VPB.t9 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X33 a_1960_413.t1 a_1610_159.t5 VPWR.t12 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X34 a_1226_119.t1 SCD.t1 VGND.t5 VNB.t5 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X35 VGND.t7 a_791_264.t5 a_2177_47.t0 VNB.t11 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X36 a_1446_413.t1 a_193_47.t5 a_915_47.t2 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X37 a_915_47.t1 a_885_21.t3 a_299_47.t5 VNB.t19 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X38 VPWR.t11 a_2051_413.t7 a_791_264.t1 VPB.t12 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X39 VGND.t0 CLK.t1 a_27_47.t0 VNB.t6 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X40 VGND.t2 DE.t3 a_381_47.t0 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X41 a_1610_159.t0 a_1446_413.t5 VGND.t1 VNB.t10 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
R0 a_27_47.n1 a_27_47.t2 443.438
R1 a_27_47.n0 a_27_47.t5 269.985
R2 a_27_47.n3 a_27_47.t6 263.405
R3 a_27_47.n1 a_27_47.t7 254.388
R4 a_27_47.t1 a_27_47.n5 244.156
R5 a_27_47.n3 a_27_47.t4 228.059
R6 a_27_47.n4 a_27_47.t0 195.871
R7 a_27_47.n0 a_27_47.t3 142.49
R8 a_27_47.n2 a_27_47.n1 113.844
R9 a_27_47.n4 a_27_47.n3 76
R10 a_27_47.n5 a_27_47.n4 35.339
R11 a_27_47.n5 a_27_47.n2 10.69
R12 a_27_47.n2 a_27_47.n0 2.9
R13 a_2051_413.n4 a_2051_413.n3 398.525
R14 a_2051_413.n2 a_2051_413.t7 269.919
R15 a_2051_413.n1 a_2051_413.t6 212.079
R16 a_2051_413.n2 a_2051_413.t4 176.733
R17 a_2051_413.n3 a_2051_413.n2 176.181
R18 a_2051_413.n3 a_2051_413.n0 159.603
R19 a_2051_413.n1 a_2051_413.t5 139.779
R20 a_2051_413.n0 a_2051_413.t3 76.666
R21 a_2051_413.n2 a_2051_413.n1 70.839
R22 a_2051_413.t1 a_2051_413.n4 63.321
R23 a_2051_413.n4 a_2051_413.t2 63.321
R24 a_2051_413.n0 a_2051_413.t0 50
R25 a_2177_47.t0 a_2177_47.t1 93.059
R26 VNB.t19 VNB.t9 8836.4
R27 VNB.t11 VNB.t16 6082.35
R28 VNB.t4 VNB.t7 6082.35
R29 VNB.t13 VNB.t3 6082.35
R30 VNB.t10 VNB.t17 5346.86
R31 VNB VNB.t6 4270.59
R32 VNB.t8 VNB.t12 4015.64
R33 VNB.t1 VNB.t14 3429.41
R34 VNB.t0 VNB.t18 3429.41
R35 VNB.t20 VNB.t2 3300
R36 VNB.t17 VNB.t1 3138.24
R37 VNB.t18 VNB.t10 3130.33
R38 VNB.t14 VNB.t11 3073.53
R39 VNB.t12 VNB.t0 2847.06
R40 VNB.t7 VNB.t20 2847.06
R41 VNB.t9 VNB.t5 2717.65
R42 VNB.t2 VNB.t19 2717.65
R43 VNB.t6 VNB.t13 2717.65
R44 VNB.t5 VNB.t8 2329.41
R45 VNB.t3 VNB.t4 2329.41
R46 VNB.t16 VNB.t15 2303.7
R47 D.n0 D.t1 216.76
R48 D.n0 D.t0 215.106
R49 D D.n0 34.479
R50 a_299_47.n1 a_299_47.t3 321.627
R51 a_299_47.n3 a_299_47.n2 233.623
R52 a_299_47.n1 a_299_47.t4 139.932
R53 a_299_47.n3 a_299_47.t2 53.867
R54 a_299_47.t1 a_299_47.n3 41.554
R55 a_299_47.n0 a_299_47.t5 37.55
R56 a_299_47.n0 a_299_47.t0 36.873
R57 a_299_47.n2 a_299_47.n1 8.177
R58 a_299_47.n2 a_299_47.n0 8.115
R59 a_381_369.t0 a_381_369.t1 64.64
R60 VPB.t9 VPB.t8 622.849
R61 VPB.t0 VPB.t5 556.386
R62 VPB.t11 VPB.t14 556.386
R63 VPB.t1 VPB.t2 383.22
R64 VPB.t8 VPB.t10 351.016
R65 VPB.t10 VPB.t1 309.152
R66 VPB.t6 VPB.t4 301.869
R67 VPB.t4 VPB.t9 272.274
R68 VPB.t5 VPB.t6 260.436
R69 VPB.t7 VPB.t11 248.598
R70 VPB.t14 VPB.t0 213.084
R71 VPB VPB.t7 142.056
R72 VPB.t3 VPB.t13 18.759
R73 VPB.t2 VPB.t12 10.958
R74 VPB.t12 VPB.t3 8.254
R75 a_1446_413.n3 a_1446_413.n2 388.236
R76 a_1446_413.n0 a_1446_413.t5 230.482
R77 a_1446_413.n0 a_1446_413.t4 196.013
R78 a_1446_413.n2 a_1446_413.n1 183.768
R79 a_1446_413.n2 a_1446_413.n0 95.938
R80 a_1446_413.n3 a_1446_413.t3 72.702
R81 a_1446_413.t1 a_1446_413.n3 70.357
R82 a_1446_413.n1 a_1446_413.t0 51.666
R83 a_1446_413.n1 a_1446_413.t2 45
R84 a_1537_413.t0 a_1537_413.t1 171.202
R85 DE.n0 DE.t2 319.725
R86 DE.n2 DE.n1 238.689
R87 DE.n0 DE.t0 178.339
R88 DE.n1 DE.n0 147.813
R89 DE.n2 DE.t3 130.384
R90 DE.n1 DE.t1 130.14
R91 DE DE.n2 82.892
R92 a_423_343.n1 a_423_343.t3 299.566
R93 a_423_343.n0 a_423_343.t2 258.036
R94 a_423_343.t1 a_423_343.n1 230.699
R95 a_423_343.n0 a_423_343.t0 151.679
R96 a_423_343.n1 a_423_343.n0 11.133
R97 VPWR.n2 VPWR.t1 378.842
R98 VPWR.n11 VPWR.t12 375.462
R99 VPWR.n53 VPWR.n52 311.893
R100 VPWR.n29 VPWR.n28 306.598
R101 VPWR.n44 VPWR.t5 228.681
R102 VPWR.n40 VPWR.n39 176.72
R103 VPWR.n16 VPWR.n15 171.436
R104 VPWR.n1 VPWR.n0 144.883
R105 VPWR.n15 VPWR.t0 106.098
R106 VPWR.n0 VPWR.t11 61.912
R107 VPWR.n28 VPWR.t8 61.562
R108 VPWR.n28 VPWR.t7 60.023
R109 VPWR.n39 VPWR.t3 44.632
R110 VPWR.n39 VPWR.t4 44.632
R111 VPWR.n15 VPWR.t2 43.34
R112 VPWR.n52 VPWR.t9 41.554
R113 VPWR.n52 VPWR.t6 41.554
R114 VPWR.n0 VPWR.t10 30.241
R115 VPWR.n4 VPWR.n3 4.65
R116 VPWR.n6 VPWR.n5 4.65
R117 VPWR.n8 VPWR.n7 4.65
R118 VPWR.n10 VPWR.n9 4.65
R119 VPWR.n12 VPWR.n11 4.65
R120 VPWR.n14 VPWR.n13 4.65
R121 VPWR.n17 VPWR.n16 4.65
R122 VPWR.n19 VPWR.n18 4.65
R123 VPWR.n21 VPWR.n20 4.65
R124 VPWR.n23 VPWR.n22 4.65
R125 VPWR.n25 VPWR.n24 4.65
R126 VPWR.n27 VPWR.n26 4.65
R127 VPWR.n30 VPWR.n29 4.65
R128 VPWR.n32 VPWR.n31 4.65
R129 VPWR.n34 VPWR.n33 4.65
R130 VPWR.n36 VPWR.n35 4.65
R131 VPWR.n38 VPWR.n37 4.65
R132 VPWR.n41 VPWR.n40 4.65
R133 VPWR.n43 VPWR.n42 4.65
R134 VPWR.n45 VPWR.n44 4.65
R135 VPWR.n47 VPWR.n46 4.65
R136 VPWR.n49 VPWR.n48 4.65
R137 VPWR.n51 VPWR.n50 4.65
R138 VPWR.n54 VPWR.n53 3.932
R139 VPWR.n3 VPWR.n2 0.752
R140 VPWR.n4 VPWR.n1 0.3
R141 VPWR.n54 VPWR.n51 0.137
R142 VPWR VPWR.n54 0.123
R143 VPWR.n6 VPWR.n4 0.119
R144 VPWR.n8 VPWR.n6 0.119
R145 VPWR.n10 VPWR.n8 0.119
R146 VPWR.n12 VPWR.n10 0.119
R147 VPWR.n14 VPWR.n12 0.119
R148 VPWR.n17 VPWR.n14 0.119
R149 VPWR.n19 VPWR.n17 0.119
R150 VPWR.n21 VPWR.n19 0.119
R151 VPWR.n23 VPWR.n21 0.119
R152 VPWR.n25 VPWR.n23 0.119
R153 VPWR.n27 VPWR.n25 0.119
R154 VPWR.n30 VPWR.n27 0.119
R155 VPWR.n32 VPWR.n30 0.119
R156 VPWR.n34 VPWR.n32 0.119
R157 VPWR.n36 VPWR.n34 0.119
R158 VPWR.n38 VPWR.n36 0.119
R159 VPWR.n41 VPWR.n38 0.119
R160 VPWR.n43 VPWR.n41 0.119
R161 VPWR.n45 VPWR.n43 0.119
R162 VPWR.n47 VPWR.n45 0.119
R163 VPWR.n49 VPWR.n47 0.119
R164 VPWR.n51 VPWR.n49 0.119
R165 CLK.n0 CLK.t0 292.947
R166 CLK.n0 CLK.t1 209.401
R167 CLK CLK.n0 78.067
R168 SCE.t1 SCE.t2 604.106
R169 SCE.n1 SCE.t3 352.394
R170 SCE.n0 SCE.t0 189.586
R171 SCE.n0 SCE.t1 142.029
R172 SCE SCE.n1 77.631
R173 SCE.n1 SCE.n0 74.085
R174 a_885_21.n0 a_885_21.t3 495.544
R175 a_885_21.n1 a_885_21.t2 351.552
R176 a_885_21.t1 a_885_21.n1 226.125
R177 a_885_21.n0 a_885_21.t0 131.071
R178 a_885_21.n1 a_885_21.n0 74.939
R179 VGND.n11 VGND.t11 152.016
R180 VGND.n0 VGND.t7 149.356
R181 VGND.n46 VGND.t2 145.81
R182 VGND.n30 VGND.n29 130.388
R183 VGND.n42 VGND.n41 109.76
R184 VGND.n55 VGND.n54 107.239
R185 VGND.n17 VGND.n16 106.11
R186 VGND.n2 VGND.n1 76.596
R187 VGND.n16 VGND.t1 74.865
R188 VGND.n1 VGND.t9 57.781
R189 VGND.n41 VGND.t4 41.428
R190 VGND.n41 VGND.t3 41.428
R191 VGND.n16 VGND.t12 40
R192 VGND.n29 VGND.t5 38.571
R193 VGND.n29 VGND.t6 38.571
R194 VGND.n54 VGND.t8 38.571
R195 VGND.n54 VGND.t0 38.571
R196 VGND.n1 VGND.t10 24.78
R197 VGND.n2 VGND.n0 8.863
R198 VGND.n4 VGND.n3 4.65
R199 VGND.n6 VGND.n5 4.65
R200 VGND.n8 VGND.n7 4.65
R201 VGND.n10 VGND.n9 4.65
R202 VGND.n13 VGND.n12 4.65
R203 VGND.n15 VGND.n14 4.65
R204 VGND.n18 VGND.n17 4.65
R205 VGND.n20 VGND.n19 4.65
R206 VGND.n22 VGND.n21 4.65
R207 VGND.n24 VGND.n23 4.65
R208 VGND.n26 VGND.n25 4.65
R209 VGND.n28 VGND.n27 4.65
R210 VGND.n32 VGND.n31 4.65
R211 VGND.n34 VGND.n33 4.65
R212 VGND.n36 VGND.n35 4.65
R213 VGND.n38 VGND.n37 4.65
R214 VGND.n40 VGND.n39 4.65
R215 VGND.n43 VGND.n42 4.65
R216 VGND.n45 VGND.n44 4.65
R217 VGND.n47 VGND.n46 4.65
R218 VGND.n49 VGND.n48 4.65
R219 VGND.n51 VGND.n50 4.65
R220 VGND.n53 VGND.n52 4.65
R221 VGND.n56 VGND.n55 3.932
R222 VGND.n12 VGND.n11 2.635
R223 VGND.n31 VGND.n30 0.752
R224 VGND.n4 VGND.n2 0.3
R225 VGND.n56 VGND.n53 0.137
R226 VGND VGND.n56 0.123
R227 VGND.n6 VGND.n4 0.119
R228 VGND.n8 VGND.n6 0.119
R229 VGND.n10 VGND.n8 0.119
R230 VGND.n13 VGND.n10 0.119
R231 VGND.n15 VGND.n13 0.119
R232 VGND.n18 VGND.n15 0.119
R233 VGND.n20 VGND.n18 0.119
R234 VGND.n22 VGND.n20 0.119
R235 VGND.n24 VGND.n22 0.119
R236 VGND.n26 VGND.n24 0.119
R237 VGND.n28 VGND.n26 0.119
R238 VGND.n32 VGND.n28 0.119
R239 VGND.n34 VGND.n32 0.119
R240 VGND.n36 VGND.n34 0.119
R241 VGND.n38 VGND.n36 0.119
R242 VGND.n40 VGND.n38 0.119
R243 VGND.n43 VGND.n40 0.119
R244 VGND.n45 VGND.n43 0.119
R245 VGND.n47 VGND.n45 0.119
R246 VGND.n49 VGND.n47 0.119
R247 VGND.n51 VGND.n49 0.119
R248 VGND.n53 VGND.n51 0.119
R249 a_1610_159.n1 a_1610_159.t2 406.399
R250 a_1610_159.n0 a_1610_159.t5 318.12
R251 a_1610_159.t1 a_1610_159.n3 262.563
R252 a_1610_159.n0 a_1610_159.t3 194.476
R253 a_1610_159.n1 a_1610_159.t4 130.052
R254 a_1610_159.n2 a_1610_159.n1 100.533
R255 a_1610_159.n2 a_1610_159.t0 93.987
R256 a_1610_159.n3 a_1610_159.n0 92.484
R257 a_1610_159.n3 a_1610_159.n2 9.323
R258 a_193_47.n1 a_193_47.t2 389.542
R259 a_193_47.n1 a_193_47.t5 273.571
R260 a_193_47.t1 a_193_47.n3 249.337
R261 a_193_47.n0 a_193_47.t4 232.651
R262 a_193_47.n0 a_193_47.t3 222.372
R263 a_193_47.n3 a_193_47.t0 207.871
R264 a_193_47.n2 a_193_47.n1 93.104
R265 a_193_47.n3 a_193_47.n2 9.98
R266 a_193_47.n2 a_193_47.n0 7.6
R267 a_1561_47.t1 a_1561_47.t0 111.393
R268 a_791_264.n2 a_791_264.t5 382.743
R269 a_791_264.n0 a_791_264.t2 310.621
R270 a_791_264.t1 a_791_264.n3 216.537
R271 a_791_264.n0 a_791_264.t3 194.941
R272 a_791_264.n1 a_791_264.t0 149.821
R273 a_791_264.n2 a_791_264.t4 138.53
R274 a_791_264.n1 a_791_264.n0 135.659
R275 a_791_264.n3 a_791_264.n2 98.016
R276 a_791_264.n3 a_791_264.n1 48.37
R277 a_1974_47.n0 a_1974_47.t0 70
R278 a_1974_47.n0 a_1974_47.t1 26.393
R279 a_1974_47.n1 a_1974_47.n0 14.4
R280 a_1231_369.t0 a_1231_369.t1 101.578
R281 a_915_47.n0 a_915_47.t4 305.928
R282 a_915_47.n5 a_915_47.n4 221.84
R283 a_915_47.n5 a_915_47.t2 117.17
R284 a_915_47.n2 a_915_47.n1 97.479
R285 a_915_47.n4 a_915_47.n3 92.5
R286 a_915_47.n1 a_915_47.t5 75.384
R287 a_915_47.t0 a_915_47.n5 61.587
R288 a_915_47.n0 a_915_47.t1 46.679
R289 a_915_47.n3 a_915_47.t3 32.197
R290 a_915_47.n4 a_915_47.n2 9.521
R291 a_915_47.n2 a_915_47.n0 7.415
R292 a_729_47.t0 a_729_47.t1 102.857
R293 a_729_369.t0 a_729_369.t1 110.812
R294 Q Q.t1 153.46
R295 Q Q.t0 100.27
R296 a_2135_413.t0 a_2135_413.t1 197
R297 SCD.n0 SCD.t1 206.188
R298 SCD.n0 SCD.t0 183.694
R299 SCD SCD.n0 87.674
R300 a_1226_119.t0 a_1226_119.t1 60
R301 a_1960_413.t0 a_1960_413.t1 143.059
R302 a_381_47.t0 a_381_47.t1 60
C0 VPWR Q 0.21fF
C1 D DE 0.13fF
C2 VGND Q 0.15fF
C3 VPB VPWR 0.28fF
C4 VPWR VGND 0.12fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__sedfxtp_2.ext - technology: sky130A

.subckt sky130_fd_sc_hd__sedfxtp_2 VPWR VGND CLK SCD DE D Q SCE VNB VPB
X0 a_2177_47.t0 a_27_47.t2 a_2051_413.t2 VNB.t16 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X1 a_381_369.t1 D.t0 a_299_47.t3 VPB.t16 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X2 a_1537_413.t1 a_27_47.t3 a_1446_413.t3 VPB.t13 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3 VPWR.t7 DE.t0 a_423_343.t1 VPB.t10 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X4 VPWR.t2 CLK.t0 a_27_47.t0 VPB.t5 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X5 VPWR.t3 SCE.t0 a_885_21.t1 VPB.t7 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X6 VGND.t13 SCE.t1 a_885_21.t0 VNB.t8 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7 VPWR.t0 a_1610_159.t2 a_1537_413.t0 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 a_1610_159.t1 a_1446_413.t4 VPWR.t8 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X9 a_1561_47.t1 a_193_47.t2 a_1446_413.t1 VNB.t6 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X10 VGND.t9 a_2051_413.t4 a_791_264.t0 VNB.t21 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11 VGND.t5 DE.t1 a_423_343.t0 VNB.t10 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12 a_1974_47.t0 a_1610_159.t3 VGND.t0 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13 VGND.t11 a_2051_413.t5 Q.t1 VNB.t20 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14 a_915_47.t2 a_885_21.t2 a_1231_369.t1 VPB.t6 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X15 a_193_47.t0 a_27_47.t4 VGND.t2 VNB.t15 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16 a_2051_413.t0 a_193_47.t3 a_1974_47.t1 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X17 a_729_47.t1 a_423_343.t2 VGND.t12 VNB.t13 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18 a_729_369.t1 DE.t2 VPWR.t6 VPB.t9 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X19 Q.t0 a_2051_413.t6 VGND.t10 VNB.t19 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X20 a_299_47.t1 a_791_264.t2 a_729_47.t0 VNB.t5 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21 a_1446_413.t2 a_27_47.t5 a_915_47.t0 VNB.t14 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X22 a_2135_413.t1 a_193_47.t4 a_2051_413.t1 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23 a_193_47.t1 a_27_47.t6 VPWR.t4 VPB.t12 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X24 a_1231_369.t0 SCD.t0 VPWR.t5 VPB.t15 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X25 a_915_47.t3 SCE.t2 a_1226_119.t0 VNB.t9 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X26 VPWR.t12 a_2051_413.t7 Q.t3 VPB.t21 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X27 a_2051_413.t3 a_27_47.t7 a_1960_413.t0 VPB.t11 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X28 a_299_47.t5 a_791_264.t3 a_729_369.t0 VPB.t17 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X29 a_381_47.t1 D.t1 a_299_47.t4 VNB.t11 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X30 VPWR.t9 a_791_264.t4 a_2135_413.t0 VPB.t18 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X31 VGND.t1 a_1610_159.t4 a_1561_47.t0 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X32 Q.t2 a_2051_413.t8 VPWR.t11 VPB.t20 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X33 VPWR.t13 a_423_343.t3 a_381_369.t0 VPB.t14 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X34 a_915_47.t4 SCE.t3 a_299_47.t2 VPB.t8 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X35 a_1960_413.t1 a_1610_159.t5 VPWR.t1 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X36 a_1226_119.t1 SCD.t1 VGND.t3 VNB.t17 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X37 VGND.t7 a_791_264.t5 a_2177_47.t1 VNB.t18 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X38 a_1446_413.t0 a_193_47.t5 a_915_47.t5 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X39 a_915_47.t1 a_885_21.t3 a_299_47.t0 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X40 VPWR.t10 a_2051_413.t9 a_791_264.t1 VPB.t19 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X41 VGND.t8 CLK.t1 a_27_47.t1 VNB.t7 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X42 VGND.t4 DE.t3 a_381_47.t0 VNB.t12 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X43 a_1610_159.t0 a_1446_413.t5 VGND.t6 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
R0 a_27_47.n1 a_27_47.t2 443.438
R1 a_27_47.n0 a_27_47.t5 269.985
R2 a_27_47.n3 a_27_47.t6 263.405
R3 a_27_47.n1 a_27_47.t7 254.388
R4 a_27_47.t0 a_27_47.n5 244.156
R5 a_27_47.n3 a_27_47.t4 228.059
R6 a_27_47.n4 a_27_47.t1 195.871
R7 a_27_47.n0 a_27_47.t3 142.49
R8 a_27_47.n2 a_27_47.n1 113.844
R9 a_27_47.n4 a_27_47.n3 76
R10 a_27_47.n5 a_27_47.n4 35.339
R11 a_27_47.n5 a_27_47.n2 10.69
R12 a_27_47.n2 a_27_47.n0 2.9
R13 a_2051_413.n5 a_2051_413.n4 398.525
R14 a_2051_413.n3 a_2051_413.t9 269.919
R15 a_2051_413.n1 a_2051_413.t7 212.079
R16 a_2051_413.n2 a_2051_413.t8 212.079
R17 a_2051_413.n3 a_2051_413.t4 176.733
R18 a_2051_413.n4 a_2051_413.n3 176.181
R19 a_2051_413.n4 a_2051_413.n0 159.603
R20 a_2051_413.n1 a_2051_413.t5 139.779
R21 a_2051_413.n2 a_2051_413.t6 139.779
R22 a_2051_413.n0 a_2051_413.t2 76.666
R23 a_2051_413.n3 a_2051_413.n2 70.839
R24 a_2051_413.t1 a_2051_413.n5 63.321
R25 a_2051_413.n5 a_2051_413.t3 63.321
R26 a_2051_413.n2 a_2051_413.n1 61.345
R27 a_2051_413.n0 a_2051_413.t0 50
R28 a_2177_47.t1 a_2177_47.t0 93.059
R29 VNB.t4 VNB.t8 8836.4
R30 VNB.t18 VNB.t21 6082.35
R31 VNB.t12 VNB.t10 6082.35
R32 VNB.t15 VNB.t11 6082.35
R33 VNB.t3 VNB.t1 5346.86
R34 VNB VNB.t7 4270.59
R35 VNB.t9 VNB.t14 4015.64
R36 VNB.t0 VNB.t16 3429.41
R37 VNB.t6 VNB.t2 3429.41
R38 VNB.t13 VNB.t5 3300
R39 VNB.t1 VNB.t0 3138.24
R40 VNB.t2 VNB.t3 3130.33
R41 VNB.t16 VNB.t18 3073.53
R42 VNB.t14 VNB.t6 2847.06
R43 VNB.t10 VNB.t13 2847.06
R44 VNB.t8 VNB.t17 2717.65
R45 VNB.t5 VNB.t4 2717.65
R46 VNB.t7 VNB.t15 2717.65
R47 VNB.t17 VNB.t9 2329.41
R48 VNB.t11 VNB.t12 2329.41
R49 VNB.t21 VNB.t19 2303.7
R50 VNB.t19 VNB.t20 2030.77
R51 D.n0 D.t1 216.76
R52 D.n0 D.t0 215.106
R53 D D.n0 34.479
R54 a_299_47.n1 a_299_47.t3 321.627
R55 a_299_47.n3 a_299_47.n2 233.623
R56 a_299_47.n1 a_299_47.t4 139.932
R57 a_299_47.t2 a_299_47.n3 53.867
R58 a_299_47.n3 a_299_47.t5 41.554
R59 a_299_47.n0 a_299_47.t0 37.55
R60 a_299_47.n0 a_299_47.t1 36.873
R61 a_299_47.n2 a_299_47.n1 8.177
R62 a_299_47.n2 a_299_47.n0 8.115
R63 a_381_369.t0 a_381_369.t1 64.64
R64 VPB.t18 VPB.t19 624.454
R65 VPB.t8 VPB.t7 622.849
R66 VPB.t4 VPB.t3 556.386
R67 VPB.t14 VPB.t10 556.386
R68 VPB.t12 VPB.t16 556.386
R69 VPB.t2 VPB.t4 390.654
R70 VPB.t6 VPB.t1 383.22
R71 VPB.t7 VPB.t15 351.016
R72 VPB.t0 VPB.t18 337.383
R73 VPB.t15 VPB.t6 309.152
R74 VPB.t13 VPB.t2 304.828
R75 VPB.t9 VPB.t17 301.869
R76 VPB.t19 VPB.t20 287.071
R77 VPB.t17 VPB.t8 272.274
R78 VPB.t3 VPB.t11 269.314
R79 VPB.t10 VPB.t9 260.436
R80 VPB.t1 VPB.t13 256.559
R81 VPB.t20 VPB.t21 248.598
R82 VPB.t11 VPB.t0 248.598
R83 VPB.t5 VPB.t12 248.598
R84 VPB.t16 VPB.t14 213.084
R85 VPB VPB.t5 142.056
R86 a_1446_413.n3 a_1446_413.n2 388.236
R87 a_1446_413.n0 a_1446_413.t5 230.482
R88 a_1446_413.n0 a_1446_413.t4 196.013
R89 a_1446_413.n2 a_1446_413.n1 183.768
R90 a_1446_413.n2 a_1446_413.n0 95.938
R91 a_1446_413.n3 a_1446_413.t3 72.702
R92 a_1446_413.t0 a_1446_413.n3 70.357
R93 a_1446_413.n1 a_1446_413.t1 51.666
R94 a_1446_413.n1 a_1446_413.t2 45
R95 a_1537_413.t0 a_1537_413.t1 171.202
R96 DE.n0 DE.t2 319.725
R97 DE.n2 DE.n1 238.689
R98 DE.n0 DE.t0 178.339
R99 DE.n1 DE.n0 147.813
R100 DE.n2 DE.t3 130.384
R101 DE.n1 DE.t1 130.14
R102 DE DE.n2 82.892
R103 a_423_343.n1 a_423_343.t3 299.566
R104 a_423_343.n0 a_423_343.t2 258.036
R105 a_423_343.t1 a_423_343.n1 230.699
R106 a_423_343.n0 a_423_343.t0 151.679
R107 a_423_343.n1 a_423_343.n0 11.133
R108 VPWR.n7 VPWR.t9 378.842
R109 VPWR.n16 VPWR.t1 375.462
R110 VPWR.n58 VPWR.n57 311.893
R111 VPWR.n34 VPWR.n33 306.598
R112 VPWR.n49 VPWR.t13 228.681
R113 VPWR.n45 VPWR.n44 176.72
R114 VPWR.n21 VPWR.n20 171.436
R115 VPWR.n2 VPWR.t12 160.596
R116 VPWR.n1 VPWR.n0 140.629
R117 VPWR.n20 VPWR.t0 106.098
R118 VPWR.n0 VPWR.t10 61.911
R119 VPWR.n33 VPWR.t5 61.562
R120 VPWR.n33 VPWR.t3 60.023
R121 VPWR.n44 VPWR.t6 44.632
R122 VPWR.n44 VPWR.t7 44.632
R123 VPWR.n20 VPWR.t8 43.34
R124 VPWR.n57 VPWR.t4 41.554
R125 VPWR.n57 VPWR.t2 41.554
R126 VPWR.n0 VPWR.t11 30.242
R127 VPWR.n2 VPWR.n1 8.848
R128 VPWR.n4 VPWR.n3 4.65
R129 VPWR.n6 VPWR.n5 4.65
R130 VPWR.n9 VPWR.n8 4.65
R131 VPWR.n11 VPWR.n10 4.65
R132 VPWR.n13 VPWR.n12 4.65
R133 VPWR.n15 VPWR.n14 4.65
R134 VPWR.n17 VPWR.n16 4.65
R135 VPWR.n19 VPWR.n18 4.65
R136 VPWR.n22 VPWR.n21 4.65
R137 VPWR.n24 VPWR.n23 4.65
R138 VPWR.n26 VPWR.n25 4.65
R139 VPWR.n28 VPWR.n27 4.65
R140 VPWR.n30 VPWR.n29 4.65
R141 VPWR.n32 VPWR.n31 4.65
R142 VPWR.n35 VPWR.n34 4.65
R143 VPWR.n37 VPWR.n36 4.65
R144 VPWR.n39 VPWR.n38 4.65
R145 VPWR.n41 VPWR.n40 4.65
R146 VPWR.n43 VPWR.n42 4.65
R147 VPWR.n46 VPWR.n45 4.65
R148 VPWR.n48 VPWR.n47 4.65
R149 VPWR.n50 VPWR.n49 4.65
R150 VPWR.n52 VPWR.n51 4.65
R151 VPWR.n54 VPWR.n53 4.65
R152 VPWR.n56 VPWR.n55 4.65
R153 VPWR.n59 VPWR.n58 3.932
R154 VPWR.n8 VPWR.n7 0.752
R155 VPWR.n4 VPWR.n2 0.315
R156 VPWR.n59 VPWR.n56 0.137
R157 VPWR VPWR.n59 0.123
R158 VPWR.n6 VPWR.n4 0.119
R159 VPWR.n9 VPWR.n6 0.119
R160 VPWR.n11 VPWR.n9 0.119
R161 VPWR.n13 VPWR.n11 0.119
R162 VPWR.n15 VPWR.n13 0.119
R163 VPWR.n17 VPWR.n15 0.119
R164 VPWR.n19 VPWR.n17 0.119
R165 VPWR.n22 VPWR.n19 0.119
R166 VPWR.n24 VPWR.n22 0.119
R167 VPWR.n26 VPWR.n24 0.119
R168 VPWR.n28 VPWR.n26 0.119
R169 VPWR.n30 VPWR.n28 0.119
R170 VPWR.n32 VPWR.n30 0.119
R171 VPWR.n35 VPWR.n32 0.119
R172 VPWR.n37 VPWR.n35 0.119
R173 VPWR.n39 VPWR.n37 0.119
R174 VPWR.n41 VPWR.n39 0.119
R175 VPWR.n43 VPWR.n41 0.119
R176 VPWR.n46 VPWR.n43 0.119
R177 VPWR.n48 VPWR.n46 0.119
R178 VPWR.n50 VPWR.n48 0.119
R179 VPWR.n52 VPWR.n50 0.119
R180 VPWR.n54 VPWR.n52 0.119
R181 VPWR.n56 VPWR.n54 0.119
R182 CLK.n0 CLK.t0 292.947
R183 CLK.n0 CLK.t1 209.401
R184 CLK CLK.n0 78.067
R185 SCE.t1 SCE.t2 604.106
R186 SCE.n1 SCE.t3 352.394
R187 SCE.n0 SCE.t0 189.586
R188 SCE.n0 SCE.t1 142.029
R189 SCE SCE.n1 77.631
R190 SCE.n1 SCE.n0 74.085
R191 a_885_21.n0 a_885_21.t3 495.544
R192 a_885_21.n1 a_885_21.t2 351.552
R193 a_885_21.t1 a_885_21.n1 226.125
R194 a_885_21.n0 a_885_21.t0 131.071
R195 a_885_21.n1 a_885_21.n0 74.939
R196 VGND.n16 VGND.t0 152.016
R197 VGND.n5 VGND.t7 149.356
R198 VGND.n51 VGND.t4 145.81
R199 VGND.n35 VGND.n34 130.388
R200 VGND.n2 VGND.t11 110.253
R201 VGND.n47 VGND.n46 109.76
R202 VGND.n60 VGND.n59 107.239
R203 VGND.n22 VGND.n21 106.11
R204 VGND.n21 VGND.t6 74.865
R205 VGND.n1 VGND.n0 72.154
R206 VGND.n0 VGND.t9 57.779
R207 VGND.n46 VGND.t12 41.428
R208 VGND.n46 VGND.t5 41.428
R209 VGND.n21 VGND.t1 40
R210 VGND.n34 VGND.t3 38.571
R211 VGND.n34 VGND.t13 38.571
R212 VGND.n59 VGND.t2 38.571
R213 VGND.n59 VGND.t8 38.571
R214 VGND.n0 VGND.t10 24.782
R215 VGND.n2 VGND.n1 8.848
R216 VGND.n6 VGND.n5 4.894
R217 VGND.n4 VGND.n3 4.65
R218 VGND.n7 VGND.n6 4.65
R219 VGND.n9 VGND.n8 4.65
R220 VGND.n11 VGND.n10 4.65
R221 VGND.n13 VGND.n12 4.65
R222 VGND.n15 VGND.n14 4.65
R223 VGND.n18 VGND.n17 4.65
R224 VGND.n20 VGND.n19 4.65
R225 VGND.n23 VGND.n22 4.65
R226 VGND.n25 VGND.n24 4.65
R227 VGND.n27 VGND.n26 4.65
R228 VGND.n29 VGND.n28 4.65
R229 VGND.n31 VGND.n30 4.65
R230 VGND.n33 VGND.n32 4.65
R231 VGND.n37 VGND.n36 4.65
R232 VGND.n39 VGND.n38 4.65
R233 VGND.n41 VGND.n40 4.65
R234 VGND.n43 VGND.n42 4.65
R235 VGND.n45 VGND.n44 4.65
R236 VGND.n48 VGND.n47 4.65
R237 VGND.n50 VGND.n49 4.65
R238 VGND.n52 VGND.n51 4.65
R239 VGND.n54 VGND.n53 4.65
R240 VGND.n56 VGND.n55 4.65
R241 VGND.n58 VGND.n57 4.65
R242 VGND.n61 VGND.n60 3.932
R243 VGND.n17 VGND.n16 2.635
R244 VGND.n36 VGND.n35 0.752
R245 VGND.n4 VGND.n2 0.315
R246 VGND.n61 VGND.n58 0.137
R247 VGND VGND.n61 0.123
R248 VGND.n7 VGND.n4 0.119
R249 VGND.n9 VGND.n7 0.119
R250 VGND.n11 VGND.n9 0.119
R251 VGND.n13 VGND.n11 0.119
R252 VGND.n15 VGND.n13 0.119
R253 VGND.n18 VGND.n15 0.119
R254 VGND.n20 VGND.n18 0.119
R255 VGND.n23 VGND.n20 0.119
R256 VGND.n25 VGND.n23 0.119
R257 VGND.n27 VGND.n25 0.119
R258 VGND.n29 VGND.n27 0.119
R259 VGND.n31 VGND.n29 0.119
R260 VGND.n33 VGND.n31 0.119
R261 VGND.n37 VGND.n33 0.119
R262 VGND.n39 VGND.n37 0.119
R263 VGND.n41 VGND.n39 0.119
R264 VGND.n43 VGND.n41 0.119
R265 VGND.n45 VGND.n43 0.119
R266 VGND.n48 VGND.n45 0.119
R267 VGND.n50 VGND.n48 0.119
R268 VGND.n52 VGND.n50 0.119
R269 VGND.n54 VGND.n52 0.119
R270 VGND.n56 VGND.n54 0.119
R271 VGND.n58 VGND.n56 0.119
R272 a_1610_159.n1 a_1610_159.t2 406.399
R273 a_1610_159.n0 a_1610_159.t5 318.12
R274 a_1610_159.t1 a_1610_159.n3 262.563
R275 a_1610_159.n0 a_1610_159.t3 194.476
R276 a_1610_159.n1 a_1610_159.t4 130.052
R277 a_1610_159.n2 a_1610_159.n1 100.533
R278 a_1610_159.n2 a_1610_159.t0 93.987
R279 a_1610_159.n3 a_1610_159.n0 92.484
R280 a_1610_159.n3 a_1610_159.n2 9.323
R281 a_193_47.n1 a_193_47.t2 389.542
R282 a_193_47.n1 a_193_47.t5 273.571
R283 a_193_47.t1 a_193_47.n3 249.337
R284 a_193_47.n0 a_193_47.t4 232.651
R285 a_193_47.n0 a_193_47.t3 222.372
R286 a_193_47.n3 a_193_47.t0 207.871
R287 a_193_47.n2 a_193_47.n1 93.104
R288 a_193_47.n3 a_193_47.n2 9.98
R289 a_193_47.n2 a_193_47.n0 7.6
R290 a_1561_47.t0 a_1561_47.t1 111.393
R291 a_791_264.n2 a_791_264.t5 382.743
R292 a_791_264.n0 a_791_264.t2 310.621
R293 a_791_264.t1 a_791_264.n3 216.537
R294 a_791_264.n0 a_791_264.t3 194.941
R295 a_791_264.n1 a_791_264.t0 149.821
R296 a_791_264.n2 a_791_264.t4 138.53
R297 a_791_264.n1 a_791_264.n0 135.659
R298 a_791_264.n3 a_791_264.n2 98.016
R299 a_791_264.n3 a_791_264.n1 48.37
R300 a_1974_47.n0 a_1974_47.t1 70
R301 a_1974_47.n0 a_1974_47.t0 26.393
R302 a_1974_47.n1 a_1974_47.n0 14.4
R303 Q Q.n0 124.895
R304 Q Q.n1 63.679
R305 Q.n0 Q.t3 26.595
R306 Q.n0 Q.t2 26.595
R307 Q.n1 Q.t1 24.923
R308 Q.n1 Q.t0 24.923
R309 a_1231_369.t0 a_1231_369.t1 101.578
R310 a_915_47.n0 a_915_47.t4 305.928
R311 a_915_47.n5 a_915_47.n4 221.84
R312 a_915_47.n5 a_915_47.t5 117.17
R313 a_915_47.n2 a_915_47.n1 97.479
R314 a_915_47.n4 a_915_47.n3 92.5
R315 a_915_47.n1 a_915_47.t0 75.384
R316 a_915_47.t2 a_915_47.n5 61.587
R317 a_915_47.n0 a_915_47.t1 46.679
R318 a_915_47.n3 a_915_47.t3 32.197
R319 a_915_47.n4 a_915_47.n2 9.521
R320 a_915_47.n2 a_915_47.n0 7.415
R321 a_729_47.t0 a_729_47.t1 102.857
R322 a_729_369.t0 a_729_369.t1 110.812
R323 a_2135_413.t0 a_2135_413.t1 197
R324 SCD.n0 SCD.t1 206.188
R325 SCD.n0 SCD.t0 183.694
R326 SCD SCD.n0 87.674
R327 a_1226_119.t0 a_1226_119.t1 60
R328 a_1960_413.t0 a_1960_413.t1 143.059
R329 a_381_47.t0 a_381_47.t1 60
C0 VPWR Q 0.37fF
C1 D DE 0.13fF
C2 VGND Q 0.25fF
C3 VPB VPWR 0.30fF
C4 VPWR VGND 0.15fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__sedfxtp_4.ext - technology: sky130A

.subckt sky130_fd_sc_hd__sedfxtp_4 VPWR VGND CLK SCD DE D Q SCE VNB VPB
X0 a_2177_47.t0 a_27_47.t2 a_2051_413.t2 VNB.t16 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X1 a_381_369.t1 D.t0 a_299_47.t2 VPB.t15 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X2 a_1537_413.t1 a_27_47.t3 a_1446_413.t3 VPB.t14 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3 VPWR.t15 DE.t0 a_423_343.t1 VPB.t11 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X4 VPWR.t3 CLK.t0 a_27_47.t1 VPB.t5 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X5 VPWR.t4 SCE.t0 a_885_21.t1 VPB.t6 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X6 VGND.t13 SCE.t1 a_885_21.t0 VNB.t9 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7 VPWR.t1 a_1610_159.t2 a_1537_413.t0 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 a_1610_159.t0 a_1446_413.t4 VPWR.t0 VPB.t8 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X9 a_1561_47.t1 a_193_47.t2 a_1446_413.t1 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X10 VPWR.t12 a_2051_413.t4 Q.t3 VPB.t21 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 VGND.t12 a_2051_413.t5 a_791_264.t1 VNB.t22 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12 VGND.t14 DE.t1 a_423_343.t0 VNB.t12 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13 a_1974_47.t0 a_1610_159.t3 VGND.t2 VNB.t5 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14 Q.t2 a_2051_413.t6 VPWR.t11 VPB.t20 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 VGND.t11 a_2051_413.t7 Q.t7 VNB.t21 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X16 a_915_47.t5 a_885_21.t2 a_1231_369.t1 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X17 a_193_47.t1 a_27_47.t4 VGND.t4 VNB.t15 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18 a_2051_413.t1 a_193_47.t3 a_1974_47.t1 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X19 a_729_47.t0 a_423_343.t2 VGND.t6 VNB.t13 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20 a_729_369.t1 DE.t2 VPWR.t14 VPB.t9 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X21 Q.t6 a_2051_413.t8 VGND.t10 VNB.t20 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X22 a_299_47.t4 a_791_264.t2 a_729_47.t1 VNB.t23 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23 a_1446_413.t2 a_27_47.t5 a_915_47.t0 VNB.t14 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X24 a_2135_413.t1 a_193_47.t4 a_2051_413.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X25 Q.t5 a_2051_413.t9 VGND.t9 VNB.t19 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X26 a_193_47.t0 a_27_47.t6 VPWR.t5 VPB.t13 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X27 a_1231_369.t0 SCD.t0 VPWR.t13 VPB.t23 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X28 a_915_47.t1 SCE.t2 a_1226_119.t0 VNB.t10 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X29 VPWR.t10 a_2051_413.t10 Q.t1 VPB.t19 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X30 a_2051_413.t3 a_27_47.t7 a_1960_413.t0 VPB.t12 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X31 a_299_47.t5 a_791_264.t3 a_729_369.t0 VPB.t22 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X32 a_381_47.t0 D.t1 a_299_47.t3 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X33 VPWR.t7 a_791_264.t4 a_2135_413.t0 VPB.t16 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X34 VGND.t3 a_1610_159.t4 a_1561_47.t0 VNB.t6 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X35 Q.t0 a_2051_413.t11 VPWR.t9 VPB.t18 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X36 VPWR.t6 a_423_343.t3 a_381_369.t0 VPB.t10 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X37 a_915_47.t2 SCE.t3 a_299_47.t1 VPB.t7 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X38 a_1960_413.t1 a_1610_159.t5 VPWR.t2 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X39 a_1226_119.t1 SCD.t1 VGND.t0 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X40 VGND.t7 a_791_264.t5 a_2177_47.t1 VNB.t17 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X41 a_1446_413.t0 a_193_47.t5 a_915_47.t3 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X42 a_915_47.t4 a_885_21.t3 a_299_47.t0 VNB.t8 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X43 VPWR.t8 a_2051_413.t12 a_791_264.t0 VPB.t17 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X44 VGND.t8 a_2051_413.t13 Q.t4 VNB.t18 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X45 VGND.t5 CLK.t1 a_27_47.t0 VNB.t7 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X46 VGND.t15 DE.t3 a_381_47.t1 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X47 a_1610_159.t1 a_1446_413.t5 VGND.t1 VNB.t11 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
R0 a_27_47.n1 a_27_47.t2 443.438
R1 a_27_47.n0 a_27_47.t5 269.985
R2 a_27_47.n3 a_27_47.t6 263.405
R3 a_27_47.n1 a_27_47.t7 254.388
R4 a_27_47.t1 a_27_47.n5 244.156
R5 a_27_47.n3 a_27_47.t4 228.059
R6 a_27_47.n4 a_27_47.t0 195.871
R7 a_27_47.n0 a_27_47.t3 142.49
R8 a_27_47.n2 a_27_47.n1 113.844
R9 a_27_47.n4 a_27_47.n3 76
R10 a_27_47.n5 a_27_47.n4 35.339
R11 a_27_47.n5 a_27_47.n2 10.69
R12 a_27_47.n2 a_27_47.n0 2.9
R13 a_2051_413.n7 a_2051_413.n6 398.525
R14 a_2051_413.n5 a_2051_413.t12 269.919
R15 a_2051_413.n1 a_2051_413.t4 212.079
R16 a_2051_413.n2 a_2051_413.t6 212.079
R17 a_2051_413.n3 a_2051_413.t10 212.079
R18 a_2051_413.n4 a_2051_413.t11 212.079
R19 a_2051_413.n5 a_2051_413.t5 176.733
R20 a_2051_413.n6 a_2051_413.n5 176.181
R21 a_2051_413.n6 a_2051_413.n0 159.603
R22 a_2051_413.n1 a_2051_413.t13 139.779
R23 a_2051_413.n2 a_2051_413.t9 139.779
R24 a_2051_413.n3 a_2051_413.t7 139.779
R25 a_2051_413.n4 a_2051_413.t8 139.779
R26 a_2051_413.n0 a_2051_413.t2 76.666
R27 a_2051_413.n5 a_2051_413.n4 70.839
R28 a_2051_413.t0 a_2051_413.n7 63.321
R29 a_2051_413.n7 a_2051_413.t3 63.321
R30 a_2051_413.n2 a_2051_413.n1 61.345
R31 a_2051_413.n3 a_2051_413.n2 61.345
R32 a_2051_413.n4 a_2051_413.n3 61.345
R33 a_2051_413.n0 a_2051_413.t1 50
R34 a_2177_47.t1 a_2177_47.t0 93.059
R35 VNB.t8 VNB.t9 8836.4
R36 VNB.t17 VNB.t22 6082.35
R37 VNB.t0 VNB.t12 6082.35
R38 VNB.t15 VNB.t4 6082.35
R39 VNB.t11 VNB.t5 5346.86
R40 VNB VNB.t7 4270.59
R41 VNB.t10 VNB.t14 4015.64
R42 VNB.t3 VNB.t16 3429.41
R43 VNB.t2 VNB.t6 3429.41
R44 VNB.t13 VNB.t23 3300
R45 VNB.t5 VNB.t3 3138.24
R46 VNB.t6 VNB.t11 3130.33
R47 VNB.t16 VNB.t17 3073.53
R48 VNB.t14 VNB.t2 2847.06
R49 VNB.t12 VNB.t13 2847.06
R50 VNB.t9 VNB.t1 2717.65
R51 VNB.t23 VNB.t8 2717.65
R52 VNB.t7 VNB.t15 2717.65
R53 VNB.t1 VNB.t10 2329.41
R54 VNB.t4 VNB.t0 2329.41
R55 VNB.t22 VNB.t20 2303.7
R56 VNB.t19 VNB.t18 2030.77
R57 VNB.t21 VNB.t19 2030.77
R58 VNB.t20 VNB.t21 2030.77
R59 D.n0 D.t1 216.76
R60 D.n0 D.t0 215.106
R61 D D.n0 34.479
R62 a_299_47.n1 a_299_47.t2 321.627
R63 a_299_47.n3 a_299_47.n2 233.623
R64 a_299_47.n1 a_299_47.t3 139.932
R65 a_299_47.t1 a_299_47.n3 53.867
R66 a_299_47.n3 a_299_47.t5 41.554
R67 a_299_47.n0 a_299_47.t0 37.55
R68 a_299_47.n0 a_299_47.t4 36.873
R69 a_299_47.n2 a_299_47.n1 8.177
R70 a_299_47.n2 a_299_47.n0 8.115
R71 a_381_369.t0 a_381_369.t1 64.64
R72 VPB.t16 VPB.t17 624.454
R73 VPB.t7 VPB.t6 622.849
R74 VPB.t8 VPB.t3 556.386
R75 VPB.t10 VPB.t11 556.386
R76 VPB.t13 VPB.t15 556.386
R77 VPB.t2 VPB.t8 390.654
R78 VPB.t4 VPB.t1 383.22
R79 VPB.t6 VPB.t23 351.016
R80 VPB.t0 VPB.t16 337.383
R81 VPB.t23 VPB.t4 309.152
R82 VPB.t14 VPB.t2 304.828
R83 VPB.t9 VPB.t22 301.869
R84 VPB.t17 VPB.t18 287.071
R85 VPB.t22 VPB.t7 272.274
R86 VPB.t3 VPB.t12 269.314
R87 VPB.t11 VPB.t9 260.436
R88 VPB.t1 VPB.t14 256.559
R89 VPB.t20 VPB.t21 248.598
R90 VPB.t19 VPB.t20 248.598
R91 VPB.t18 VPB.t19 248.598
R92 VPB.t12 VPB.t0 248.598
R93 VPB.t5 VPB.t13 248.598
R94 VPB.t15 VPB.t10 213.084
R95 VPB VPB.t5 142.056
R96 a_1446_413.n3 a_1446_413.n2 388.236
R97 a_1446_413.n0 a_1446_413.t5 230.482
R98 a_1446_413.n0 a_1446_413.t4 196.013
R99 a_1446_413.n2 a_1446_413.n1 183.768
R100 a_1446_413.n2 a_1446_413.n0 95.938
R101 a_1446_413.n3 a_1446_413.t3 72.702
R102 a_1446_413.t0 a_1446_413.n3 70.357
R103 a_1446_413.n1 a_1446_413.t1 51.666
R104 a_1446_413.n1 a_1446_413.t2 45
R105 a_1537_413.t0 a_1537_413.t1 171.202
R106 DE.n0 DE.t2 319.725
R107 DE.n2 DE.n1 238.689
R108 DE.n0 DE.t0 178.339
R109 DE.n1 DE.n0 147.813
R110 DE.n2 DE.t3 130.384
R111 DE.n1 DE.t1 130.14
R112 DE DE.n2 82.892
R113 a_423_343.n1 a_423_343.t3 299.566
R114 a_423_343.n0 a_423_343.t2 258.036
R115 a_423_343.t1 a_423_343.n1 230.699
R116 a_423_343.n0 a_423_343.t0 151.679
R117 a_423_343.n1 a_423_343.n0 11.133
R118 VPWR.n13 VPWR.t7 378.842
R119 VPWR.n22 VPWR.t2 375.462
R120 VPWR.n64 VPWR.n63 311.893
R121 VPWR.n40 VPWR.n39 306.598
R122 VPWR.n55 VPWR.t6 228.681
R123 VPWR.n51 VPWR.n50 176.72
R124 VPWR.n27 VPWR.n26 171.436
R125 VPWR.n2 VPWR.t12 160.503
R126 VPWR.n6 VPWR.n5 140.629
R127 VPWR.n1 VPWR.n0 135.124
R128 VPWR.n26 VPWR.t1 106.098
R129 VPWR.n5 VPWR.t8 61.911
R130 VPWR.n39 VPWR.t13 61.562
R131 VPWR.n39 VPWR.t4 60.023
R132 VPWR.n50 VPWR.t14 44.632
R133 VPWR.n50 VPWR.t15 44.632
R134 VPWR.n26 VPWR.t0 43.34
R135 VPWR.n63 VPWR.t5 41.554
R136 VPWR.n63 VPWR.t3 41.554
R137 VPWR.n5 VPWR.t9 30.242
R138 VPWR.n0 VPWR.t11 26.595
R139 VPWR.n0 VPWR.t10 26.595
R140 VPWR.n2 VPWR.n1 21.148
R141 VPWR.n7 VPWR.n6 4.894
R142 VPWR.n4 VPWR.n3 4.65
R143 VPWR.n8 VPWR.n7 4.65
R144 VPWR.n10 VPWR.n9 4.65
R145 VPWR.n12 VPWR.n11 4.65
R146 VPWR.n15 VPWR.n14 4.65
R147 VPWR.n17 VPWR.n16 4.65
R148 VPWR.n19 VPWR.n18 4.65
R149 VPWR.n21 VPWR.n20 4.65
R150 VPWR.n23 VPWR.n22 4.65
R151 VPWR.n25 VPWR.n24 4.65
R152 VPWR.n28 VPWR.n27 4.65
R153 VPWR.n30 VPWR.n29 4.65
R154 VPWR.n32 VPWR.n31 4.65
R155 VPWR.n34 VPWR.n33 4.65
R156 VPWR.n36 VPWR.n35 4.65
R157 VPWR.n38 VPWR.n37 4.65
R158 VPWR.n41 VPWR.n40 4.65
R159 VPWR.n43 VPWR.n42 4.65
R160 VPWR.n45 VPWR.n44 4.65
R161 VPWR.n47 VPWR.n46 4.65
R162 VPWR.n49 VPWR.n48 4.65
R163 VPWR.n52 VPWR.n51 4.65
R164 VPWR.n54 VPWR.n53 4.65
R165 VPWR.n56 VPWR.n55 4.65
R166 VPWR.n58 VPWR.n57 4.65
R167 VPWR.n60 VPWR.n59 4.65
R168 VPWR.n62 VPWR.n61 4.65
R169 VPWR.n65 VPWR.n64 3.932
R170 VPWR.n14 VPWR.n13 0.752
R171 VPWR.n4 VPWR.n2 0.438
R172 VPWR.n65 VPWR.n62 0.137
R173 VPWR VPWR.n65 0.123
R174 VPWR.n8 VPWR.n4 0.119
R175 VPWR.n10 VPWR.n8 0.119
R176 VPWR.n12 VPWR.n10 0.119
R177 VPWR.n15 VPWR.n12 0.119
R178 VPWR.n17 VPWR.n15 0.119
R179 VPWR.n19 VPWR.n17 0.119
R180 VPWR.n21 VPWR.n19 0.119
R181 VPWR.n23 VPWR.n21 0.119
R182 VPWR.n25 VPWR.n23 0.119
R183 VPWR.n28 VPWR.n25 0.119
R184 VPWR.n30 VPWR.n28 0.119
R185 VPWR.n32 VPWR.n30 0.119
R186 VPWR.n34 VPWR.n32 0.119
R187 VPWR.n36 VPWR.n34 0.119
R188 VPWR.n38 VPWR.n36 0.119
R189 VPWR.n41 VPWR.n38 0.119
R190 VPWR.n43 VPWR.n41 0.119
R191 VPWR.n45 VPWR.n43 0.119
R192 VPWR.n47 VPWR.n45 0.119
R193 VPWR.n49 VPWR.n47 0.119
R194 VPWR.n52 VPWR.n49 0.119
R195 VPWR.n54 VPWR.n52 0.119
R196 VPWR.n56 VPWR.n54 0.119
R197 VPWR.n58 VPWR.n56 0.119
R198 VPWR.n60 VPWR.n58 0.119
R199 VPWR.n62 VPWR.n60 0.119
R200 CLK.n0 CLK.t0 292.947
R201 CLK.n0 CLK.t1 209.401
R202 CLK CLK.n0 78.067
R203 SCE.t1 SCE.t2 604.106
R204 SCE.n1 SCE.t3 352.394
R205 SCE.n0 SCE.t0 189.586
R206 SCE.n0 SCE.t1 142.029
R207 SCE SCE.n1 77.631
R208 SCE.n1 SCE.n0 74.085
R209 a_885_21.n0 a_885_21.t3 495.544
R210 a_885_21.n1 a_885_21.t2 351.552
R211 a_885_21.t1 a_885_21.n1 226.125
R212 a_885_21.n0 a_885_21.t0 131.071
R213 a_885_21.n1 a_885_21.n0 74.939
R214 VGND.n22 VGND.t2 152.016
R215 VGND.n11 VGND.t7 149.356
R216 VGND.n57 VGND.t15 145.81
R217 VGND.n41 VGND.n40 130.388
R218 VGND.n2 VGND.t8 110.159
R219 VGND.n53 VGND.n52 109.76
R220 VGND.n66 VGND.n65 107.239
R221 VGND.n28 VGND.n27 106.11
R222 VGND.n1 VGND.n0 75.214
R223 VGND.n27 VGND.t1 74.865
R224 VGND.n6 VGND.n5 72.154
R225 VGND.n5 VGND.t12 57.779
R226 VGND.n52 VGND.t6 41.428
R227 VGND.n52 VGND.t14 41.428
R228 VGND.n27 VGND.t3 40
R229 VGND.n40 VGND.t0 38.571
R230 VGND.n40 VGND.t13 38.571
R231 VGND.n65 VGND.t4 38.571
R232 VGND.n65 VGND.t5 38.571
R233 VGND.n0 VGND.t9 24.923
R234 VGND.n0 VGND.t11 24.923
R235 VGND.n5 VGND.t10 24.782
R236 VGND.n2 VGND.n1 21.148
R237 VGND.n7 VGND.n6 4.894
R238 VGND.n12 VGND.n11 4.894
R239 VGND.n4 VGND.n3 4.65
R240 VGND.n8 VGND.n7 4.65
R241 VGND.n10 VGND.n9 4.65
R242 VGND.n13 VGND.n12 4.65
R243 VGND.n15 VGND.n14 4.65
R244 VGND.n17 VGND.n16 4.65
R245 VGND.n19 VGND.n18 4.65
R246 VGND.n21 VGND.n20 4.65
R247 VGND.n24 VGND.n23 4.65
R248 VGND.n26 VGND.n25 4.65
R249 VGND.n29 VGND.n28 4.65
R250 VGND.n31 VGND.n30 4.65
R251 VGND.n33 VGND.n32 4.65
R252 VGND.n35 VGND.n34 4.65
R253 VGND.n37 VGND.n36 4.65
R254 VGND.n39 VGND.n38 4.65
R255 VGND.n43 VGND.n42 4.65
R256 VGND.n45 VGND.n44 4.65
R257 VGND.n47 VGND.n46 4.65
R258 VGND.n49 VGND.n48 4.65
R259 VGND.n51 VGND.n50 4.65
R260 VGND.n54 VGND.n53 4.65
R261 VGND.n56 VGND.n55 4.65
R262 VGND.n58 VGND.n57 4.65
R263 VGND.n60 VGND.n59 4.65
R264 VGND.n62 VGND.n61 4.65
R265 VGND.n64 VGND.n63 4.65
R266 VGND.n67 VGND.n66 3.932
R267 VGND.n23 VGND.n22 2.635
R268 VGND.n42 VGND.n41 0.752
R269 VGND.n4 VGND.n2 0.438
R270 VGND.n67 VGND.n64 0.137
R271 VGND VGND.n67 0.123
R272 VGND.n8 VGND.n4 0.119
R273 VGND.n10 VGND.n8 0.119
R274 VGND.n13 VGND.n10 0.119
R275 VGND.n15 VGND.n13 0.119
R276 VGND.n17 VGND.n15 0.119
R277 VGND.n19 VGND.n17 0.119
R278 VGND.n21 VGND.n19 0.119
R279 VGND.n24 VGND.n21 0.119
R280 VGND.n26 VGND.n24 0.119
R281 VGND.n29 VGND.n26 0.119
R282 VGND.n31 VGND.n29 0.119
R283 VGND.n33 VGND.n31 0.119
R284 VGND.n35 VGND.n33 0.119
R285 VGND.n37 VGND.n35 0.119
R286 VGND.n39 VGND.n37 0.119
R287 VGND.n43 VGND.n39 0.119
R288 VGND.n45 VGND.n43 0.119
R289 VGND.n47 VGND.n45 0.119
R290 VGND.n49 VGND.n47 0.119
R291 VGND.n51 VGND.n49 0.119
R292 VGND.n54 VGND.n51 0.119
R293 VGND.n56 VGND.n54 0.119
R294 VGND.n58 VGND.n56 0.119
R295 VGND.n60 VGND.n58 0.119
R296 VGND.n62 VGND.n60 0.119
R297 VGND.n64 VGND.n62 0.119
R298 a_1610_159.n1 a_1610_159.t2 406.399
R299 a_1610_159.n0 a_1610_159.t5 318.12
R300 a_1610_159.t0 a_1610_159.n3 262.563
R301 a_1610_159.n0 a_1610_159.t3 194.476
R302 a_1610_159.n1 a_1610_159.t4 130.052
R303 a_1610_159.n2 a_1610_159.n1 100.533
R304 a_1610_159.n2 a_1610_159.t1 93.987
R305 a_1610_159.n3 a_1610_159.n0 92.484
R306 a_1610_159.n3 a_1610_159.n2 9.323
R307 a_193_47.n1 a_193_47.t2 389.542
R308 a_193_47.n1 a_193_47.t5 273.571
R309 a_193_47.t0 a_193_47.n3 249.337
R310 a_193_47.n0 a_193_47.t4 232.651
R311 a_193_47.n0 a_193_47.t3 222.372
R312 a_193_47.n3 a_193_47.t1 207.871
R313 a_193_47.n2 a_193_47.n1 93.104
R314 a_193_47.n3 a_193_47.n2 9.98
R315 a_193_47.n2 a_193_47.n0 7.6
R316 a_1561_47.t0 a_1561_47.t1 111.393
R317 Q.n2 Q.n0 121.986
R318 Q.n4 Q.n3 121.986
R319 Q.n2 Q.n1 66.588
R320 Q Q.n5 63.679
R321 Q.n4 Q.n2 29.013
R322 Q.n3 Q.t1 26.595
R323 Q.n3 Q.t0 26.595
R324 Q.n0 Q.t3 26.595
R325 Q.n0 Q.t2 26.595
R326 Q.n5 Q.t7 24.923
R327 Q.n5 Q.t6 24.923
R328 Q.n1 Q.t4 24.923
R329 Q.n1 Q.t5 24.923
R330 Q Q.n4 2.909
R331 a_791_264.n2 a_791_264.t5 382.743
R332 a_791_264.n0 a_791_264.t2 310.621
R333 a_791_264.t0 a_791_264.n3 216.537
R334 a_791_264.n0 a_791_264.t3 194.941
R335 a_791_264.n1 a_791_264.t1 149.821
R336 a_791_264.n2 a_791_264.t4 138.53
R337 a_791_264.n1 a_791_264.n0 135.659
R338 a_791_264.n3 a_791_264.n2 98.016
R339 a_791_264.n3 a_791_264.n1 48.37
R340 a_1974_47.n0 a_1974_47.t1 70
R341 a_1974_47.n0 a_1974_47.t0 26.393
R342 a_1974_47.n1 a_1974_47.n0 14.4
R343 a_1231_369.t0 a_1231_369.t1 101.578
R344 a_915_47.t2 a_915_47.n5 305.929
R345 a_915_47.n2 a_915_47.n0 221.84
R346 a_915_47.n0 a_915_47.t3 117.17
R347 a_915_47.n4 a_915_47.n3 97.479
R348 a_915_47.n2 a_915_47.n1 92.5
R349 a_915_47.n3 a_915_47.t0 75.384
R350 a_915_47.n0 a_915_47.t5 61.587
R351 a_915_47.n5 a_915_47.t4 46.68
R352 a_915_47.n1 a_915_47.t1 32.197
R353 a_915_47.n4 a_915_47.n2 9.521
R354 a_915_47.n5 a_915_47.n4 7.415
R355 a_729_47.t0 a_729_47.t1 102.857
R356 a_729_369.t0 a_729_369.t1 110.812
R357 a_2135_413.t0 a_2135_413.t1 197
R358 SCD.n0 SCD.t1 206.188
R359 SCD.n0 SCD.t0 183.694
R360 SCD SCD.n0 87.674
R361 a_1226_119.t0 a_1226_119.t1 60
R362 a_1960_413.t0 a_1960_413.t1 143.059
R363 a_381_47.t0 a_381_47.t1 60
C0 VPB VGND 0.10fF
C1 VPWR Q 0.78fF
C2 D DE 0.13fF
C3 VGND Q 0.59fF
C4 VPB VPWR 0.32fF
C5 VPWR VGND 0.20fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__tap_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__tap_1 VGND VPWR VNB VPB
.ends

* NGSPICE file created from sky130_fd_sc_hd__tap_2.ext - technology: sky130A

.subckt sky130_fd_sc_hd__tap_2 VGND VPWR VPB VNB
C0 VPB VPWR 0.14fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__tapvgnd2_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__tapvgnd2_1 VPB VGND VPWR
.ends

* NGSPICE file created from sky130_fd_sc_hd__tapvgnd_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__tapvgnd_1 VPB VGND VPWR
C0 VPB VPWR 0.16fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__tapvpwrvgnd_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VPWR VGND
.ends

* NGSPICE file created from sky130_fd_sc_hd__xnor2_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__xnor2_1 VGND VPWR B Y A VNB VPB
X0 a_377_297.t1 A.t0 VPWR.t3 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_47_47.t0 B.t0 VPWR.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 a_129_47.t0 B.t1 a_47_47.t1 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 a_285_47.t1 B.t2 VGND.t0 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 Y.t1 a_47_47.t3 a_285_47.t0 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 VGND.t1 A.t1 a_129_47.t1 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 VPWR.t2 A.t2 a_47_47.t2 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 VPWR.t1 a_47_47.t4 Y.t0 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 Y.t2 B.t3 a_377_297.t0 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 a_285_47.t2 A.t3 VGND.t2 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
R0 A.n1 A.t0 266.851
R1 A.n2 A.t2 212.079
R2 A.n2 A.t1 139.779
R3 A.n0 A.t3 139.779
R4 A.n4 A.n1 97.76
R5 A.n4 A.n3 76
R6 A.n3 A.n2 24.1
R7 A.n1 A.n0 12.415
R8 A A.n4 1.92
R9 VPWR.n9 VPWR.t0 541.829
R10 VPWR.n2 VPWR.t1 481.98
R11 VPWR.n4 VPWR.n3 292.5
R12 VPWR.n1 VPWR.n0 292.5
R13 VPWR.n0 VPWR.t3 26.595
R14 VPWR.n3 VPWR.t2 26.595
R15 VPWR.n6 VPWR.n5 4.65
R16 VPWR.n8 VPWR.n7 4.65
R17 VPWR.n10 VPWR.n9 4.65
R18 VPWR.n2 VPWR.n1 4.264
R19 VPWR.n5 VPWR.n4 0.188
R20 VPWR.n6 VPWR.n2 0.144
R21 VPWR.n8 VPWR.n6 0.119
R22 VPWR.n10 VPWR.n8 0.119
R23 VPWR VPWR.n10 0.022
R24 a_377_297.t0 a_377_297.t1 41.37
R25 VPB.t3 VPB.t4 520.872
R26 VPB.t1 VPB.t2 284.112
R27 VPB.t0 VPB.t3 248.598
R28 VPB VPB.t0 216.043
R29 VPB.t4 VPB.t1 213.084
R30 B.n1 B.t0 241.534
R31 B.n0 B.t3 241.534
R32 B.n2 B.n0 208.515
R33 B.n1 B.t1 169.234
R34 B.n0 B.t2 169.234
R35 B B.n1 90.889
R36 B B.n2 4.894
R37 B.n2 B 4.44
R38 a_47_47.n1 a_47_47.n0 247.669
R39 a_47_47.n0 a_47_47.t4 241.534
R40 a_47_47.n1 a_47_47.t1 191.644
R41 a_47_47.n0 a_47_47.t3 169.234
R42 a_47_47.n2 a_47_47.n1 152.966
R43 a_47_47.n2 a_47_47.t2 26.595
R44 a_47_47.t0 a_47_47.n2 26.595
R45 a_129_47.t0 a_129_47.t1 38.769
R46 VNB VNB.t2 6561.6
R47 VNB.t3 VNB.t1 4545.05
R48 VNB.t1 VNB.t0 2030.77
R49 VNB.t4 VNB.t3 2030.77
R50 VNB.t2 VNB.t4 1740.66
R51 VGND.n1 VGND.t0 188.788
R52 VGND.n1 VGND.n0 79.097
R53 VGND.n0 VGND.t2 24.923
R54 VGND.n0 VGND.t1 24.923
R55 VGND VGND.n1 0.317
R56 a_285_47.n0 a_285_47.t2 242.797
R57 a_285_47.t0 a_285_47.n0 24.923
R58 a_285_47.n0 a_285_47.t1 24.923
R59 Y Y.n0 336.415
R60 Y Y.t1 214.91
R61 Y.n0 Y.t2 38.415
R62 Y.n0 Y.t0 26.595
C0 B A 0.36fF
C1 VPWR Y 0.16fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__xnor2_2.ext - technology: sky130A

.subckt sky130_fd_sc_hd__xnor2_2 VGND VPWR Y A B VNB VPB
X0 a_27_297.t5 B.t0 VPWR.t7 VPB.t7 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_560_47.t1 A.t0 VGND.t2 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 VGND.t5 B.t1 a_560_47.t3 VNB.t7 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 Y.t1 B.t2 a_474_297.t3 VPB.t6 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 VGND.t0 A.t1 a_27_47.t1 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 Y.t3 a_27_297.t6 a_560_47.t5 VNB.t9 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 a_474_297.t2 B.t3 Y.t0 VPB.t5 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 VGND.t1 A.t2 a_560_47.t0 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 a_27_47.t3 B.t4 a_27_297.t3 VNB.t6 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 a_27_297.t2 B.t5 a_27_47.t2 VNB.t5 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 a_27_47.t0 A.t3 VGND.t3 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 VPWR.t6 B.t6 a_27_297.t4 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 a_474_297.t1 A.t4 VPWR.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13 a_560_47.t4 a_27_297.t7 Y.t2 VNB.t8 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14 VPWR.t1 A.t5 a_474_297.t0 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 Y.t5 a_27_297.t8 VPWR.t4 VPB.t9 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16 VPWR.t5 a_27_297.t9 Y.t4 VPB.t8 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17 a_560_47.t2 B.t7 VGND.t4 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X18 a_27_297.t0 A.t6 VPWR.t2 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X19 VPWR.t3 A.t7 a_27_297.t1 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
R0 B B.n2 279.974
R1 B.n3 B.t0 212.079
R2 B.n4 B.t6 212.079
R3 B.n0 B.t3 212.079
R4 B.n1 B.t2 212.079
R5 B.n3 B.t4 139.779
R6 B.n4 B.t5 139.779
R7 B.n0 B.t1 139.779
R8 B.n1 B.t7 139.779
R9 B B.n5 116.066
R10 B.n2 B.n0 38.706
R11 B.n5 B.n3 37.245
R12 B.n2 B.n1 27.751
R13 B.n5 B.n4 24.1
R14 VPWR.n0 VPWR.t4 552.677
R15 VPWR.n9 VPWR.n8 314.004
R16 VPWR.n16 VPWR.n15 314.004
R17 VPWR.n21 VPWR.n20 314.004
R18 VPWR.n1 VPWR.t5 191.559
R19 VPWR.n8 VPWR.t0 26.595
R20 VPWR.n8 VPWR.t1 26.595
R21 VPWR.n15 VPWR.t2 26.595
R22 VPWR.n15 VPWR.t3 26.595
R23 VPWR.n20 VPWR.t7 26.595
R24 VPWR.n20 VPWR.t6 26.595
R25 VPWR.n3 VPWR.n2 4.65
R26 VPWR.n5 VPWR.n4 4.65
R27 VPWR.n7 VPWR.n6 4.65
R28 VPWR.n10 VPWR.n9 4.65
R29 VPWR.n12 VPWR.n11 4.65
R30 VPWR.n14 VPWR.n13 4.65
R31 VPWR.n17 VPWR.n16 4.65
R32 VPWR.n19 VPWR.n18 4.65
R33 VPWR.n22 VPWR.n21 4.017
R34 VPWR.n1 VPWR.n0 3.977
R35 VPWR.n3 VPWR.n1 0.248
R36 VPWR.n22 VPWR.n19 0.135
R37 VPWR VPWR.n22 0.125
R38 VPWR.n5 VPWR.n3 0.119
R39 VPWR.n7 VPWR.n5 0.119
R40 VPWR.n10 VPWR.n7 0.119
R41 VPWR.n12 VPWR.n10 0.119
R42 VPWR.n14 VPWR.n12 0.119
R43 VPWR.n17 VPWR.n14 0.119
R44 VPWR.n19 VPWR.n17 0.119
R45 a_27_297.n5 a_27_297.n4 333.759
R46 a_27_297.n2 a_27_297.t9 212.079
R47 a_27_297.n3 a_27_297.t8 212.079
R48 a_27_297.n5 a_27_297.t0 181.424
R49 a_27_297.n1 a_27_297.t4 179.673
R50 a_27_297.n1 a_27_297.n0 171.031
R51 a_27_297.n7 a_27_297.n6 154.828
R52 a_27_297.n2 a_27_297.t6 139.779
R53 a_27_297.n3 a_27_297.t7 139.779
R54 a_27_297.n6 a_27_297.n1 41.955
R55 a_27_297.n6 a_27_297.n5 41.955
R56 a_27_297.n4 a_27_297.n2 36.515
R57 a_27_297.n7 a_27_297.t1 26.595
R58 a_27_297.t5 a_27_297.n7 26.595
R59 a_27_297.n0 a_27_297.t3 24.923
R60 a_27_297.n0 a_27_297.t2 24.923
R61 a_27_297.n4 a_27_297.n3 24.83
R62 VPB.t2 VPB.t1 580.062
R63 VPB.t5 VPB.t9 556.386
R64 VPB.t6 VPB.t5 269.314
R65 VPB.t9 VPB.t8 248.598
R66 VPB.t0 VPB.t6 248.598
R67 VPB.t1 VPB.t0 248.598
R68 VPB.t3 VPB.t2 248.598
R69 VPB.t7 VPB.t3 248.598
R70 VPB.t4 VPB.t7 248.598
R71 VPB VPB.t4 201.246
R72 A.n0 A.t4 212.079
R73 A.n1 A.t5 212.079
R74 A.n5 A.t6 212.079
R75 A.n3 A.t7 212.079
R76 A.n0 A.t2 139.779
R77 A.n1 A.t0 139.779
R78 A.n5 A.t3 139.779
R79 A.n3 A.t1 139.779
R80 A.n7 A.n4 97.76
R81 A.n7 A.n6 76
R82 A.n2 A.n1 61.586
R83 A.n1 A.n0 61.345
R84 A A.n2 40.429
R85 A A.n7 14.4
R86 A.n4 A.n3 13.875
R87 A.n6 A.n5 2.19
R88 VGND.n2 VGND.t5 203.574
R89 VGND.n1 VGND.n0 115.464
R90 VGND.n11 VGND.n10 115.464
R91 VGND.n5 VGND.t2 111.584
R92 VGND.n0 VGND.t4 24.923
R93 VGND.n0 VGND.t1 24.923
R94 VGND.n10 VGND.t3 24.923
R95 VGND.n10 VGND.t0 24.923
R96 VGND.n2 VGND.n1 11.125
R97 VGND.n12 VGND.n11 5.647
R98 VGND.n4 VGND.n3 4.65
R99 VGND.n7 VGND.n6 4.65
R100 VGND.n9 VGND.n8 4.65
R101 VGND.n13 VGND.n12 4.65
R102 VGND.n6 VGND.n5 1.129
R103 VGND.n4 VGND.n2 0.301
R104 VGND VGND.n14 0.247
R105 VGND.n14 VGND.n13 0.134
R106 VGND.n7 VGND.n4 0.119
R107 VGND.n9 VGND.n7 0.119
R108 VGND.n13 VGND.n9 0.119
R109 a_560_47.n2 a_560_47.n0 173.867
R110 a_560_47.n3 a_560_47.n2 88.889
R111 a_560_47.n2 a_560_47.n1 52.031
R112 a_560_47.n1 a_560_47.t2 31.384
R113 a_560_47.n0 a_560_47.t5 24.923
R114 a_560_47.n0 a_560_47.t4 24.923
R115 a_560_47.n1 a_560_47.t3 24.923
R116 a_560_47.n3 a_560_47.t0 24.923
R117 a_560_47.t1 a_560_47.n3 24.923
R118 VNB VNB.t5 6150.61
R119 VNB.t0 VNB.t3 4738.46
R120 VNB.t7 VNB.t8 4545.05
R121 VNB.t4 VNB.t7 2200
R122 VNB.t8 VNB.t9 2030.77
R123 VNB.t1 VNB.t4 2030.77
R124 VNB.t3 VNB.t1 2030.77
R125 VNB.t2 VNB.t0 2030.77
R126 VNB.t6 VNB.t2 2030.77
R127 VNB.t5 VNB.t6 2030.77
R128 a_474_297.n0 a_474_297.t2 580.787
R129 a_474_297.n0 a_474_297.t0 204.237
R130 a_474_297.t1 a_474_297.n1 36.097
R131 a_474_297.n1 a_474_297.t3 16.306
R132 a_474_297.n1 a_474_297.n0 9.963
R133 Y.n2 Y.n0 387.479
R134 Y.n3 Y.t2 233.211
R135 Y.n2 Y.n1 144.013
R136 Y.n3 Y.t3 82.78
R137 Y.n0 Y.t1 33.49
R138 Y Y.n3 28.869
R139 Y Y.n2 26.845
R140 Y.n1 Y.t4 26.595
R141 Y.n1 Y.t5 26.595
R142 Y.n0 Y.t0 26.595
R143 a_27_47.n0 a_27_47.t2 219.844
R144 a_27_47.n0 a_27_47.t0 137.72
R145 a_27_47.n1 a_27_47.n0 42.273
R146 a_27_47.t1 a_27_47.n1 24.923
R147 a_27_47.n1 a_27_47.t3 24.923
C0 VPWR VGND 0.11fF
C1 Y VGND 0.20fF
C2 VPB VPWR 0.12fF
C3 B A 0.53fF
C4 VPWR Y 0.24fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__xnor2_4.ext - technology: sky130A

.subckt sky130_fd_sc_hd__xnor2_4 Y B A VGND VPWR VNB VPB
X0 VGND.t11 A.t0 a_902_47.t11 VNB.t19 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 Y.t7 a_38_297.t12 VPWR.t7 VPB.t11 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 a_38_297.t0 B.t0 VPWR.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 a_820_297.t3 B.t1 Y.t0 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 VPWR.t6 a_38_297.t13 Y.t6 VPB.t10 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 VGND.t10 A.t1 a_902_47.t10 VNB.t18 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 VGND.t0 B.t2 a_902_47.t0 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 VGND.t1 B.t3 a_902_47.t1 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 Y.t1 B.t4 a_820_297.t2 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 a_38_297.t11 A.t2 VPWR.t15 VPB.t19 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 a_38_297.t1 B.t5 a_38_47.t3 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 VGND.t7 A.t3 a_38_47.t7 VNB.t17 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 a_902_47.t2 B.t6 VGND.t2 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 a_820_297.t1 B.t7 Y.t2 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14 a_902_47.t3 B.t8 VGND.t3 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X15 VPWR.t14 A.t4 a_38_297.t10 VPB.t18 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16 Y.t11 a_38_297.t14 a_902_47.t4 VNB.t8 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X17 Y.t10 a_38_297.t15 a_902_47.t5 VNB.t9 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X18 a_38_47.t2 B.t9 a_38_297.t2 VNB.t5 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X19 a_38_47.t1 B.t10 a_38_297.t3 VNB.t6 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X20 a_38_297.t4 B.t11 a_38_47.t0 VNB.t7 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X21 a_38_47.t6 A.t5 VGND.t6 VNB.t16 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X22 VPWR.t1 B.t12 a_38_297.t5 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X23 a_38_47.t5 A.t6 VGND.t5 VNB.t15 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X24 a_902_47.t6 a_38_297.t16 Y.t9 VNB.t10 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X25 a_902_47.t7 a_38_297.t17 Y.t8 VNB.t11 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X26 Y.t3 B.t13 a_820_297.t0 VPB.t5 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X27 a_38_297.t9 A.t7 VPWR.t13 VPB.t17 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X28 a_820_297.t7 A.t8 VPWR.t11 VPB.t16 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X29 VPWR.t12 A.t9 a_38_297.t8 VPB.t15 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X30 VGND.t4 A.t10 a_38_47.t4 VNB.t14 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X31 VPWR.t10 A.t11 a_820_297.t6 VPB.t14 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X32 a_902_47.t9 A.t12 VGND.t9 VNB.t13 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X33 a_820_297.t5 A.t13 VPWR.t9 VPB.t13 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X34 Y.t5 a_38_297.t18 VPWR.t5 VPB.t9 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X35 a_902_47.t8 A.t14 VGND.t8 VNB.t12 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X36 a_38_297.t6 B.t14 VPWR.t2 VPB.t6 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X37 VPWR.t8 A.t15 a_820_297.t4 VPB.t12 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X38 VPWR.t4 a_38_297.t19 Y.t4 VPB.t8 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X39 VPWR.t3 B.t15 a_38_297.t7 VPB.t7 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
R0 A.n7 A.t2 212.079
R1 A.n14 A.t4 212.079
R2 A.n11 A.t7 212.079
R3 A.n9 A.t9 212.079
R4 A.n0 A.t8 212.079
R5 A.n1 A.t11 212.079
R6 A.n2 A.t13 212.079
R7 A.n4 A.t15 212.079
R8 A.n7 A.t6 139.779
R9 A.n14 A.t10 139.779
R10 A.n11 A.t5 139.779
R11 A.n9 A.t3 139.779
R12 A.n0 A.t0 139.779
R13 A.n1 A.t12 139.779
R14 A.n2 A.t1 139.779
R15 A.n4 A.t14 139.779
R16 A.n13 A.n10 97.76
R17 A.n6 A.n5 76
R18 A.n17 A.n8 76
R19 A.n16 A.n15 76
R20 A.n13 A.n12 76
R21 A.n1 A.n0 61.345
R22 A.n6 A.n3 55.015
R23 A A.n6 46.08
R24 A A.n17 29.12
R25 A.n3 A.n1 29.033
R26 A.n17 A.n16 21.76
R27 A.n16 A.n13 21.76
R28 A.n3 A.n2 21.274
R29 A.n10 A.n9 18.257
R30 A.n8 A.n7 16.796
R31 A.n5 A.n4 16.066
R32 A.n12 A.n11 6.572
R33 A.n15 A.n14 5.112
R34 a_902_47.n4 a_902_47.t7 228.604
R35 a_902_47.n4 a_902_47.n3 92.5
R36 a_902_47.n2 a_902_47.n0 88.89
R37 a_902_47.n5 a_902_47.t4 81.34
R38 a_902_47.n5 a_902_47.n4 65.13
R39 a_902_47.n7 a_902_47.n5 59.907
R40 a_902_47.n7 a_902_47.n6 52.624
R41 a_902_47.n2 a_902_47.n1 52.624
R42 a_902_47.n9 a_902_47.n8 52.623
R43 a_902_47.n8 a_902_47.n2 36.266
R44 a_902_47.n8 a_902_47.n7 36.266
R45 a_902_47.n3 a_902_47.t5 24.923
R46 a_902_47.n3 a_902_47.t6 24.923
R47 a_902_47.n6 a_902_47.t1 24.923
R48 a_902_47.n6 a_902_47.t3 24.923
R49 a_902_47.n0 a_902_47.t10 24.923
R50 a_902_47.n0 a_902_47.t8 24.923
R51 a_902_47.n1 a_902_47.t11 24.923
R52 a_902_47.n1 a_902_47.t9 24.923
R53 a_902_47.t0 a_902_47.n9 24.923
R54 a_902_47.n9 a_902_47.t2 24.923
R55 VGND.n0 VGND.t1 192.535
R56 VGND.n2 VGND.n1 115.464
R57 VGND.n8 VGND.n7 115.464
R58 VGND.n12 VGND.n11 115.464
R59 VGND.n23 VGND.n22 115.464
R60 VGND.n29 VGND.n28 115.464
R61 VGND.n17 VGND.t8 107.415
R62 VGND.n1 VGND.t3 24.923
R63 VGND.n1 VGND.t0 24.923
R64 VGND.n7 VGND.t2 24.923
R65 VGND.n7 VGND.t11 24.923
R66 VGND.n11 VGND.t9 24.923
R67 VGND.n11 VGND.t10 24.923
R68 VGND.n22 VGND.t5 24.923
R69 VGND.n22 VGND.t4 24.923
R70 VGND.n28 VGND.t6 24.923
R71 VGND.n28 VGND.t7 24.923
R72 VGND.n13 VGND.n12 16.941
R73 VGND.n24 VGND.n23 13.176
R74 VGND.n9 VGND.n8 11.67
R75 VGND.n30 VGND.n29 7.152
R76 VGND.n3 VGND.n2 5.647
R77 VGND.n4 VGND.n3 4.65
R78 VGND.n6 VGND.n5 4.65
R79 VGND.n10 VGND.n9 4.65
R80 VGND.n14 VGND.n13 4.65
R81 VGND.n16 VGND.n15 4.65
R82 VGND.n19 VGND.n18 4.65
R83 VGND.n21 VGND.n20 4.65
R84 VGND.n25 VGND.n24 4.65
R85 VGND.n27 VGND.n26 4.65
R86 VGND.n31 VGND.n30 4.65
R87 VGND.n18 VGND.n17 4.517
R88 VGND.n4 VGND.n0 0.635
R89 VGND VGND.n32 0.486
R90 VGND.n32 VGND.n31 0.134
R91 VGND.n6 VGND.n4 0.119
R92 VGND.n10 VGND.n6 0.119
R93 VGND.n14 VGND.n10 0.119
R94 VGND.n16 VGND.n14 0.119
R95 VGND.n19 VGND.n16 0.119
R96 VGND.n21 VGND.n19 0.119
R97 VGND.n25 VGND.n21 0.119
R98 VGND.n27 VGND.n25 0.119
R99 VGND.n31 VGND.n27 0.119
R100 VNB VNB.t7 6440.72
R101 VNB.t1 VNB.t8 4641.76
R102 VNB.t15 VNB.t12 4593.41
R103 VNB.t9 VNB.t11 2030.77
R104 VNB.t10 VNB.t9 2030.77
R105 VNB.t8 VNB.t10 2030.77
R106 VNB.t4 VNB.t1 2030.77
R107 VNB.t0 VNB.t4 2030.77
R108 VNB.t3 VNB.t0 2030.77
R109 VNB.t19 VNB.t3 2030.77
R110 VNB.t13 VNB.t19 2030.77
R111 VNB.t18 VNB.t13 2030.77
R112 VNB.t12 VNB.t18 2030.77
R113 VNB.t14 VNB.t15 2030.77
R114 VNB.t16 VNB.t14 2030.77
R115 VNB.t17 VNB.t16 2030.77
R116 VNB.t6 VNB.t17 2030.77
R117 VNB.t2 VNB.t6 2030.77
R118 VNB.t5 VNB.t2 2030.77
R119 VNB.t7 VNB.t5 2030.77
R120 a_38_297.n3 a_38_297.t11 214.727
R121 a_38_297.n11 a_38_297.t18 212.079
R122 a_38_297.n13 a_38_297.t19 212.079
R123 a_38_297.n16 a_38_297.t12 212.079
R124 a_38_297.n19 a_38_297.t13 212.079
R125 a_38_297.n22 a_38_297.n21 183.534
R126 a_38_297.n3 a_38_297.n2 153.805
R127 a_38_297.n5 a_38_297.n4 153.805
R128 a_38_297.n11 a_38_297.t17 139.779
R129 a_38_297.n13 a_38_297.t15 139.779
R130 a_38_297.n16 a_38_297.t16 139.779
R131 a_38_297.n19 a_38_297.t14 139.779
R132 a_38_297.n9 a_38_297.n7 133.853
R133 a_38_297.n10 a_38_297.t5 133.386
R134 a_38_297.n15 a_38_297.n12 97.76
R135 a_38_297.n9 a_38_297.n8 92.5
R136 a_38_297.n21 a_38_297.n20 76
R137 a_38_297.n15 a_38_297.n14 76
R138 a_38_297.n18 a_38_297.n17 76
R139 a_38_297.n10 a_38_297.n9 59.636
R140 a_38_297.n22 a_38_297.n10 45.399
R141 a_38_297.n6 a_38_297.n5 38.703
R142 a_38_297.n5 a_38_297.n3 34.327
R143 a_38_297.n2 a_38_297.t10 26.595
R144 a_38_297.n2 a_38_297.t9 26.595
R145 a_38_297.n4 a_38_297.t8 26.595
R146 a_38_297.n4 a_38_297.t6 26.595
R147 a_38_297.n7 a_38_297.t3 24.923
R148 a_38_297.n7 a_38_297.t1 24.923
R149 a_38_297.n8 a_38_297.t2 24.923
R150 a_38_297.n8 a_38_297.t4 24.923
R151 a_38_297.t0 a_38_297.n24 23.64
R152 a_38_297.n18 a_38_297.n15 21.76
R153 a_38_297.n21 a_38_297.n18 21.76
R154 a_38_297.n12 a_38_297.n11 18.987
R155 a_38_297.n20 a_38_297.n19 16.066
R156 a_38_297.n1 a_38_297.n0 13.79
R157 a_38_297.n0 a_38_297.t7 12.805
R158 a_38_297.n23 a_38_297.n6 11.635
R159 a_38_297.n24 a_38_297.n23 9.3
R160 a_38_297.n14 a_38_297.n13 7.303
R161 a_38_297.n17 a_38_297.n16 4.381
R162 a_38_297.n24 a_38_297.n1 2.955
R163 a_38_297.n23 a_38_297.n22 0.889
R164 VPWR.n17 VPWR.n16 311.956
R165 VPWR.n21 VPWR.n20 311.956
R166 VPWR.n29 VPWR.n28 311.956
R167 VPWR.n35 VPWR.n34 311.956
R168 VPWR.n40 VPWR.n39 311.956
R169 VPWR.n3 VPWR.n2 173.549
R170 VPWR.n45 VPWR.n44 169.933
R171 VPWR.n1 VPWR.n0 169.933
R172 VPWR.n2 VPWR.t5 26.595
R173 VPWR.n2 VPWR.t4 26.595
R174 VPWR.n0 VPWR.t7 26.595
R175 VPWR.n0 VPWR.t6 26.595
R176 VPWR.n16 VPWR.t11 26.595
R177 VPWR.n16 VPWR.t10 26.595
R178 VPWR.n20 VPWR.t9 26.595
R179 VPWR.n20 VPWR.t8 26.595
R180 VPWR.n28 VPWR.t15 26.595
R181 VPWR.n28 VPWR.t14 26.595
R182 VPWR.n34 VPWR.t13 26.595
R183 VPWR.n34 VPWR.t12 26.595
R184 VPWR.n39 VPWR.t2 26.595
R185 VPWR.n39 VPWR.t3 26.595
R186 VPWR.n44 VPWR.t0 26.595
R187 VPWR.n44 VPWR.t1 26.595
R188 VPWR.n18 VPWR.n17 5.27
R189 VPWR.n5 VPWR.n4 4.65
R190 VPWR.n7 VPWR.n6 4.65
R191 VPWR.n9 VPWR.n8 4.65
R192 VPWR.n11 VPWR.n10 4.65
R193 VPWR.n13 VPWR.n12 4.65
R194 VPWR.n15 VPWR.n14 4.65
R195 VPWR.n19 VPWR.n18 4.65
R196 VPWR.n23 VPWR.n22 4.65
R197 VPWR.n25 VPWR.n24 4.65
R198 VPWR.n27 VPWR.n26 4.65
R199 VPWR.n31 VPWR.n30 4.65
R200 VPWR.n33 VPWR.n32 4.65
R201 VPWR.n36 VPWR.n35 4.65
R202 VPWR.n38 VPWR.n37 4.65
R203 VPWR.n41 VPWR.n40 4.65
R204 VPWR.n43 VPWR.n42 4.65
R205 VPWR.n22 VPWR.n21 4.517
R206 VPWR.n46 VPWR.n45 4.09
R207 VPWR.n3 VPWR.n1 3.847
R208 VPWR.n30 VPWR.n29 3.764
R209 VPWR.n5 VPWR.n3 0.232
R210 VPWR.n46 VPWR.n43 0.133
R211 VPWR VPWR.n46 0.127
R212 VPWR.n7 VPWR.n5 0.119
R213 VPWR.n9 VPWR.n7 0.119
R214 VPWR.n11 VPWR.n9 0.119
R215 VPWR.n13 VPWR.n11 0.119
R216 VPWR.n15 VPWR.n13 0.119
R217 VPWR.n19 VPWR.n15 0.119
R218 VPWR.n23 VPWR.n19 0.119
R219 VPWR.n25 VPWR.n23 0.119
R220 VPWR.n27 VPWR.n25 0.119
R221 VPWR.n31 VPWR.n27 0.119
R222 VPWR.n33 VPWR.n31 0.119
R223 VPWR.n36 VPWR.n33 0.119
R224 VPWR.n38 VPWR.n36 0.119
R225 VPWR.n41 VPWR.n38 0.119
R226 VPWR.n43 VPWR.n41 0.119
R227 Y.n2 Y.n1 333.853
R228 Y.n2 Y.n0 292.5
R229 Y.n8 Y.n7 133.853
R230 Y.n10 Y.t5 126.817
R231 Y.n3 Y.t6 123.727
R232 Y.n5 Y.n4 109.992
R233 Y.n8 Y.n6 92.5
R234 Y.n9 Y.n8 61.968
R235 Y.n5 Y.n3 45.521
R236 Y.n3 Y.n2 43.462
R237 Y.n9 Y.n5 34.327
R238 Y.n1 Y.t2 26.595
R239 Y.n1 Y.t3 26.595
R240 Y.n0 Y.t0 26.595
R241 Y.n0 Y.t1 26.595
R242 Y.n4 Y.t4 26.595
R243 Y.n4 Y.t7 26.595
R244 Y.n6 Y.t8 24.923
R245 Y.n6 Y.t10 24.923
R246 Y.n7 Y.t9 24.923
R247 Y.n7 Y.t11 24.923
R248 Y.n10 Y.n9 6.176
R249 Y Y.n10 2.039
R250 VPB.t1 VPB.t10 568.224
R251 VPB.t19 VPB.t12 562.305
R252 VPB.t8 VPB.t9 248.598
R253 VPB.t11 VPB.t8 248.598
R254 VPB.t10 VPB.t11 248.598
R255 VPB.t2 VPB.t1 248.598
R256 VPB.t3 VPB.t2 248.598
R257 VPB.t5 VPB.t3 248.598
R258 VPB.t16 VPB.t5 248.598
R259 VPB.t14 VPB.t16 248.598
R260 VPB.t13 VPB.t14 248.598
R261 VPB.t12 VPB.t13 248.598
R262 VPB.t18 VPB.t19 248.598
R263 VPB.t17 VPB.t18 248.598
R264 VPB.t15 VPB.t17 248.598
R265 VPB.t6 VPB.t15 248.598
R266 VPB.t7 VPB.t6 248.598
R267 VPB.t0 VPB.t7 248.598
R268 VPB.t4 VPB.t0 248.598
R269 VPB VPB.t4 236.76
R270 B.n13 B.n10 361.524
R271 B.n11 B.t14 212.079
R272 B.n14 B.t15 212.079
R273 B.n19 B.t0 212.079
R274 B.n17 B.t12 212.079
R275 B.n0 B.t1 212.079
R276 B.n2 B.t4 212.079
R277 B.n5 B.t7 212.079
R278 B.n8 B.t13 212.079
R279 B.n11 B.t10 139.779
R280 B.n14 B.t5 139.779
R281 B.n19 B.t9 139.779
R282 B.n17 B.t11 139.779
R283 B.n0 B.t3 139.779
R284 B.n2 B.t8 139.779
R285 B.n5 B.t2 139.779
R286 B.n8 B.t6 139.779
R287 B.n4 B.n1 97.76
R288 B.n21 B.n18 97.76
R289 B.n10 B.n9 76
R290 B.n4 B.n3 76
R291 B.n7 B.n6 76
R292 B.n13 B.n12 76
R293 B.n16 B.n15 76
R294 B.n21 B.n20 76
R295 B.n7 B.n4 21.76
R296 B.n10 B.n7 21.76
R297 B.n16 B.n13 21.76
R298 B.n12 B.n11 18.987
R299 B.n9 B.n8 18.257
R300 B B.n16 17.28
R301 B.n1 B.n0 16.796
R302 B.n18 B.n17 16.066
R303 B.n15 B.n14 7.303
R304 B.n6 B.n5 6.572
R305 B.n3 B.n2 5.112
R306 B B.n21 4.48
R307 B.n20 B.n19 4.381
R308 a_820_297.t3 a_820_297.n5 574.181
R309 a_820_297.n5 a_820_297.n0 292.5
R310 a_820_297.n2 a_820_297.t4 213.188
R311 a_820_297.n2 a_820_297.n1 153.805
R312 a_820_297.n4 a_820_297.n3 143.164
R313 a_820_297.n5 a_820_297.n4 49.748
R314 a_820_297.n4 a_820_297.n2 47.203
R315 a_820_297.n0 a_820_297.t2 26.595
R316 a_820_297.n0 a_820_297.t1 26.595
R317 a_820_297.n3 a_820_297.t0 26.595
R318 a_820_297.n3 a_820_297.t7 26.595
R319 a_820_297.n1 a_820_297.t6 26.595
R320 a_820_297.n1 a_820_297.t5 26.595
R321 a_38_47.n4 a_38_47.t0 214.229
R322 a_38_47.n1 a_38_47.t5 128.218
R323 a_38_47.n5 a_38_47.n4 92.5
R324 a_38_47.n4 a_38_47.n3 53.163
R325 a_38_47.n1 a_38_47.n0 52.624
R326 a_38_47.n3 a_38_47.n1 48.574
R327 a_38_47.n3 a_38_47.n2 42.273
R328 a_38_47.n2 a_38_47.t7 24.923
R329 a_38_47.n2 a_38_47.t1 24.923
R330 a_38_47.n0 a_38_47.t4 24.923
R331 a_38_47.n0 a_38_47.t6 24.923
R332 a_38_47.t3 a_38_47.n5 24.923
R333 a_38_47.n5 a_38_47.t2 24.923
C0 VPB B 0.12fF
C1 VPWR VGND 0.12fF
C2 B A 0.99fF
C3 VPB VPWR 0.19fF
C4 A VGND 0.12fF
C5 VPWR Y 0.65fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__xnor3_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__xnor3_1 X B C A VGND VPWR VNB VPB
X0 a_841_297.t1 a_735_297.t2 a_355_49.t1 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=600000u l=150000u
X1 a_1106_49.t5 a_841_297.t6 VGND.t4 VNB.t10 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X2 a_78_199.t3 C.t0 a_355_49.t4 VNB.t8 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X3 a_1106_49.t1 a_735_297.t3 a_355_49.t0 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X4 a_735_297.t0 B.t0 VGND.t1 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 a_1106_49.t4 a_841_297.t7 VPWR.t1 VPB.t7 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 VPWR.t0 A.t0 a_841_297.t5 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 a_331_325.t4 B.t1 a_841_297.t3 VNB.t5 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X8 a_355_49.t3 B.t2 a_841_297.t4 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X9 a_216_93.t1 C.t1 VPWR.t4 VPB.t10 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X10 a_735_297.t1 B.t3 VPWR.t3 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 VPWR.t2 a_78_199.t4 X.t1 VPB.t8 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 a_355_49.t2 B.t4 a_1106_49.t2 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X13 a_331_325.t3 B.t5 a_1106_49.t3 VPB.t6 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X14 a_331_325.t2 a_216_93.t2 a_78_199.t0 VNB.t9 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X15 a_78_199.t2 C.t2 a_331_325.t5 VPB.t9 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X16 a_355_49.t5 a_216_93.t3 a_78_199.t1 VPB.t5 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X17 VGND.t0 A.t1 a_841_297.t2 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X18 a_216_93.t0 C.t3 VGND.t3 VNB.t7 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19 a_1106_49.t0 a_735_297.t4 a_331_325.t0 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20 a_841_297.t0 a_735_297.t5 a_331_325.t1 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X21 VGND.t2 a_78_199.t5 X.t0 VNB.t6 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
R0 a_735_297.t1 a_735_297.n3 599.237
R1 a_735_297.n0 a_735_297.t5 283.255
R2 a_735_297.n1 a_735_297.t4 173.52
R3 a_735_297.n0 a_735_297.t2 161.201
R4 a_735_297.n1 a_735_297.t3 154.239
R5 a_735_297.n2 a_735_297.n1 143.387
R6 a_735_297.n2 a_735_297.n0 94.522
R7 a_735_297.n3 a_735_297.t0 94.135
R8 a_735_297.n3 a_735_297.n2 2.703
R9 a_355_49.n1 a_355_49.t4 287.572
R10 a_355_49.n2 a_355_49.n0 250.115
R11 a_355_49.n1 a_355_49.t5 176.167
R12 a_355_49.n3 a_355_49.n2 151.6
R13 a_355_49.n3 a_355_49.t0 83.109
R14 a_355_49.n0 a_355_49.t1 51.386
R15 a_355_49.n4 a_355_49.t3 40.516
R16 a_355_49.n5 a_355_49.n4 39.797
R17 a_355_49.n4 a_355_49.n3 27.703
R18 a_355_49.n0 a_355_49.t2 25.321
R19 a_355_49.n2 a_355_49.n1 8.28
R20 a_841_297.n5 a_841_297.t4 468.615
R21 a_841_297.n9 a_841_297.n8 349.224
R22 a_841_297.n1 a_841_297.t7 241.534
R23 a_841_297.n1 a_841_297.t6 170.841
R24 a_841_297.n8 a_841_297.n1 76
R25 a_841_297.n8 a_841_297.n7 55.794
R26 a_841_297.n5 a_841_297.t3 52.25
R27 a_841_297.n0 a_841_297.t0 50.422
R28 a_841_297.n4 a_841_297.t1 42
R29 a_841_297.n10 a_841_297.n9 38.696
R30 a_841_297.n0 a_841_297.t5 28.87
R31 a_841_297.n9 a_841_297.n0 17.589
R32 a_841_297.n3 a_841_297.n2 13.805
R33 a_841_297.n6 a_841_297.n4 9.3
R34 a_841_297.n2 a_841_297.t2 9.275
R35 a_841_297.n6 a_841_297.n5 7.566
R36 a_841_297.n7 a_841_297.n6 3.71
R37 a_841_297.n4 a_841_297.n3 1
R38 VNB VNB.t6 6078.09
R39 VNB.t9 VNB.t3 5888.96
R40 VNB.t7 VNB.t8 5451.11
R41 VNB.t3 VNB.t5 4522.22
R42 VNB.t0 VNB.t4 3886.67
R43 VNB.t5 VNB.t0 3691.11
R44 VNB.t4 VNB.t1 2836.76
R45 VNB.t6 VNB.t7 2538.73
R46 VNB.t1 VNB.t2 2444.44
R47 VNB.t8 VNB.t9 2151.11
R48 VNB.t2 VNB.t10 2053.33
R49 VGND.n16 VGND.n15 151.577
R50 VGND.n1 VGND.n0 122.581
R51 VGND.n2 VGND.t1 108.528
R52 VGND.n15 VGND.t3 65.714
R53 VGND.n0 VGND.t4 25.312
R54 VGND.n0 VGND.t0 25.312
R55 VGND.n15 VGND.t2 20.091
R56 VGND.n3 VGND.n2 8.282
R57 VGND.n4 VGND.n3 4.65
R58 VGND.n6 VGND.n5 4.65
R59 VGND.n8 VGND.n7 4.65
R60 VGND.n10 VGND.n9 4.65
R61 VGND.n12 VGND.n11 4.65
R62 VGND.n14 VGND.n13 4.65
R63 VGND.n17 VGND.n16 3.932
R64 VGND.n17 VGND.n14 0.137
R65 VGND.n4 VGND.n1 0.134
R66 VGND VGND.n17 0.123
R67 VGND.n6 VGND.n4 0.119
R68 VGND.n8 VGND.n6 0.119
R69 VGND.n10 VGND.n8 0.119
R70 VGND.n12 VGND.n10 0.119
R71 VGND.n14 VGND.n12 0.119
R72 a_1106_49.n2 a_1106_49.n0 297.655
R73 a_1106_49.n3 a_1106_49.t5 226.304
R74 a_1106_49.n0 a_1106_49.t1 209.825
R75 a_1106_49.n2 a_1106_49.n1 192.264
R76 a_1106_49.t4 a_1106_49.n3 176.793
R77 a_1106_49.n3 a_1106_49.n2 130.955
R78 a_1106_49.n1 a_1106_49.t0 94.776
R79 a_1106_49.n0 a_1106_49.t3 41.555
R80 a_1106_49.n1 a_1106_49.t2 38.437
R81 C.n0 C.t2 269.92
R82 C.n1 C.t1 154.239
R83 C.n0 C.t0 143.284
R84 C.n2 C.n1 132.915
R85 C.n1 C.t3 102.826
R86 C C.n2 79.584
R87 C.n2 C.n0 24.83
R88 a_78_199.n3 a_78_199.n2 482.376
R89 a_78_199.n2 a_78_199.n1 258.911
R90 a_78_199.n0 a_78_199.t4 236.179
R91 a_78_199.n0 a_78_199.t5 163.879
R92 a_78_199.n2 a_78_199.n0 76
R93 a_78_199.n5 a_78_199.n4 55.16
R94 a_78_199.n3 a_78_199.t2 32.611
R95 a_78_199.n4 a_78_199.t1 30.341
R96 a_78_199.n1 a_78_199.t0 27.187
R97 a_78_199.n1 a_78_199.t3 27.187
R98 a_78_199.n4 a_78_199.n3 21.107
R99 VPB.t2 VPB.t3 651.09
R100 VPB.t5 VPB.t2 627.414
R101 VPB.t10 VPB.t9 621.495
R102 VPB.t1 VPB.t6 517.912
R103 VPB.t3 VPB.t1 446.884
R104 VPB.t6 VPB.t0 304.828
R105 VPB.t8 VPB.t10 304.828
R106 VPB.t0 VPB.t4 298.909
R107 VPB.t9 VPB.t5 287.071
R108 VPB.t4 VPB.t7 248.598
R109 VPB VPB.t8 204.205
R110 B.t5 B.t2 864.385
R111 B.n1 B.n0 298.84
R112 B.n0 B.t3 295.625
R113 B.n2 B.t5 235.107
R114 B.t2 B.n1 215.293
R115 B.n0 B.t0 168.699
R116 B.n2 B.t4 167.627
R117 B.n1 B.t1 167.092
R118 B B.n2 118.163
R119 VPWR.n0 VPWR.t3 490.559
R120 VPWR.n14 VPWR.n13 427.426
R121 VPWR.n2 VPWR.n1 310.72
R122 VPWR.n13 VPWR.t4 67.718
R123 VPWR.n13 VPWR.t2 30.376
R124 VPWR.n1 VPWR.t1 26.595
R125 VPWR.n1 VPWR.t0 26.595
R126 VPWR.n4 VPWR.n3 4.65
R127 VPWR.n6 VPWR.n5 4.65
R128 VPWR.n8 VPWR.n7 4.65
R129 VPWR.n10 VPWR.n9 4.65
R130 VPWR.n12 VPWR.n11 4.65
R131 VPWR.n2 VPWR.n0 4.027
R132 VPWR.n15 VPWR.n14 3.966
R133 VPWR.n4 VPWR.n2 0.137
R134 VPWR.n15 VPWR.n12 0.137
R135 VPWR VPWR.n15 0.124
R136 VPWR.n6 VPWR.n4 0.119
R137 VPWR.n8 VPWR.n6 0.119
R138 VPWR.n10 VPWR.n8 0.119
R139 VPWR.n12 VPWR.n10 0.119
R140 A.n0 A.t0 239.503
R141 A.n0 A.t1 168.81
R142 A A.n0 87.52
R143 a_331_325.n3 a_331_325.n2 490.648
R144 a_331_325.n1 a_331_325.t5 435.971
R145 a_331_325.n1 a_331_325.t2 262.941
R146 a_331_325.n2 a_331_325.n0 221.036
R147 a_331_325.n2 a_331_325.n1 116.704
R148 a_331_325.n0 a_331_325.t0 98.437
R149 a_331_325.n3 a_331_325.t3 67.718
R150 a_331_325.t1 a_331_325.n3 34.368
R151 a_331_325.n0 a_331_325.t4 25.312
R152 a_216_93.t1 a_216_93.n1 433.577
R153 a_216_93.n1 a_216_93.t0 230.852
R154 a_216_93.n0 a_216_93.t3 215.828
R155 a_216_93.n1 a_216_93.n0 180.432
R156 a_216_93.n0 a_216_93.t2 167.627
R157 X.n1 X.t0 170.526
R158 X X.n0 158.036
R159 X.n0 X.t1 26.595
R160 X X.n1 7.542
C0 VPB VPWR 0.16fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__xnor3_2.ext - technology: sky130A

.subckt sky130_fd_sc_hd__xnor3_2 X B C A VGND VPWR VNB VPB
X0 X.t1 a_87_21.t4 VPWR.t1 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_1198_49.t5 a_933_297.t6 VGND.t5 VNB.t11 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X2 a_87_21.t2 C.t0 a_423_325.t5 VPB.t6 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X3 a_447_49.t5 a_308_93.t2 a_87_21.t0 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X4 a_447_49.t3 B.t0 a_1198_49.t3 VNB.t7 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X5 a_87_21.t3 C.t1 a_447_49.t4 VNB.t6 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X6 a_827_297.t1 B.t1 VGND.t3 VNB.t8 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 a_933_297.t0 a_827_297.t2 a_423_325.t0 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X8 X.t3 a_87_21.t5 VGND.t1 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 a_423_325.t2 a_308_93.t3 a_87_21.t1 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X10 a_1198_49.t0 a_827_297.t3 a_423_325.t1 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11 VGND.t4 A.t0 a_933_297.t5 VNB.t10 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X12 a_308_93.t1 C.t2 VGND.t2 VNB.t5 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13 a_1198_49.t1 a_827_297.t4 a_447_49.t0 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X14 a_1198_49.t4 a_933_297.t7 VPWR.t4 VPB.t10 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 a_933_297.t1 a_827_297.t5 a_447_49.t1 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=600000u l=150000u
X16 VPWR.t0 a_87_21.t6 X.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17 VPWR.t3 A.t1 a_933_297.t2 VPB.t7 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X18 a_827_297.t0 B.t2 VPWR.t5 VPB.t11 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X19 a_423_325.t4 B.t3 a_933_297.t4 VNB.t9 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X20 VGND.t0 a_87_21.t7 X.t2 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X21 a_308_93.t0 C.t3 VPWR.t2 VPB.t5 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X22 a_447_49.t2 B.t4 a_933_297.t3 VPB.t8 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X23 a_423_325.t3 B.t5 a_1198_49.t2 VPB.t9 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
R0 a_87_21.n5 a_87_21.n4 482.376
R1 a_87_21.n4 a_87_21.n3 258.911
R2 a_87_21.n2 a_87_21.t6 212.079
R3 a_87_21.n0 a_87_21.t4 212.079
R4 a_87_21.n0 a_87_21.t5 142.7
R5 a_87_21.n1 a_87_21.t7 139.779
R6 a_87_21.n4 a_87_21.n2 89.875
R7 a_87_21.n1 a_87_21.n0 58.424
R8 a_87_21.n7 a_87_21.n6 55.16
R9 a_87_21.n5 a_87_21.t2 32.611
R10 a_87_21.n6 a_87_21.t0 30.341
R11 a_87_21.n3 a_87_21.t1 27.187
R12 a_87_21.n3 a_87_21.t3 27.187
R13 a_87_21.n6 a_87_21.n5 21.107
R14 a_87_21.n2 a_87_21.n1 2.921
R15 VPWR.n1 VPWR.t5 490.559
R16 VPWR.n14 VPWR.n13 427.426
R17 VPWR.n2 VPWR.n0 310.714
R18 VPWR.n18 VPWR.t1 160.645
R19 VPWR.n13 VPWR.t2 67.718
R20 VPWR.n13 VPWR.t0 30.376
R21 VPWR.n0 VPWR.t4 26.595
R22 VPWR.n0 VPWR.t3 26.595
R23 VPWR.n4 VPWR.n3 4.65
R24 VPWR.n6 VPWR.n5 4.65
R25 VPWR.n8 VPWR.n7 4.65
R26 VPWR.n10 VPWR.n9 4.65
R27 VPWR.n12 VPWR.n11 4.65
R28 VPWR.n15 VPWR.n14 4.65
R29 VPWR.n17 VPWR.n16 4.65
R30 VPWR.n19 VPWR.n18 4.65
R31 VPWR.n2 VPWR.n1 4.027
R32 VPWR.n4 VPWR.n2 0.137
R33 VPWR.n6 VPWR.n4 0.119
R34 VPWR.n8 VPWR.n6 0.119
R35 VPWR.n10 VPWR.n8 0.119
R36 VPWR.n12 VPWR.n10 0.119
R37 VPWR.n15 VPWR.n12 0.119
R38 VPWR.n17 VPWR.n15 0.119
R39 VPWR.n19 VPWR.n17 0.119
R40 VPWR VPWR.n19 0.022
R41 X X.n0 158.036
R42 X.n2 X.n1 145.603
R43 X.n0 X.t0 26.595
R44 X.n0 X.t1 26.595
R45 X.n1 X.t2 24.923
R46 X.n1 X.t3 24.923
R47 X X.n2 7.542
R48 VPB.t11 VPB.t8 651.09
R49 VPB.t4 VPB.t11 627.414
R50 VPB.t5 VPB.t6 621.495
R51 VPB.t3 VPB.t9 517.912
R52 VPB.t8 VPB.t3 446.884
R53 VPB.t9 VPB.t2 304.828
R54 VPB.t0 VPB.t5 304.828
R55 VPB.t2 VPB.t7 298.909
R56 VPB.t6 VPB.t4 287.071
R57 VPB.t7 VPB.t10 248.598
R58 VPB.t1 VPB.t0 248.598
R59 VPB VPB.t1 227.881
R60 a_933_297.n5 a_933_297.t3 468.615
R61 a_933_297.n9 a_933_297.n8 349.224
R62 a_933_297.n1 a_933_297.t7 241.534
R63 a_933_297.n1 a_933_297.t6 170.841
R64 a_933_297.n8 a_933_297.n1 76
R65 a_933_297.n8 a_933_297.n7 55.794
R66 a_933_297.n5 a_933_297.t4 52.25
R67 a_933_297.n0 a_933_297.t0 50.422
R68 a_933_297.n4 a_933_297.t1 42
R69 a_933_297.n10 a_933_297.n9 38.696
R70 a_933_297.n0 a_933_297.t2 28.87
R71 a_933_297.n9 a_933_297.n0 17.589
R72 a_933_297.n3 a_933_297.n2 13.805
R73 a_933_297.n6 a_933_297.n4 9.3
R74 a_933_297.n2 a_933_297.t5 9.275
R75 a_933_297.n6 a_933_297.n5 7.566
R76 a_933_297.n7 a_933_297.n6 3.71
R77 a_933_297.n4 a_933_297.n3 1
R78 VGND.n16 VGND.n15 151.577
R79 VGND.n20 VGND.t1 149.524
R80 VGND.n1 VGND.n0 122.581
R81 VGND.n2 VGND.t3 108.529
R82 VGND.n15 VGND.t2 65.714
R83 VGND.n0 VGND.t5 25.312
R84 VGND.n0 VGND.t4 25.312
R85 VGND.n15 VGND.t0 20.091
R86 VGND.n3 VGND.n2 8.282
R87 VGND.n21 VGND.n20 4.65
R88 VGND.n4 VGND.n3 4.65
R89 VGND.n6 VGND.n5 4.65
R90 VGND.n8 VGND.n7 4.65
R91 VGND.n10 VGND.n9 4.65
R92 VGND.n12 VGND.n11 4.65
R93 VGND.n14 VGND.n13 4.65
R94 VGND.n17 VGND.n16 4.65
R95 VGND.n19 VGND.n18 4.65
R96 VGND.n4 VGND.n1 0.134
R97 VGND.n6 VGND.n4 0.119
R98 VGND.n8 VGND.n6 0.119
R99 VGND.n10 VGND.n8 0.119
R100 VGND.n12 VGND.n10 0.119
R101 VGND.n14 VGND.n12 0.119
R102 VGND.n17 VGND.n14 0.119
R103 VGND.n19 VGND.n17 0.119
R104 VGND.n21 VGND.n19 0.119
R105 VGND VGND.n21 0.02
R106 a_1198_49.n2 a_1198_49.n0 297.655
R107 a_1198_49.n3 a_1198_49.t5 226.304
R108 a_1198_49.n0 a_1198_49.t1 209.825
R109 a_1198_49.n2 a_1198_49.n1 192.264
R110 a_1198_49.t4 a_1198_49.n3 176.793
R111 a_1198_49.n3 a_1198_49.n2 130.955
R112 a_1198_49.n1 a_1198_49.t0 94.776
R113 a_1198_49.n0 a_1198_49.t2 41.555
R114 a_1198_49.n1 a_1198_49.t3 38.437
R115 VNB VNB.t1 6247.32
R116 VNB.t4 VNB.t8 5888.96
R117 VNB.t5 VNB.t6 5451.11
R118 VNB.t8 VNB.t9 4522.22
R119 VNB.t2 VNB.t7 3886.67
R120 VNB.t9 VNB.t2 3691.11
R121 VNB.t7 VNB.t3 2836.76
R122 VNB.t0 VNB.t5 2538.73
R123 VNB.t3 VNB.t10 2444.44
R124 VNB.t6 VNB.t4 2151.11
R125 VNB.t10 VNB.t11 2053.33
R126 VNB.t1 VNB.t0 2030.77
R127 C.n0 C.t0 269.92
R128 C.n1 C.t3 154.239
R129 C.n0 C.t1 143.284
R130 C.n2 C.n1 132.915
R131 C.n1 C.t2 102.826
R132 C C.n2 79.584
R133 C.n2 C.n0 24.83
R134 a_423_325.n3 a_423_325.n2 490.648
R135 a_423_325.n1 a_423_325.t5 435.971
R136 a_423_325.n1 a_423_325.t2 262.941
R137 a_423_325.n2 a_423_325.n0 221.036
R138 a_423_325.n2 a_423_325.n1 116.704
R139 a_423_325.n0 a_423_325.t1 98.437
R140 a_423_325.n3 a_423_325.t3 67.718
R141 a_423_325.t0 a_423_325.n3 34.368
R142 a_423_325.n0 a_423_325.t4 25.312
R143 a_308_93.t0 a_308_93.n1 433.577
R144 a_308_93.n1 a_308_93.t1 230.852
R145 a_308_93.n0 a_308_93.t2 215.828
R146 a_308_93.n1 a_308_93.n0 180.432
R147 a_308_93.n0 a_308_93.t3 167.627
R148 a_447_49.n1 a_447_49.t4 287.572
R149 a_447_49.n2 a_447_49.n0 250.115
R150 a_447_49.n1 a_447_49.t5 176.167
R151 a_447_49.n3 a_447_49.n2 151.6
R152 a_447_49.n3 a_447_49.t0 83.109
R153 a_447_49.n0 a_447_49.t1 51.386
R154 a_447_49.n4 a_447_49.t2 40.516
R155 a_447_49.n5 a_447_49.n4 39.797
R156 a_447_49.n4 a_447_49.n3 27.703
R157 a_447_49.n0 a_447_49.t3 25.321
R158 a_447_49.n2 a_447_49.n1 8.28
R159 B.t5 B.t4 864.385
R160 B.n1 B.n0 298.84
R161 B.n0 B.t2 295.625
R162 B.n2 B.t5 235.107
R163 B.t4 B.n1 215.293
R164 B.n0 B.t1 168.699
R165 B.n2 B.t0 167.627
R166 B.n1 B.t3 167.092
R167 B B.n2 118.163
R168 a_827_297.t0 a_827_297.n3 599.237
R169 a_827_297.n0 a_827_297.t2 283.255
R170 a_827_297.n1 a_827_297.t3 173.52
R171 a_827_297.n0 a_827_297.t5 161.201
R172 a_827_297.n1 a_827_297.t4 154.239
R173 a_827_297.n2 a_827_297.n1 143.387
R174 a_827_297.n2 a_827_297.n0 94.522
R175 a_827_297.n3 a_827_297.t1 94.135
R176 a_827_297.n3 a_827_297.n2 2.703
R177 A.n0 A.t1 239.503
R178 A.n0 A.t0 168.81
R179 A A.n0 87.52
C0 VPWR VGND 0.12fF
C1 VPB VPWR 0.17fF
C2 X VGND 0.12fF
C3 VPWR X 0.20fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__xnor3_4.ext - technology: sky130A

.subckt sky130_fd_sc_hd__xnor3_4 X B C A VGND VPWR VNB VPB
X0 a_1382_49.t1 a_1011_297.t2 a_631_49.t2 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1 a_1382_49.t2 a_1117_297.t6 VGND.t0 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X2 a_1117_297.t3 a_1011_297.t3 a_631_49.t1 VNB.t5 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=600000u l=150000u
X3 a_1011_297.t0 B.t0 VGND.t7 VNB.t11 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 a_1382_49.t3 a_1117_297.t7 VPWR.t0 VPB.t10 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 a_101_21.t3 C.t0 a_631_49.t0 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X6 VPWR.t1 A.t0 a_1117_297.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 VPWR.t3 a_101_21.t4 X.t3 VPB.t5 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 a_1011_297.t1 B.t1 VPWR.t7 VPB.t11 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 a_607_325.t3 B.t2 a_1117_297.t4 VNB.t13 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X10 X.t2 a_101_21.t5 VPWR.t4 VPB.t6 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 VPWR.t5 a_101_21.t6 X.t1 VPB.t7 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 a_492_93.t0 C.t1 VPWR.t2 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X13 a_631_49.t5 B.t3 a_1117_297.t5 VPB.t12 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X14 X.t7 a_101_21.t7 VGND.t3 VNB.t6 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X15 X.t6 a_101_21.t8 VGND.t4 VNB.t7 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X16 a_607_325.t4 B.t4 a_1382_49.t5 VPB.t13 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X17 X.t0 a_101_21.t9 VPWR.t6 VPB.t8 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X18 a_631_49.t4 B.t5 a_1382_49.t4 VNB.t12 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X19 a_101_21.t2 C.t2 a_607_325.t5 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X20 VGND.t5 a_101_21.t10 X.t5 VNB.t8 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X21 a_631_49.t3 a_492_93.t2 a_101_21.t0 VPB.t9 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X22 VGND.t6 a_101_21.t11 X.t4 VNB.t9 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X23 a_607_325.t2 a_492_93.t3 a_101_21.t1 VNB.t10 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X24 VGND.t2 A.t1 a_1117_297.t1 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X25 a_1117_297.t2 a_1011_297.t4 a_607_325.t0 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X26 a_1382_49.t0 a_1011_297.t5 a_607_325.t1 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X27 a_492_93.t1 C.t3 VGND.t1 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
R0 a_1011_297.t1 a_1011_297.n3 599.237
R1 a_1011_297.n0 a_1011_297.t4 283.255
R2 a_1011_297.n1 a_1011_297.t5 173.52
R3 a_1011_297.n0 a_1011_297.t3 161.201
R4 a_1011_297.n1 a_1011_297.t2 154.239
R5 a_1011_297.n2 a_1011_297.n1 143.387
R6 a_1011_297.n2 a_1011_297.n0 94.522
R7 a_1011_297.n3 a_1011_297.t0 94.135
R8 a_1011_297.n3 a_1011_297.n2 2.703
R9 a_631_49.n3 a_631_49.t0 287.572
R10 a_631_49.n2 a_631_49.n0 250.115
R11 a_631_49.t3 a_631_49.n3 176.167
R12 a_631_49.n2 a_631_49.n1 151.601
R13 a_631_49.n4 a_631_49.t3 108.512
R14 a_631_49.n1 a_631_49.t5 85.161
R15 a_631_49.n1 a_631_49.t2 83.109
R16 a_631_49.n0 a_631_49.t1 51.386
R17 a_631_49.n0 a_631_49.t4 25.321
R18 a_631_49.n3 a_631_49.n2 8.28
R19 a_1382_49.n2 a_1382_49.n0 297.655
R20 a_1382_49.n3 a_1382_49.t2 226.304
R21 a_1382_49.n0 a_1382_49.t1 209.825
R22 a_1382_49.n2 a_1382_49.n1 192.264
R23 a_1382_49.t3 a_1382_49.n3 176.793
R24 a_1382_49.n3 a_1382_49.n2 130.955
R25 a_1382_49.n1 a_1382_49.t0 94.776
R26 a_1382_49.n0 a_1382_49.t5 41.555
R27 a_1382_49.n1 a_1382_49.t4 38.437
R28 VPB.t11 VPB.t12 651.09
R29 VPB.t9 VPB.t11 627.414
R30 VPB.t1 VPB.t2 621.495
R31 VPB.t4 VPB.t13 517.912
R32 VPB.t12 VPB.t4 446.884
R33 VPB.t13 VPB.t3 304.828
R34 VPB.t5 VPB.t1 304.828
R35 VPB.t3 VPB.t0 298.909
R36 VPB.t2 VPB.t9 287.071
R37 VPB.t7 VPB.t6 266.355
R38 VPB VPB.t8 257.476
R39 VPB.t0 VPB.t10 248.598
R40 VPB.t6 VPB.t5 248.598
R41 VPB.t8 VPB.t7 248.598
R42 a_1117_297.n5 a_1117_297.t5 468.615
R43 a_1117_297.n9 a_1117_297.n8 349.224
R44 a_1117_297.n1 a_1117_297.t7 241.534
R45 a_1117_297.n1 a_1117_297.t6 170.841
R46 a_1117_297.n8 a_1117_297.n1 76
R47 a_1117_297.n8 a_1117_297.n7 55.794
R48 a_1117_297.n5 a_1117_297.t4 52.25
R49 a_1117_297.n0 a_1117_297.t2 50.422
R50 a_1117_297.n4 a_1117_297.t3 42
R51 a_1117_297.n10 a_1117_297.n9 38.696
R52 a_1117_297.n0 a_1117_297.t0 28.87
R53 a_1117_297.n9 a_1117_297.n0 17.589
R54 a_1117_297.n3 a_1117_297.n2 13.805
R55 a_1117_297.n6 a_1117_297.n4 9.3
R56 a_1117_297.n2 a_1117_297.t1 9.275
R57 a_1117_297.n6 a_1117_297.n5 7.566
R58 a_1117_297.n7 a_1117_297.n6 3.71
R59 a_1117_297.n4 a_1117_297.n3 1
R60 VGND.n26 VGND.t4 153.187
R61 VGND.n16 VGND.n15 151.577
R62 VGND.n21 VGND.n20 128.264
R63 VGND.n1 VGND.n0 122.581
R64 VGND.n2 VGND.t7 108.529
R65 VGND.n15 VGND.t1 65.714
R66 VGND.n20 VGND.t3 26.769
R67 VGND.n0 VGND.t0 25.312
R68 VGND.n0 VGND.t2 25.312
R69 VGND.n20 VGND.t6 24.923
R70 VGND.n15 VGND.t5 20.091
R71 VGND.n27 VGND.n26 15.191
R72 VGND.n3 VGND.n2 8.282
R73 VGND.n4 VGND.n3 4.65
R74 VGND.n6 VGND.n5 4.65
R75 VGND.n8 VGND.n7 4.65
R76 VGND.n10 VGND.n9 4.65
R77 VGND.n12 VGND.n11 4.65
R78 VGND.n14 VGND.n13 4.65
R79 VGND.n17 VGND.n16 4.65
R80 VGND.n19 VGND.n18 4.65
R81 VGND.n23 VGND.n22 4.65
R82 VGND.n25 VGND.n24 4.65
R83 VGND.n22 VGND.n21 4.517
R84 VGND.n4 VGND.n1 0.134
R85 VGND.n6 VGND.n4 0.119
R86 VGND.n8 VGND.n6 0.119
R87 VGND.n10 VGND.n8 0.119
R88 VGND.n12 VGND.n10 0.119
R89 VGND.n14 VGND.n12 0.119
R90 VGND.n17 VGND.n14 0.119
R91 VGND.n19 VGND.n17 0.119
R92 VGND.n23 VGND.n19 0.119
R93 VGND.n25 VGND.n23 0.119
R94 VGND.n27 VGND.n25 0.119
R95 VGND VGND.n27 0.022
R96 VNB VNB.t7 6609.95
R97 VNB.t10 VNB.t11 5888.96
R98 VNB.t2 VNB.t1 5451.11
R99 VNB.t11 VNB.t13 4522.22
R100 VNB.t4 VNB.t12 3886.67
R101 VNB.t13 VNB.t4 3691.11
R102 VNB.t12 VNB.t5 2836.76
R103 VNB.t8 VNB.t2 2538.73
R104 VNB.t5 VNB.t3 2444.44
R105 VNB.t1 VNB.t10 2151.11
R106 VNB.t9 VNB.t6 2079.12
R107 VNB.t3 VNB.t0 2053.33
R108 VNB.t6 VNB.t8 2030.77
R109 VNB.t7 VNB.t9 2030.77
R110 B.t4 B.t3 864.385
R111 B.n1 B.n0 298.84
R112 B.n0 B.t1 295.625
R113 B.n2 B.t4 235.107
R114 B.t3 B.n1 215.293
R115 B.n0 B.t0 168.699
R116 B.n2 B.t5 167.627
R117 B.n1 B.t2 167.092
R118 B B.n2 118.163
R119 VPWR.n1 VPWR.t7 490.559
R120 VPWR.n14 VPWR.n13 427.426
R121 VPWR.n2 VPWR.n0 310.714
R122 VPWR.n24 VPWR.t6 159.459
R123 VPWR.n19 VPWR.n18 132.865
R124 VPWR.n13 VPWR.t2 67.718
R125 VPWR.n18 VPWR.t4 32.505
R126 VPWR.n13 VPWR.t3 30.376
R127 VPWR.n18 VPWR.t5 26.595
R128 VPWR.n0 VPWR.t0 26.595
R129 VPWR.n0 VPWR.t1 26.595
R130 VPWR.n25 VPWR.n24 15.191
R131 VPWR.n4 VPWR.n3 4.65
R132 VPWR.n6 VPWR.n5 4.65
R133 VPWR.n8 VPWR.n7 4.65
R134 VPWR.n10 VPWR.n9 4.65
R135 VPWR.n12 VPWR.n11 4.65
R136 VPWR.n15 VPWR.n14 4.65
R137 VPWR.n17 VPWR.n16 4.65
R138 VPWR.n21 VPWR.n20 4.65
R139 VPWR.n23 VPWR.n22 4.65
R140 VPWR.n20 VPWR.n19 4.517
R141 VPWR.n2 VPWR.n1 4.027
R142 VPWR.n4 VPWR.n2 0.137
R143 VPWR.n6 VPWR.n4 0.119
R144 VPWR.n8 VPWR.n6 0.119
R145 VPWR.n10 VPWR.n8 0.119
R146 VPWR.n12 VPWR.n10 0.119
R147 VPWR.n15 VPWR.n12 0.119
R148 VPWR.n17 VPWR.n15 0.119
R149 VPWR.n21 VPWR.n17 0.119
R150 VPWR.n23 VPWR.n21 0.119
R151 VPWR.n25 VPWR.n23 0.119
R152 VPWR VPWR.n25 0.022
R153 C.n0 C.t2 269.92
R154 C.n1 C.t1 154.239
R155 C.n0 C.t0 143.284
R156 C.n2 C.n1 132.915
R157 C.n1 C.t3 102.826
R158 C C.n2 79.584
R159 C.n2 C.n0 24.83
R160 a_101_21.n8 a_101_21.n7 482.376
R161 a_101_21.n7 a_101_21.n6 258.911
R162 a_101_21.n5 a_101_21.t4 212.079
R163 a_101_21.n3 a_101_21.t5 212.079
R164 a_101_21.n1 a_101_21.t6 212.079
R165 a_101_21.n0 a_101_21.t9 212.079
R166 a_101_21.n1 a_101_21.t11 139.779
R167 a_101_21.n0 a_101_21.t8 139.779
R168 a_101_21.n2 a_101_21.t7 139.779
R169 a_101_21.n4 a_101_21.t10 139.779
R170 a_101_21.n7 a_101_21.n5 89.875
R171 a_101_21.n2 a_101_21.n1 62.806
R172 a_101_21.n1 a_101_21.n0 61.345
R173 a_101_21.n4 a_101_21.n3 58.424
R174 a_101_21.n10 a_101_21.n9 55.16
R175 a_101_21.n8 a_101_21.t2 32.611
R176 a_101_21.n9 a_101_21.t0 30.341
R177 a_101_21.n6 a_101_21.t1 27.187
R178 a_101_21.n6 a_101_21.t3 27.187
R179 a_101_21.n9 a_101_21.n8 21.107
R180 a_101_21.n5 a_101_21.n4 2.921
R181 a_101_21.n3 a_101_21.n2 2.921
R182 A.n0 A.t0 239.503
R183 A.n0 A.t1 168.81
R184 A A.n0 87.52
R185 X X.n0 158.036
R186 X.n4 X.n2 117.525
R187 X.n4 X.n3 116.323
R188 X.n5 X.n1 114.126
R189 X.n5 X.n4 30.836
R190 X.n0 X.t3 26.595
R191 X.n0 X.t2 26.595
R192 X.n2 X.t1 26.595
R193 X.n2 X.t0 26.595
R194 X.n1 X.t5 24.923
R195 X.n1 X.t7 24.923
R196 X.n3 X.t4 24.923
R197 X.n3 X.t6 24.923
R198 X.n6 X.n5 14.236
R199 X X.n6 7.542
R200 a_607_325.n3 a_607_325.n2 490.648
R201 a_607_325.n1 a_607_325.t5 435.971
R202 a_607_325.n1 a_607_325.t2 262.941
R203 a_607_325.n2 a_607_325.n0 221.036
R204 a_607_325.n2 a_607_325.n1 116.704
R205 a_607_325.n0 a_607_325.t1 98.437
R206 a_607_325.n3 a_607_325.t4 67.718
R207 a_607_325.t0 a_607_325.n3 34.368
R208 a_607_325.n0 a_607_325.t3 25.312
R209 a_492_93.t0 a_492_93.n1 433.577
R210 a_492_93.n1 a_492_93.t1 230.852
R211 a_492_93.n0 a_492_93.t2 215.828
R212 a_492_93.n1 a_492_93.n0 180.432
R213 a_492_93.n0 a_492_93.t3 167.627
C0 VPWR X 0.61fF
C1 VPWR VGND 0.14fF
C2 VPB VPWR 0.19fF
C3 X VGND 0.29fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__xor2_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__xor2_1 B X A VPWR VGND VNB VPB
X0 X.t1 a_35_297.t3 a_285_297.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 X.t2 B.t0 a_285_47.t0 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 a_35_297.t1 B.t1 VGND.t1 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 a_117_297.t1 B.t2 a_35_297.t2 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 VPWR.t1 B.t3 a_285_297.t1 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 VGND.t2 A.t0 a_35_297.t0 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 VGND.t0 a_35_297.t4 X.t0 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 a_285_297.t2 A.t1 VPWR.t2 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 VPWR.t0 A.t2 a_117_297.t0 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 a_285_47.t1 A.t3 VGND.t3 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
R0 a_35_297.t2 a_35_297.n2 296.59
R1 a_35_297.n2 a_35_297.n1 267.921
R2 a_35_297.n1 a_35_297.t3 215.48
R3 a_35_297.n1 a_35_297.t4 139.779
R4 a_35_297.n2 a_35_297.n0 104.17
R5 a_35_297.n0 a_35_297.t0 24.923
R6 a_35_297.n0 a_35_297.t1 24.923
R7 a_285_297.t0 a_285_297.n0 369.053
R8 a_285_297.n0 a_285_297.t1 26.595
R9 a_285_297.n0 a_285_297.t2 26.595
R10 X.n1 X.t1 138.138
R11 X.n1 X.n0 129.705
R12 X.n0 X.t2 63.067
R13 X.n0 X.t0 52.034
R14 X X.n1 0.2
R15 VPB.t1 VPB.t0 556.386
R16 VPB.t4 VPB.t1 248.598
R17 VPB.t2 VPB.t4 248.598
R18 VPB.t3 VPB.t2 248.598
R19 VPB VPB.t3 216.043
R20 B.n1 B.t2 241.534
R21 B.n0 B.t3 241.534
R22 B.n2 B.n0 173.88
R23 B.n1 B.t1 169.234
R24 B.n0 B.t0 169.234
R25 B B.n1 90.889
R26 B B.n2 4.894
R27 B.n2 B 4.44
R28 a_285_47.t0 a_285_47.t1 49.846
R29 VNB VNB.t1 6271.49
R30 VNB.t2 VNB.t0 4448.35
R31 VNB.t4 VNB.t2 2030.77
R32 VNB.t3 VNB.t4 2030.77
R33 VNB.t1 VNB.t3 2030.77
R34 VGND.n5 VGND.t1 186.088
R35 VGND.n1 VGND.n0 107.627
R36 VGND.n2 VGND.t0 102.907
R37 VGND.n0 VGND.t3 24.923
R38 VGND.n0 VGND.t2 24.923
R39 VGND.n6 VGND.n5 4.65
R40 VGND.n4 VGND.n3 4.65
R41 VGND.n2 VGND.n1 3.952
R42 VGND.n4 VGND.n2 0.14
R43 VGND.n6 VGND.n4 0.119
R44 VGND VGND.n6 0.022
R45 a_117_297.t0 a_117_297.t1 53.19
R46 VPWR.n1 VPWR.t1 557.792
R47 VPWR.n1 VPWR.n0 182.569
R48 VPWR.n0 VPWR.t2 26.595
R49 VPWR.n0 VPWR.t0 26.595
R50 VPWR VPWR.n1 0.369
R51 A.n0 A.t1 212.079
R52 A.n1 A.t2 212.079
R53 A.n0 A.t3 139.779
R54 A.n1 A.t0 139.779
R55 A A.n2 77.28
R56 A.n2 A.n0 37.245
R57 A.n2 A.n1 24.1
C0 X VGND 0.26fF
C1 B A 0.33fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__xor2_2.ext - technology: sky130A

.subckt sky130_fd_sc_hd__xor2_2 VPWR VGND X B A VNB VPB
X0 a_27_297.t1 A.t0 VPWR.t3 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_470_47.t1 A.t1 VGND.t3 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 a_470_297.t1 A.t2 VPWR.t1 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 VPWR.t0 A.t3 a_470_297.t0 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 a_112_47.t1 B.t0 VGND.t6 VNB.t7 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 a_470_47.t3 B.t1 X.t1 VNB.t8 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 VGND.t1 A.t4 a_112_47.t5 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 a_112_47.t4 A.t5 VGND.t0 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 VGND.t7 B.t2 a_112_47.t0 VNB.t9 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 VPWR.t2 A.t6 a_27_297.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 a_470_297.t4 B.t3 VPWR.t4 VPB.t8 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 X.t3 a_112_47.t6 VGND.t4 VNB.t5 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 VPWR.t5 B.t4 a_470_297.t5 VPB.t9 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13 VGND.t5 a_112_47.t7 X.t2 VNB.t6 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14 VGND.t2 A.t7 a_470_47.t0 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X15 a_27_297.t2 B.t5 a_112_47.t3 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16 X.t5 a_112_47.t8 a_470_297.t3 VPB.t7 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17 a_470_297.t2 a_112_47.t9 X.t4 VPB.t6 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X18 X.t0 B.t6 a_470_47.t2 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X19 a_112_47.t2 B.t7 a_27_297.t3 VPB.t5 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
R0 A.n3 A.t0 212.079
R1 A.n4 A.t6 212.079
R2 A.n0 A.t2 212.079
R3 A.n1 A.t3 212.079
R4 A A.n2 160.539
R5 A.n3 A.t4 139.779
R6 A.n4 A.t5 139.779
R7 A.n0 A.t1 139.779
R8 A.n1 A.t7 139.779
R9 A A.n5 113.965
R10 A.n5 A.n4 32.863
R11 A.n5 A.n3 28.481
R12 A.n2 A.n0 27.572
R13 A.n2 A.n1 22.735
R14 VPWR.n1 VPWR.n0 314.004
R15 VPWR.n13 VPWR.n12 314.004
R16 VPWR.n3 VPWR.n2 313.497
R17 VPWR.n2 VPWR.t5 37.43
R18 VPWR.n2 VPWR.t4 26.595
R19 VPWR.n0 VPWR.t1 26.595
R20 VPWR.n0 VPWR.t0 26.595
R21 VPWR.n12 VPWR.t3 26.595
R22 VPWR.n12 VPWR.t2 26.595
R23 VPWR.n5 VPWR.n4 4.65
R24 VPWR.n7 VPWR.n6 4.65
R25 VPWR.n9 VPWR.n8 4.65
R26 VPWR.n11 VPWR.n10 4.65
R27 VPWR.n14 VPWR.n13 4.017
R28 VPWR.n3 VPWR.n1 3.998
R29 VPWR.n5 VPWR.n3 0.241
R30 VPWR.n14 VPWR.n11 0.135
R31 VPWR VPWR.n14 0.125
R32 VPWR.n7 VPWR.n5 0.119
R33 VPWR.n9 VPWR.n7 0.119
R34 VPWR.n11 VPWR.n9 0.119
R35 a_27_297.n0 a_27_297.t2 583.515
R36 a_27_297.n1 a_27_297.t0 208.715
R37 a_27_297.n2 a_27_297.t3 23.64
R38 a_27_297.n4 a_27_297.n3 13.79
R39 a_27_297.t1 a_27_297.n4 12.805
R40 a_27_297.n2 a_27_297.n1 9.3
R41 a_27_297.n1 a_27_297.n0 3.327
R42 a_27_297.n3 a_27_297.n2 2.955
R43 VPB.t8 VPB.t7 556.386
R44 VPB.t4 VPB.t1 556.386
R45 VPB.t9 VPB.t8 281.152
R46 VPB.t7 VPB.t6 248.598
R47 VPB.t2 VPB.t9 248.598
R48 VPB.t1 VPB.t2 248.598
R49 VPB.t5 VPB.t4 248.598
R50 VPB.t3 VPB.t5 248.598
R51 VPB.t0 VPB.t3 248.598
R52 VPB VPB.t0 201.246
R53 VGND.n1 VGND.t5 204.432
R54 VGND.n0 VGND.t4 193.925
R55 VGND.n14 VGND.t7 193.925
R56 VGND.n25 VGND.t0 189.645
R57 VGND.n9 VGND.n8 115.464
R58 VGND.n20 VGND.n19 115.464
R59 VGND.n8 VGND.t3 24.923
R60 VGND.n8 VGND.t2 24.923
R61 VGND.n19 VGND.t6 24.923
R62 VGND.n19 VGND.t1 24.923
R63 VGND.n1 VGND.n0 11.464
R64 VGND.n15 VGND.n14 8.658
R65 VGND.n26 VGND.n25 8.038
R66 VGND.n10 VGND.n9 7.152
R67 VGND.n3 VGND.n2 4.65
R68 VGND.n5 VGND.n4 4.65
R69 VGND.n7 VGND.n6 4.65
R70 VGND.n11 VGND.n10 4.65
R71 VGND.n13 VGND.n12 4.65
R72 VGND.n16 VGND.n15 4.65
R73 VGND.n18 VGND.n17 4.65
R74 VGND.n22 VGND.n21 4.65
R75 VGND.n24 VGND.n23 4.65
R76 VGND.n21 VGND.n20 2.635
R77 VGND.n3 VGND.n1 0.339
R78 VGND.n5 VGND.n3 0.119
R79 VGND.n7 VGND.n5 0.119
R80 VGND.n11 VGND.n7 0.119
R81 VGND.n13 VGND.n11 0.119
R82 VGND.n16 VGND.n13 0.119
R83 VGND.n18 VGND.n16 0.119
R84 VGND.n22 VGND.n18 0.119
R85 VGND.n24 VGND.n22 0.119
R86 VGND.n26 VGND.n24 0.119
R87 VGND VGND.n26 0.022
R88 a_470_47.n0 a_470_47.t3 227.048
R89 a_470_47.n0 a_470_47.t0 142.298
R90 a_470_47.n1 a_470_47.n0 92.5
R91 a_470_47.n1 a_470_47.t2 24.923
R92 a_470_47.t1 a_470_47.n1 24.923
R93 VNB VNB.t1 6150.61
R94 VNB.t8 VNB.t5 4545.05
R95 VNB.t9 VNB.t0 4545.05
R96 VNB.t4 VNB.t8 2296.7
R97 VNB.t5 VNB.t6 2030.77
R98 VNB.t3 VNB.t4 2030.77
R99 VNB.t0 VNB.t3 2030.77
R100 VNB.t7 VNB.t9 2030.77
R101 VNB.t2 VNB.t7 2030.77
R102 VNB.t1 VNB.t2 2030.77
R103 a_470_297.n0 a_470_297.t2 227.943
R104 a_470_297.n2 a_470_297.t0 226.924
R105 a_470_297.n1 a_470_297.t4 172.845
R106 a_470_297.n0 a_470_297.t3 172.845
R107 a_470_297.n3 a_470_297.n2 155.084
R108 a_470_297.n2 a_470_297.n1 50.916
R109 a_470_297.n3 a_470_297.t5 26.595
R110 a_470_297.t1 a_470_297.n3 26.595
R111 a_470_297.n1 a_470_297.n0 9.788
R112 B.n5 B.t3 212.079
R113 B.n3 B.t4 212.079
R114 B.n0 B.t5 212.079
R115 B.n1 B.t7 212.079
R116 B.n5 B.t1 139.779
R117 B.n3 B.t6 139.779
R118 B.n0 B.t2 139.779
R119 B.n1 B.t0 139.779
R120 B.n7 B.n2 98.993
R121 B.n2 B.n0 54.042
R122 B.n6 B.n4 48.912
R123 B.n6 B.n5 10.838
R124 B.n4 B.n3 8.763
R125 B.n7 B.n6 8.353
R126 B.n2 B.n1 7.303
R127 B B.n7 3.081
R128 a_112_47.n6 a_112_47.n2 368.326
R129 a_112_47.n7 a_112_47.n6 292.5
R130 a_112_47.n0 a_112_47.t9 212.079
R131 a_112_47.n1 a_112_47.t8 212.079
R132 a_112_47.n6 a_112_47.n5 184.803
R133 a_112_47.n0 a_112_47.t7 139.779
R134 a_112_47.n1 a_112_47.t6 139.779
R135 a_112_47.n5 a_112_47.n3 88.89
R136 a_112_47.n5 a_112_47.n4 52.624
R137 a_112_47.n2 a_112_47.n0 36.515
R138 a_112_47.t3 a_112_47.n7 26.595
R139 a_112_47.n7 a_112_47.t2 26.595
R140 a_112_47.n3 a_112_47.t0 24.923
R141 a_112_47.n3 a_112_47.t1 24.923
R142 a_112_47.n4 a_112_47.t5 24.923
R143 a_112_47.n4 a_112_47.t4 24.923
R144 a_112_47.n2 a_112_47.n1 24.83
R145 X.n3 X.n2 181.99
R146 X X.n0 170.738
R147 X.n3 X.n1 92.5
R148 X X.n3 39.879
R149 X.n2 X.t0 35.076
R150 X.n0 X.t4 26.595
R151 X.n0 X.t5 26.595
R152 X.n1 X.t2 24.923
R153 X.n1 X.t3 24.923
R154 X.n2 X.t1 24.923
C0 VPB VPWR 0.12fF
C1 A B 0.35fF
C2 B VGND 0.16fF
C3 B VPWR 0.11fF
C4 X VGND 0.15fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__xor2_4.ext - technology: sky130A

.subckt sky130_fd_sc_hd__xor2_4 X B A VGND VPWR VNB VPB
X0 a_27_297.t3 A.t0 VPWR.t7 VPB.t7 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_806_47.t7 B.t0 X.t11 VNB.t19 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 a_806_47.t6 B.t1 X.t10 VNB.t18 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 a_112_47.t3 A.t1 VGND.t7 VNB.t7 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 a_27_297.t4 B.t2 a_112_47.t7 VPB.t12 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 a_806_297.t7 a_112_47.t12 X.t0 VPB.t8 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 VGND.t8 a_112_47.t13 X.t1 VNB.t8 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 X.t9 B.t3 a_806_47.t5 VNB.t17 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 X.t2 a_112_47.t14 a_806_297.t6 VPB.t9 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 a_112_47.t6 B.t4 a_27_297.t5 VPB.t13 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 a_806_297.t11 B.t5 VPWR.t8 VPB.t14 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 VGND.t3 A.t2 a_806_47.t3 VNB.t6 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 X.t8 B.t6 a_806_47.t4 VNB.t16 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 VGND.t2 A.t3 a_806_47.t2 VNB.t5 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14 a_806_297.t5 a_112_47.t15 X.t3 VPB.t10 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 VGND.t6 A.t4 a_112_47.t2 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X16 a_112_47.t1 A.t5 VGND.t5 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X17 VGND.t4 A.t6 a_112_47.t0 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X18 VPWR.t6 A.t7 a_27_297.t2 VPB.t6 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X19 a_806_297.t10 B.t7 VPWR.t9 VPB.t15 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X20 VPWR.t10 B.t8 a_806_297.t9 VPB.t16 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X21 VGND.t15 B.t9 a_112_47.t11 VNB.t15 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X22 VGND.t14 B.t10 a_112_47.t10 VNB.t14 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X23 VPWR.t11 B.t11 a_806_297.t8 VPB.t17 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X24 a_806_47.t1 A.t8 VGND.t1 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X25 a_806_47.t0 A.t9 VGND.t0 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X26 a_27_297.t6 B.t12 a_112_47.t5 VPB.t18 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X27 a_112_47.t9 B.t13 VGND.t13 VNB.t13 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X28 VGND.t9 a_112_47.t16 X.t4 VNB.t9 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X29 a_806_297.t3 A.t10 VPWR.t3 VPB.t5 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X30 a_112_47.t8 B.t14 VGND.t12 VNB.t12 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X31 a_112_47.t4 B.t15 a_27_297.t7 VPB.t19 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X32 VPWR.t2 A.t11 a_806_297.t2 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X33 a_27_297.t1 A.t12 VPWR.t5 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X34 X.t5 a_112_47.t17 a_806_297.t4 VPB.t11 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X35 VPWR.t4 A.t13 a_27_297.t0 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X36 a_806_297.t1 A.t14 VPWR.t1 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X37 X.t6 a_112_47.t18 VGND.t10 VNB.t10 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X38 X.t7 a_112_47.t19 VGND.t11 VNB.t11 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X39 VPWR.t0 A.t15 a_806_297.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
R0 A.n13 A.n10 355.124
R1 A.n11 A.t12 212.079
R2 A.n14 A.t13 212.079
R3 A.n19 A.t0 212.079
R4 A.n17 A.t7 212.079
R5 A.n0 A.t10 212.079
R6 A.n2 A.t11 212.079
R7 A.n5 A.t14 212.079
R8 A.n8 A.t15 212.079
R9 A.n11 A.t6 139.779
R10 A.n14 A.t1 139.779
R11 A.n19 A.t4 139.779
R12 A.n17 A.t5 139.779
R13 A.n0 A.t9 139.779
R14 A.n2 A.t3 139.779
R15 A.n5 A.t8 139.779
R16 A.n8 A.t2 139.779
R17 A.n4 A.n1 97.76
R18 A.n21 A.n18 97.76
R19 A.n10 A.n9 76
R20 A.n4 A.n3 76
R21 A.n7 A.n6 76
R22 A.n13 A.n12 76
R23 A.n16 A.n15 76
R24 A.n21 A.n20 76
R25 A.n7 A.n4 21.76
R26 A.n10 A.n7 21.76
R27 A.n16 A.n13 21.76
R28 A.n12 A.n11 18.987
R29 A.n9 A.n8 18.257
R30 A.n1 A.n0 16.796
R31 A.n18 A.n17 16.066
R32 A A.n16 13.44
R33 A A.n21 8.32
R34 A.n15 A.n14 7.303
R35 A.n6 A.n5 6.572
R36 A.n3 A.n2 5.112
R37 A.n20 A.n19 4.381
R38 VPWR.n3 VPWR.n2 315.572
R39 VPWR.n1 VPWR.n0 311.956
R40 VPWR.n7 VPWR.n6 311.956
R41 VPWR.n12 VPWR.n11 311.956
R42 VPWR.n26 VPWR.n25 311.956
R43 VPWR.n31 VPWR.n30 311.956
R44 VPWR.n2 VPWR.t3 26.595
R45 VPWR.n2 VPWR.t2 26.595
R46 VPWR.n0 VPWR.t1 26.595
R47 VPWR.n0 VPWR.t0 26.595
R48 VPWR.n6 VPWR.t8 26.595
R49 VPWR.n6 VPWR.t10 26.595
R50 VPWR.n11 VPWR.t9 26.595
R51 VPWR.n11 VPWR.t11 26.595
R52 VPWR.n25 VPWR.t5 26.595
R53 VPWR.n25 VPWR.t4 26.595
R54 VPWR.n30 VPWR.t7 26.595
R55 VPWR.n30 VPWR.t6 26.595
R56 VPWR.n13 VPWR.n12 6.023
R57 VPWR.n5 VPWR.n4 4.65
R58 VPWR.n8 VPWR.n7 4.65
R59 VPWR.n10 VPWR.n9 4.65
R60 VPWR.n14 VPWR.n13 4.65
R61 VPWR.n16 VPWR.n15 4.65
R62 VPWR.n18 VPWR.n17 4.65
R63 VPWR.n20 VPWR.n19 4.65
R64 VPWR.n22 VPWR.n21 4.65
R65 VPWR.n24 VPWR.n23 4.65
R66 VPWR.n27 VPWR.n26 4.65
R67 VPWR.n29 VPWR.n28 4.65
R68 VPWR.n32 VPWR.n31 4.017
R69 VPWR.n3 VPWR.n1 3.831
R70 VPWR.n5 VPWR.n3 0.232
R71 VPWR.n32 VPWR.n29 0.135
R72 VPWR VPWR.n32 0.125
R73 VPWR.n8 VPWR.n5 0.119
R74 VPWR.n10 VPWR.n8 0.119
R75 VPWR.n14 VPWR.n10 0.119
R76 VPWR.n16 VPWR.n14 0.119
R77 VPWR.n18 VPWR.n16 0.119
R78 VPWR.n20 VPWR.n18 0.119
R79 VPWR.n22 VPWR.n20 0.119
R80 VPWR.n24 VPWR.n22 0.119
R81 VPWR.n27 VPWR.n24 0.119
R82 VPWR.n29 VPWR.n27 0.119
R83 a_27_297.n1 a_27_297.n0 292.5
R84 a_27_297.n1 a_27_297.t4 230.296
R85 a_27_297.n4 a_27_297.t2 213.188
R86 a_27_297.n5 a_27_297.n4 153.804
R87 a_27_297.n3 a_27_297.n2 142.024
R88 a_27_297.n3 a_27_297.n1 61.677
R89 a_27_297.n4 a_27_297.n3 46.108
R90 a_27_297.n2 a_27_297.t7 26.595
R91 a_27_297.n2 a_27_297.t1 26.595
R92 a_27_297.n0 a_27_297.t5 26.595
R93 a_27_297.n0 a_27_297.t6 26.595
R94 a_27_297.n5 a_27_297.t0 26.595
R95 a_27_297.t3 a_27_297.n5 26.595
R96 VPB.t5 VPB.t10 562.305
R97 VPB.t12 VPB.t17 556.386
R98 VPB.t8 VPB.t11 248.598
R99 VPB.t9 VPB.t8 248.598
R100 VPB.t10 VPB.t9 248.598
R101 VPB.t4 VPB.t5 248.598
R102 VPB.t1 VPB.t4 248.598
R103 VPB.t0 VPB.t1 248.598
R104 VPB.t14 VPB.t0 248.598
R105 VPB.t16 VPB.t14 248.598
R106 VPB.t15 VPB.t16 248.598
R107 VPB.t17 VPB.t15 248.598
R108 VPB.t13 VPB.t12 248.598
R109 VPB.t18 VPB.t13 248.598
R110 VPB.t19 VPB.t18 248.598
R111 VPB.t3 VPB.t19 248.598
R112 VPB.t2 VPB.t3 248.598
R113 VPB.t7 VPB.t2 248.598
R114 VPB.t6 VPB.t7 248.598
R115 VPB VPB.t6 201.246
R116 B.n0 B.t5 212.079
R117 B.n1 B.t8 212.079
R118 B.n2 B.t7 212.079
R119 B.n6 B.t11 212.079
R120 B.n13 B.t2 212.079
R121 B.n11 B.t4 212.079
R122 B.n10 B.t12 212.079
R123 B.n9 B.t15 212.079
R124 B.n0 B.t0 139.779
R125 B.n1 B.t3 139.779
R126 B.n2 B.t1 139.779
R127 B.n6 B.t6 139.779
R128 B.n13 B.t10 139.779
R129 B.n11 B.t14 139.779
R130 B.n10 B.t9 139.779
R131 B.n9 B.t13 139.779
R132 B.n15 B.n12 97.76
R133 B.n5 B.n3 97.76
R134 B.n5 B.n4 76
R135 B.n8 B.n7 76
R136 B.n17 B.n16 76
R137 B.n15 B.n14 76
R138 B.n1 B.n0 61.345
R139 B.n11 B.n10 61.345
R140 B.n10 B.n9 61.345
R141 B.n3 B.n1 54.042
R142 B.n7 B.n6 30.672
R143 B.n8 B.n5 21.76
R144 B.n17 B.n15 21.76
R145 B B.n8 21.12
R146 B.n12 B.n11 18.987
R147 B.n3 B.n2 7.303
R148 B.n14 B.n13 7.303
R149 B B.n17 0.64
R150 X.n1 X.t3 213.363
R151 X.n1 X.n0 153.805
R152 X.n5 X.n3 127.137
R153 X.n10 X.t5 126.335
R154 X.n8 X.n7 52.818
R155 X.n6 X.n2 52.624
R156 X.n9 X.n8 49.266
R157 X.n9 X.n1 42.979
R158 X.n8 X.n6 38.592
R159 X.n4 X.t11 33.431
R160 X.n0 X.t0 26.595
R161 X.n0 X.t2 26.595
R162 X.n2 X.t4 24.923
R163 X.n2 X.t6 24.923
R164 X.n3 X.t10 24.923
R165 X.n3 X.t8 24.923
R166 X.n7 X.t1 24.923
R167 X.n7 X.t7 24.923
R168 X.n6 X.n5 23.997
R169 X.n4 X.t9 14.347
R170 X.n5 X.n4 8.705
R171 X.n10 X.n9 5.649
R172 X X.n10 1.656
R173 a_806_47.n4 a_806_47.t4 219.833
R174 a_806_47.n1 a_806_47.t0 128.218
R175 a_806_47.n5 a_806_47.n4 92.5
R176 a_806_47.n4 a_806_47.n3 53.163
R177 a_806_47.n1 a_806_47.n0 52.624
R178 a_806_47.n3 a_806_47.n1 48.574
R179 a_806_47.n3 a_806_47.n2 42.273
R180 a_806_47.n2 a_806_47.t3 24.923
R181 a_806_47.n2 a_806_47.t7 24.923
R182 a_806_47.n0 a_806_47.t2 24.923
R183 a_806_47.n0 a_806_47.t1 24.923
R184 a_806_47.n5 a_806_47.t5 24.923
R185 a_806_47.t6 a_806_47.n5 24.923
R186 VNB VNB.t3 6150.61
R187 VNB.t0 VNB.t10 4593.41
R188 VNB.t14 VNB.t16 4545.05
R189 VNB.t11 VNB.t8 2030.77
R190 VNB.t9 VNB.t11 2030.77
R191 VNB.t10 VNB.t9 2030.77
R192 VNB.t5 VNB.t0 2030.77
R193 VNB.t1 VNB.t5 2030.77
R194 VNB.t6 VNB.t1 2030.77
R195 VNB.t19 VNB.t6 2030.77
R196 VNB.t17 VNB.t19 2030.77
R197 VNB.t18 VNB.t17 2030.77
R198 VNB.t16 VNB.t18 2030.77
R199 VNB.t12 VNB.t14 2030.77
R200 VNB.t15 VNB.t12 2030.77
R201 VNB.t13 VNB.t15 2030.77
R202 VNB.t2 VNB.t13 2030.77
R203 VNB.t7 VNB.t2 2030.77
R204 VNB.t4 VNB.t7 2030.77
R205 VNB.t3 VNB.t4 2030.77
R206 VGND.n2 VGND.t8 198.633
R207 VGND.n5 VGND.t10 193.925
R208 VGND.n51 VGND.t5 184.833
R209 VGND.n1 VGND.n0 115.464
R210 VGND.n11 VGND.n10 115.464
R211 VGND.n17 VGND.n16 115.464
R212 VGND.n34 VGND.n33 115.464
R213 VGND.n40 VGND.n39 115.464
R214 VGND.n46 VGND.n45 115.464
R215 VGND.n28 VGND.t14 107.818
R216 VGND.n0 VGND.t11 24.923
R217 VGND.n0 VGND.t9 24.923
R218 VGND.n10 VGND.t0 24.923
R219 VGND.n10 VGND.t2 24.923
R220 VGND.n16 VGND.t1 24.923
R221 VGND.n16 VGND.t3 24.923
R222 VGND.n33 VGND.t12 24.923
R223 VGND.n33 VGND.t15 24.923
R224 VGND.n39 VGND.t13 24.923
R225 VGND.n39 VGND.t4 24.923
R226 VGND.n45 VGND.t7 24.923
R227 VGND.n45 VGND.t6 24.923
R228 VGND.n35 VGND.n34 14.682
R229 VGND.n2 VGND.n1 10.348
R230 VGND.n41 VGND.n40 8.658
R231 VGND.n29 VGND.n28 6.776
R232 VGND.n52 VGND.n51 4.65
R233 VGND.n4 VGND.n3 4.65
R234 VGND.n7 VGND.n6 4.65
R235 VGND.n9 VGND.n8 4.65
R236 VGND.n13 VGND.n12 4.65
R237 VGND.n15 VGND.n14 4.65
R238 VGND.n19 VGND.n18 4.65
R239 VGND.n21 VGND.n20 4.65
R240 VGND.n23 VGND.n22 4.65
R241 VGND.n25 VGND.n24 4.65
R242 VGND.n27 VGND.n26 4.65
R243 VGND.n30 VGND.n29 4.65
R244 VGND.n32 VGND.n31 4.65
R245 VGND.n36 VGND.n35 4.65
R246 VGND.n38 VGND.n37 4.65
R247 VGND.n42 VGND.n41 4.65
R248 VGND.n44 VGND.n43 4.65
R249 VGND.n48 VGND.n47 4.65
R250 VGND.n50 VGND.n49 4.65
R251 VGND.n18 VGND.n17 3.388
R252 VGND.n12 VGND.n11 2.635
R253 VGND.n47 VGND.n46 2.635
R254 VGND.n6 VGND.n5 0.376
R255 VGND.n4 VGND.n2 0.326
R256 VGND.n7 VGND.n4 0.119
R257 VGND.n9 VGND.n7 0.119
R258 VGND.n13 VGND.n9 0.119
R259 VGND.n15 VGND.n13 0.119
R260 VGND.n19 VGND.n15 0.119
R261 VGND.n21 VGND.n19 0.119
R262 VGND.n23 VGND.n21 0.119
R263 VGND.n25 VGND.n23 0.119
R264 VGND.n27 VGND.n25 0.119
R265 VGND.n30 VGND.n27 0.119
R266 VGND.n32 VGND.n30 0.119
R267 VGND.n36 VGND.n32 0.119
R268 VGND.n38 VGND.n36 0.119
R269 VGND.n42 VGND.n38 0.119
R270 VGND.n44 VGND.n42 0.119
R271 VGND.n48 VGND.n44 0.119
R272 VGND.n50 VGND.n48 0.119
R273 VGND.n52 VGND.n50 0.119
R274 VGND VGND.n52 0.022
R275 a_112_47.n19 a_112_47.n18 341.628
R276 a_112_47.n18 a_112_47.n0 297.108
R277 a_112_47.n1 a_112_47.t17 212.079
R278 a_112_47.n3 a_112_47.t12 212.079
R279 a_112_47.n7 a_112_47.t14 212.079
R280 a_112_47.n6 a_112_47.t15 212.079
R281 a_112_47.n17 a_112_47.n16 211.014
R282 a_112_47.n1 a_112_47.t13 139.779
R283 a_112_47.n3 a_112_47.t19 139.779
R284 a_112_47.n7 a_112_47.t16 139.779
R285 a_112_47.n6 a_112_47.t18 139.779
R286 a_112_47.n17 a_112_47.n9 108.796
R287 a_112_47.n5 a_112_47.n2 97.76
R288 a_112_47.n12 a_112_47.n10 88.89
R289 a_112_47.n9 a_112_47.n8 76
R290 a_112_47.n5 a_112_47.n4 76
R291 a_112_47.n7 a_112_47.n6 61.345
R292 a_112_47.n12 a_112_47.n11 52.624
R293 a_112_47.n14 a_112_47.n13 52.624
R294 a_112_47.n16 a_112_47.n15 52.624
R295 a_112_47.n18 a_112_47.n17 37.104
R296 a_112_47.n14 a_112_47.n12 36.266
R297 a_112_47.n16 a_112_47.n14 36.266
R298 a_112_47.n0 a_112_47.t5 26.595
R299 a_112_47.n0 a_112_47.t4 26.595
R300 a_112_47.t7 a_112_47.n19 26.595
R301 a_112_47.n19 a_112_47.t6 26.595
R302 a_112_47.n15 a_112_47.t2 24.923
R303 a_112_47.n15 a_112_47.t1 24.923
R304 a_112_47.n10 a_112_47.t10 24.923
R305 a_112_47.n10 a_112_47.t8 24.923
R306 a_112_47.n11 a_112_47.t11 24.923
R307 a_112_47.n11 a_112_47.t9 24.923
R308 a_112_47.n13 a_112_47.t0 24.923
R309 a_112_47.n13 a_112_47.t3 24.923
R310 a_112_47.n9 a_112_47.n5 21.76
R311 a_112_47.n2 a_112_47.n1 18.987
R312 a_112_47.n4 a_112_47.n3 7.303
R313 a_112_47.n8 a_112_47.n7 4.381
R314 a_806_297.n4 a_806_297.t8 214.727
R315 a_806_297.n2 a_806_297.n0 198.996
R316 a_806_297.t3 a_806_297.n9 173.769
R317 a_806_297.n4 a_806_297.n3 153.805
R318 a_806_297.n6 a_806_297.n5 153.805
R319 a_806_297.n2 a_806_297.n1 152.525
R320 a_806_297.n8 a_806_297.n7 102.422
R321 a_806_297.n9 a_806_297.n2 65.255
R322 a_806_297.n9 a_806_297.n8 46.108
R323 a_806_297.n6 a_806_297.n4 34.327
R324 a_806_297.n8 a_806_297.n6 34.327
R325 a_806_297.n3 a_806_297.t9 26.595
R326 a_806_297.n3 a_806_297.t10 26.595
R327 a_806_297.n5 a_806_297.t0 26.595
R328 a_806_297.n5 a_806_297.t11 26.595
R329 a_806_297.n7 a_806_297.t2 26.595
R330 a_806_297.n7 a_806_297.t1 26.595
R331 a_806_297.n0 a_806_297.t4 26.595
R332 a_806_297.n0 a_806_297.t7 26.595
R333 a_806_297.n1 a_806_297.t6 26.595
R334 a_806_297.n1 a_806_297.t5 26.595
C0 VPB A 0.12fF
C1 VPWR VGND 0.11fF
C2 VPB B 0.11fF
C3 X VGND 0.76fF
C4 B X 0.27fF
C5 VPB VPWR 0.19fF
C6 A B 0.89fF
C7 VPWR X 0.12fF
C8 B VGND 0.10fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__xor3_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__xor3_1 X C B A VGND VPWR VNB VPB
X0 a_112_21.t2 C.t0 a_404_49.t5 VNB.t9 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1 a_1198_49.t0 a_931_365.t6 VGND.t0 VNB.t7 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X2 a_386_325.t0 B.t0 a_1198_49.t3 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X3 a_404_49.t1 a_266_93.t2 a_112_21.t0 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X4 a_931_365.t0 a_827_297.t2 a_404_49.t0 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X5 VPWR.t4 a_112_21.t4 X.t1 VPB.t10 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 a_827_297.t0 B.t1 VGND.t2 VNB.t5 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 a_1198_49.t4 a_827_297.t3 a_404_49.t4 VNB.t6 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 VGND.t1 A.t0 a_931_365.t2 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X9 a_112_21.t3 C.t1 a_386_325.t5 VPB.t9 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X10 a_1198_49.t5 a_827_297.t4 a_386_325.t4 VPB.t7 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X11 a_266_93.t1 C.t2 VPWR.t3 VPB.t8 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X12 a_1198_49.t1 a_931_365.t7 VPWR.t0 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13 a_931_365.t1 a_827_297.t5 a_386_325.t2 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=600000u l=150000u
X14 VPWR.t2 A.t1 a_931_365.t3 VPB.t6 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 a_827_297.t1 B.t2 VPWR.t1 VPB.t5 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16 VGND.t4 a_112_21.t5 X.t0 VNB.t10 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X17 a_386_325.t1 B.t3 a_931_365.t4 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X18 a_266_93.t0 C.t3 VGND.t3 VNB.t8 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19 a_404_49.t2 B.t4 a_931_365.t5 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X20 a_386_325.t3 a_266_93.t3 a_112_21.t1 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X21 a_404_49.t3 B.t5 a_1198_49.t2 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
R0 C.n0 C.t1 229.135
R1 C.n1 C.t2 154.239
R2 C.n0 C.t0 140.989
R3 C.n2 C.n1 122.135
R4 C.n1 C.t3 102.826
R5 C C.n2 31.584
R6 C.n2 C.n0 25.593
R7 a_404_49.n3 a_404_49.n2 491.4
R8 a_404_49.n1 a_404_49.t1 431.354
R9 a_404_49.n1 a_404_49.t5 407.557
R10 a_404_49.n2 a_404_49.n0 218.359
R11 a_404_49.n2 a_404_49.n1 115.951
R12 a_404_49.n0 a_404_49.t4 99.375
R13 a_404_49.n3 a_404_49.t3 67.718
R14 a_404_49.t0 a_404_49.n3 34.368
R15 a_404_49.n0 a_404_49.t2 25.312
R16 a_112_21.n3 a_112_21.n2 487.904
R17 a_112_21.n2 a_112_21.n1 259.839
R18 a_112_21.n0 a_112_21.t4 231.476
R19 a_112_21.n0 a_112_21.t5 159.176
R20 a_112_21.n2 a_112_21.n0 76
R21 a_112_21.n1 a_112_21.t1 49.687
R22 a_112_21.t0 a_112_21.n3 46.904
R23 a_112_21.n3 a_112_21.t3 42.214
R24 a_112_21.n1 a_112_21.t2 25.312
R25 VNB VNB.t10 6916.79
R26 VNB.t2 VNB.t5 6377.31
R27 VNB.t8 VNB.t9 5426.67
R28 VNB.t5 VNB.t3 4522.22
R29 VNB.t6 VNB.t4 3886.67
R30 VNB.t3 VNB.t6 3715.55
R31 VNB.t10 VNB.t8 2949.72
R32 VNB.t4 VNB.t0 2836.76
R33 VNB.t9 VNB.t2 2688.89
R34 VNB.t0 VNB.t1 2444.44
R35 VNB.t1 VNB.t7 2053.33
R36 a_931_365.n5 a_931_365.t4 483.934
R37 a_931_365.n9 a_931_365.n8 349.224
R38 a_931_365.n1 a_931_365.t7 241.534
R39 a_931_365.n1 a_931_365.t6 170.841
R40 a_931_365.n8 a_931_365.n1 76
R41 a_931_365.n8 a_931_365.n7 55.794
R42 a_931_365.n5 a_931_365.t5 51.982
R43 a_931_365.n0 a_931_365.t0 50.422
R44 a_931_365.n4 a_931_365.t1 42
R45 a_931_365.n10 a_931_365.n9 38.696
R46 a_931_365.n0 a_931_365.t3 28.87
R47 a_931_365.n9 a_931_365.n0 17.589
R48 a_931_365.n3 a_931_365.n2 13.805
R49 a_931_365.n6 a_931_365.n4 9.3
R50 a_931_365.n2 a_931_365.t2 9.275
R51 a_931_365.n6 a_931_365.n5 7.581
R52 a_931_365.n7 a_931_365.n6 3.71
R53 a_931_365.n4 a_931_365.n3 1
R54 VGND.n1 VGND.n0 122.581
R55 VGND.n18 VGND.n17 121.366
R56 VGND.n2 VGND.t2 107.354
R57 VGND.n17 VGND.t3 78.571
R58 VGND.n17 VGND.t4 36
R59 VGND.n0 VGND.t0 25.312
R60 VGND.n0 VGND.t1 25.312
R61 VGND.n19 VGND.n18 9.417
R62 VGND.n3 VGND.n2 7.905
R63 VGND.n4 VGND.n3 4.65
R64 VGND.n6 VGND.n5 4.65
R65 VGND.n8 VGND.n7 4.65
R66 VGND.n10 VGND.n9 4.65
R67 VGND.n12 VGND.n11 4.65
R68 VGND.n14 VGND.n13 4.65
R69 VGND.n16 VGND.n15 4.65
R70 VGND.n4 VGND.n1 0.134
R71 VGND.n19 VGND.n16 0.132
R72 VGND VGND.n19 0.129
R73 VGND.n6 VGND.n4 0.119
R74 VGND.n8 VGND.n6 0.119
R75 VGND.n10 VGND.n8 0.119
R76 VGND.n12 VGND.n10 0.119
R77 VGND.n14 VGND.n12 0.119
R78 VGND.n16 VGND.n14 0.119
R79 a_1198_49.n2 a_1198_49.n0 297.655
R80 a_1198_49.n3 a_1198_49.t0 226.304
R81 a_1198_49.n0 a_1198_49.t5 209.825
R82 a_1198_49.n2 a_1198_49.n1 192.264
R83 a_1198_49.t1 a_1198_49.n3 176.793
R84 a_1198_49.n3 a_1198_49.n2 130.955
R85 a_1198_49.n1 a_1198_49.t4 94.776
R86 a_1198_49.n0 a_1198_49.t2 41.555
R87 a_1198_49.n1 a_1198_49.t3 38.437
R88 B.t5 B.t3 865.992
R89 B.n1 B.n0 298.84
R90 B.n0 B.t2 294.019
R91 B.n2 B.t5 235.107
R92 B.t3 B.n1 215.293
R93 B.n0 B.t1 168.699
R94 B.n2 B.t0 167.627
R95 B.n1 B.t4 167.092
R96 B B.n2 118.163
R97 a_386_325.n1 a_386_325.t5 428.268
R98 a_386_325.n2 a_386_325.n0 250.115
R99 a_386_325.n1 a_386_325.t3 210.453
R100 a_386_325.n3 a_386_325.n2 151.6
R101 a_386_325.n3 a_386_325.t4 83.109
R102 a_386_325.n0 a_386_325.t2 51.386
R103 a_386_325.n4 a_386_325.t1 40.764
R104 a_386_325.n5 a_386_325.n4 39.4
R105 a_386_325.n4 a_386_325.n3 27.703
R106 a_386_325.n0 a_386_325.t0 25.321
R107 a_386_325.n2 a_386_325.n1 11.25
R108 a_266_93.t1 a_266_93.n1 433.201
R109 a_266_93.n0 a_266_93.t2 260.815
R110 a_266_93.n1 a_266_93.t0 229.423
R111 a_266_93.n1 a_266_93.n0 185.702
R112 a_266_93.n0 a_266_93.t3 167.627
R113 VPB.t0 VPB.t5 713.239
R114 VPB.t5 VPB.t4 648.13
R115 VPB.t8 VPB.t9 633.333
R116 VPB.t7 VPB.t3 517.912
R117 VPB.t4 VPB.t7 449.844
R118 VPB.t10 VPB.t8 355.14
R119 VPB.t9 VPB.t0 313.707
R120 VPB.t3 VPB.t2 304.828
R121 VPB VPB.t10 301.869
R122 VPB.t2 VPB.t6 298.909
R123 VPB.t6 VPB.t1 248.598
R124 a_827_297.t1 a_827_297.n3 510.56
R125 a_827_297.n0 a_827_297.t2 283.255
R126 a_827_297.n1 a_827_297.t3 173.52
R127 a_827_297.n0 a_827_297.t5 161.201
R128 a_827_297.n1 a_827_297.t4 154.239
R129 a_827_297.n2 a_827_297.n1 143.911
R130 a_827_297.n4 a_827_297.t1 102.44
R131 a_827_297.n2 a_827_297.n0 94.522
R132 a_827_297.n3 a_827_297.t0 31.795
R133 a_827_297.n3 a_827_297.n2 2.696
R134 X X.n0 152.56
R135 X.n1 X.t0 151.988
R136 X.n0 X.t1 26.595
R137 X X.n1 4.022
R138 VPWR.n0 VPWR.t1 561.841
R139 VPWR.n14 VPWR.n13 327.699
R140 VPWR.n2 VPWR.n1 310.72
R141 VPWR.n13 VPWR.t3 81.57
R142 VPWR.n13 VPWR.t4 36.445
R143 VPWR.n1 VPWR.t0 26.595
R144 VPWR.n1 VPWR.t2 26.595
R145 VPWR.n16 VPWR.n15 4.65
R146 VPWR.n4 VPWR.n3 4.65
R147 VPWR.n6 VPWR.n5 4.65
R148 VPWR.n8 VPWR.n7 4.65
R149 VPWR.n10 VPWR.n9 4.65
R150 VPWR.n12 VPWR.n11 4.65
R151 VPWR.n2 VPWR.n0 4.027
R152 VPWR.n15 VPWR.n14 2.635
R153 VPWR.n4 VPWR.n2 0.137
R154 VPWR.n17 VPWR.n16 0.132
R155 VPWR VPWR.n17 0.129
R156 VPWR.n6 VPWR.n4 0.119
R157 VPWR.n8 VPWR.n6 0.119
R158 VPWR.n10 VPWR.n8 0.119
R159 VPWR.n12 VPWR.n10 0.119
R160 VPWR.n16 VPWR.n12 0.119
R161 A.n0 A.t1 239.503
R162 A.n0 A.t0 168.81
R163 A A.n0 87.52
C0 VPWR VGND 0.10fF
C1 VPB VPWR 0.17fF
C2 X VPWR 0.13fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__xor3_2.ext - technology: sky130A

.subckt sky130_fd_sc_hd__xor3_2 X C B A VGND VPWR VNB VPB
X0 a_120_21.t2 C.t0 a_496_49.t5 VNB.t11 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1 a_1023_365.t0 a_919_297.t2 a_478_325.t0 VNB.t6 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=600000u l=150000u
X2 VGND.t4 a_120_21.t4 X.t3 VNB.t9 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 a_358_93.t0 C.t1 VGND.t5 VNB.t10 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 a_496_49.t1 B.t0 a_1023_365.t5 VNB.t5 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X5 a_496_49.t2 B.t1 a_1290_49.t5 VPB.t5 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X6 a_1290_49.t1 a_919_297.t3 a_496_49.t3 VNB.t7 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7 a_496_49.t0 a_358_93.t2 a_120_21.t0 VPB.t7 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X8 a_1023_365.t1 a_919_297.t4 a_496_49.t4 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X9 a_1290_49.t2 a_1023_365.t6 VGND.t0 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X10 VPWR.t4 a_120_21.t5 X.t1 VPB.t9 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 a_478_325.t4 B.t2 a_1290_49.t4 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X12 X.t0 a_120_21.t6 VPWR.t3 VPB.t8 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13 a_1290_49.t0 a_919_297.t5 a_478_325.t1 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X14 a_919_297.t0 B.t3 VGND.t2 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X15 a_120_21.t3 C.t2 a_478_325.t5 VPB.t11 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X16 a_358_93.t1 C.t3 VPWR.t5 VPB.t10 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X17 a_1290_49.t3 a_1023_365.t7 VPWR.t0 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X18 VGND.t1 A.t0 a_1023_365.t3 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X19 X.t2 a_120_21.t7 VGND.t3 VNB.t8 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X20 VPWR.t2 A.t1 a_1023_365.t4 VPB.t6 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X21 a_919_297.t1 B.t4 VPWR.t1 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X22 a_478_325.t3 B.t5 a_1023_365.t2 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X23 a_478_325.t2 a_358_93.t3 a_120_21.t1 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
R0 C.n0 C.t2 229.135
R1 C.n1 C.t3 154.239
R2 C.n0 C.t0 140.989
R3 C.n2 C.n1 122.135
R4 C.n1 C.t1 102.826
R5 C C.n2 31.584
R6 C.n2 C.n0 25.593
R7 a_496_49.n2 a_496_49.n1 491.4
R8 a_496_49.t0 a_496_49.n3 431.354
R9 a_496_49.n3 a_496_49.t5 407.557
R10 a_496_49.n2 a_496_49.n0 218.359
R11 a_496_49.n3 a_496_49.n2 115.951
R12 a_496_49.n0 a_496_49.t3 99.375
R13 a_496_49.n1 a_496_49.t2 67.718
R14 a_496_49.n1 a_496_49.t4 34.368
R15 a_496_49.n0 a_496_49.t1 25.312
R16 a_120_21.n5 a_120_21.n4 487.904
R17 a_120_21.n4 a_120_21.n3 259.839
R18 a_120_21.n2 a_120_21.t5 212.079
R19 a_120_21.n0 a_120_21.t6 212.079
R20 a_120_21.n0 a_120_21.t7 142.7
R21 a_120_21.n1 a_120_21.t4 139.779
R22 a_120_21.n4 a_120_21.n2 102.29
R23 a_120_21.n1 a_120_21.n0 58.424
R24 a_120_21.n3 a_120_21.t1 49.687
R25 a_120_21.t0 a_120_21.n5 46.904
R26 a_120_21.n5 a_120_21.t3 42.214
R27 a_120_21.n3 a_120_21.t2 25.312
R28 a_120_21.n2 a_120_21.n1 2.921
R29 VNB VNB.t8 7244.69
R30 VNB.t0 VNB.t4 6377.31
R31 VNB.t10 VNB.t11 5426.67
R32 VNB.t4 VNB.t5 4522.22
R33 VNB.t7 VNB.t3 3886.67
R34 VNB.t5 VNB.t7 3715.55
R35 VNB.t9 VNB.t10 2949.72
R36 VNB.t3 VNB.t6 2836.76
R37 VNB.t11 VNB.t0 2688.89
R38 VNB.t6 VNB.t2 2444.44
R39 VNB.t2 VNB.t1 2053.33
R40 VNB.t8 VNB.t9 2030.77
R41 a_919_297.t1 a_919_297.n3 510.56
R42 a_919_297.n0 a_919_297.t4 283.255
R43 a_919_297.n1 a_919_297.t3 173.52
R44 a_919_297.n0 a_919_297.t2 161.201
R45 a_919_297.n1 a_919_297.t5 154.239
R46 a_919_297.n2 a_919_297.n1 143.911
R47 a_919_297.n4 a_919_297.t1 102.44
R48 a_919_297.n2 a_919_297.n0 94.522
R49 a_919_297.n3 a_919_297.t0 31.795
R50 a_919_297.n3 a_919_297.n2 2.696
R51 a_478_325.n1 a_478_325.t5 428.268
R52 a_478_325.n2 a_478_325.n0 250.115
R53 a_478_325.n1 a_478_325.t2 210.453
R54 a_478_325.n3 a_478_325.n2 151.6
R55 a_478_325.n3 a_478_325.t1 83.109
R56 a_478_325.n0 a_478_325.t0 51.386
R57 a_478_325.n4 a_478_325.t3 40.764
R58 a_478_325.n5 a_478_325.n4 39.4
R59 a_478_325.n4 a_478_325.n3 27.703
R60 a_478_325.n0 a_478_325.t4 25.321
R61 a_478_325.n2 a_478_325.n1 11.25
R62 a_1023_365.n5 a_1023_365.t2 483.934
R63 a_1023_365.n9 a_1023_365.n8 349.224
R64 a_1023_365.n1 a_1023_365.t7 241.534
R65 a_1023_365.n1 a_1023_365.t6 170.841
R66 a_1023_365.n8 a_1023_365.n1 76
R67 a_1023_365.n8 a_1023_365.n7 55.794
R68 a_1023_365.n5 a_1023_365.t5 51.982
R69 a_1023_365.n0 a_1023_365.t1 50.422
R70 a_1023_365.n4 a_1023_365.t0 42
R71 a_1023_365.n10 a_1023_365.n9 38.696
R72 a_1023_365.n0 a_1023_365.t4 28.87
R73 a_1023_365.n9 a_1023_365.n0 17.589
R74 a_1023_365.n3 a_1023_365.n2 13.805
R75 a_1023_365.n6 a_1023_365.n4 9.3
R76 a_1023_365.n2 a_1023_365.t3 9.275
R77 a_1023_365.n6 a_1023_365.n5 7.581
R78 a_1023_365.n7 a_1023_365.n6 3.71
R79 a_1023_365.n4 a_1023_365.n3 1
R80 X.n2 X.n0 132.261
R81 X.n2 X.n1 100.072
R82 X.n1 X.t1 26.595
R83 X.n1 X.t0 26.595
R84 X.n0 X.t3 24.923
R85 X.n0 X.t2 24.923
R86 X X.n2 1.377
R87 VGND.n21 VGND.t3 190.315
R88 VGND.n1 VGND.n0 122.581
R89 VGND.n18 VGND.n17 121.366
R90 VGND.n2 VGND.t2 107.355
R91 VGND.n17 VGND.t5 78.571
R92 VGND.n17 VGND.t4 36
R93 VGND.n0 VGND.t0 25.312
R94 VGND.n0 VGND.t1 25.312
R95 VGND.n3 VGND.n2 7.905
R96 VGND.n19 VGND.n18 5.27
R97 VGND.n4 VGND.n3 4.65
R98 VGND.n6 VGND.n5 4.65
R99 VGND.n8 VGND.n7 4.65
R100 VGND.n10 VGND.n9 4.65
R101 VGND.n12 VGND.n11 4.65
R102 VGND.n14 VGND.n13 4.65
R103 VGND.n16 VGND.n15 4.65
R104 VGND.n20 VGND.n19 4.65
R105 VGND.n23 VGND.n22 4.65
R106 VGND.n22 VGND.n21 4.517
R107 VGND.n4 VGND.n1 0.134
R108 VGND.n6 VGND.n4 0.119
R109 VGND.n8 VGND.n6 0.119
R110 VGND.n10 VGND.n8 0.119
R111 VGND.n12 VGND.n10 0.119
R112 VGND.n14 VGND.n12 0.119
R113 VGND.n16 VGND.n14 0.119
R114 VGND.n20 VGND.n16 0.119
R115 VGND.n23 VGND.n20 0.119
R116 VGND.n24 VGND.n23 0.119
R117 VGND VGND.n24 0.022
R118 a_358_93.t1 a_358_93.n1 433.201
R119 a_358_93.n0 a_358_93.t2 260.815
R120 a_358_93.n1 a_358_93.t0 229.423
R121 a_358_93.n1 a_358_93.n0 185.702
R122 a_358_93.n0 a_358_93.t3 167.627
R123 B.t1 B.t5 865.992
R124 B.n1 B.n0 298.84
R125 B.n0 B.t4 294.019
R126 B.n2 B.t1 235.107
R127 B.t5 B.n1 215.293
R128 B.n0 B.t3 168.699
R129 B.n2 B.t2 167.627
R130 B.n1 B.t0 167.092
R131 B B.n2 118.163
R132 a_1290_49.n2 a_1290_49.n0 297.655
R133 a_1290_49.n3 a_1290_49.t2 226.304
R134 a_1290_49.n0 a_1290_49.t0 209.825
R135 a_1290_49.n2 a_1290_49.n1 192.264
R136 a_1290_49.t3 a_1290_49.n3 176.793
R137 a_1290_49.n3 a_1290_49.n2 130.955
R138 a_1290_49.n1 a_1290_49.t1 94.776
R139 a_1290_49.n0 a_1290_49.t5 41.555
R140 a_1290_49.n1 a_1290_49.t4 38.437
R141 VPB.t7 VPB.t4 713.239
R142 VPB.t4 VPB.t3 648.13
R143 VPB.t10 VPB.t11 633.333
R144 VPB.t0 VPB.t5 517.912
R145 VPB.t3 VPB.t0 449.844
R146 VPB.t9 VPB.t10 355.14
R147 VPB VPB.t8 325.545
R148 VPB.t11 VPB.t7 313.707
R149 VPB.t5 VPB.t1 304.828
R150 VPB.t1 VPB.t6 298.909
R151 VPB.t6 VPB.t2 248.598
R152 VPB.t8 VPB.t9 248.598
R153 VPWR.n0 VPWR.t1 561.841
R154 VPWR.n19 VPWR.t3 546.533
R155 VPWR.n14 VPWR.n13 327.699
R156 VPWR.n2 VPWR.n1 310.72
R157 VPWR.n13 VPWR.t5 81.57
R158 VPWR.n13 VPWR.t4 36.445
R159 VPWR.n1 VPWR.t0 26.595
R160 VPWR.n1 VPWR.t2 26.595
R161 VPWR.n21 VPWR.n20 4.65
R162 VPWR.n4 VPWR.n3 4.65
R163 VPWR.n6 VPWR.n5 4.65
R164 VPWR.n8 VPWR.n7 4.65
R165 VPWR.n10 VPWR.n9 4.65
R166 VPWR.n12 VPWR.n11 4.65
R167 VPWR.n16 VPWR.n15 4.65
R168 VPWR.n18 VPWR.n17 4.65
R169 VPWR.n2 VPWR.n0 4.027
R170 VPWR.n20 VPWR.n19 3.011
R171 VPWR.n15 VPWR.n14 2.635
R172 VPWR.n4 VPWR.n2 0.137
R173 VPWR.n6 VPWR.n4 0.119
R174 VPWR.n8 VPWR.n6 0.119
R175 VPWR.n10 VPWR.n8 0.119
R176 VPWR.n12 VPWR.n10 0.119
R177 VPWR.n16 VPWR.n12 0.119
R178 VPWR.n18 VPWR.n16 0.119
R179 VPWR.n21 VPWR.n18 0.119
R180 VPWR.n22 VPWR.n21 0.119
R181 VPWR VPWR.n22 0.022
R182 A.n0 A.t1 239.503
R183 A.n0 A.t0 168.81
R184 A A.n0 87.52
C0 X VGND 0.11fF
C1 VPWR X 0.17fF
C2 VPWR VGND 0.12fF
C3 VPB VPWR 0.18fF
.ends

* NGSPICE file created from sky130_fd_sc_hd__xor3_4.ext - technology: sky130A

.subckt sky130_fd_sc_hd__xor3_4 X C B A VGND VPWR VNB VPB
X0 a_602_325.t1 B.t0 a_1402_49.t1 VNB.t7 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1 a_1031_297.t0 B.t1 VPWR.t4 VPB.t9 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 a_608_49.t3 B.t2 a_1402_49.t0 VPB.t8 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X3 VGND.t7 A.t0 a_1135_365.t5 VNB.t11 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X4 a_1402_49.t4 a_1031_297.t2 a_608_49.t0 VNB.t12 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 a_480_297.t0 C.t0 VPWR.t6 VPB.t11 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X6 a_608_49.t2 a_480_297.t2 a_79_21.t0 VPB.t6 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X7 a_1135_365.t0 a_1031_297.t3 a_608_49.t1 VPB.t1 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X8 X.t3 a_79_21.t4 VPWR.t0 VPB.t2 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 a_1135_365.t1 a_1031_297.t4 a_602_325.t4 VNB.t13 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=600000u l=150000u
X10 VGND.t1 a_79_21.t5 X.t7 VNB.t0 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 VGND.t2 a_79_21.t6 X.t6 VNB.t1 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 a_1031_297.t1 B.t3 VGND.t5 VNB.t6 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 a_1402_49.t5 a_1031_297.t5 a_602_325.t5 VPB.t0 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X14 a_79_21.t3 C.t1 a_602_325.t3 VPB.t12 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X15 a_480_297.t1 C.t2 VGND.t6 VNB.t8 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16 a_608_49.t4 B.t4 a_1135_365.t2 VNB.t5 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X17 VPWR.t7 A.t1 a_1135_365.t4 VPB.t13 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X18 a_1402_49.t3 a_1135_365.t6 VGND.t0 VNB.t10 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X19 X.t5 a_79_21.t7 VGND.t3 VNB.t2 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X20 a_602_325.t2 B.t5 a_1135_365.t3 VPB.t7 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X21 VPWR.t1 a_79_21.t8 X.t2 VPB.t3 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X22 a_602_325.t0 a_480_297.t3 a_79_21.t1 VNB.t4 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X23 X.t1 a_79_21.t9 VPWR.t2 VPB.t4 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X24 a_79_21.t2 C.t3 a_608_49.t5 VNB.t9 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X25 VPWR.t3 a_79_21.t10 X.t0 VPB.t5 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X26 X.t4 a_79_21.t11 VGND.t4 VNB.t3 sky130_fd_pr__nshort ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X27 a_1402_49.t2 a_1135_365.t7 VPWR.t5 VPB.t10 sky130_fd_pr__phighvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
R0 B.t2 B.t5 865.992
R1 B.n1 B.n0 298.84
R2 B.n0 B.t1 294.019
R3 B.n2 B.t2 235.107
R4 B.t5 B.n1 215.293
R5 B.n0 B.t3 168.699
R6 B.n2 B.t0 167.627
R7 B.n1 B.t4 167.092
R8 B B.n2 118.163
R9 a_1402_49.n2 a_1402_49.n0 297.655
R10 a_1402_49.n3 a_1402_49.t3 227.966
R11 a_1402_49.n0 a_1402_49.t5 209.825
R12 a_1402_49.n2 a_1402_49.n1 192.264
R13 a_1402_49.t2 a_1402_49.n3 176.196
R14 a_1402_49.n3 a_1402_49.n2 132.994
R15 a_1402_49.n1 a_1402_49.t4 94.776
R16 a_1402_49.n0 a_1402_49.t0 41.555
R17 a_1402_49.n1 a_1402_49.t1 38.437
R18 a_602_325.n1 a_602_325.t3 428.268
R19 a_602_325.n2 a_602_325.n0 250.115
R20 a_602_325.n1 a_602_325.t0 210.453
R21 a_602_325.n3 a_602_325.n2 151.6
R22 a_602_325.n3 a_602_325.t5 83.109
R23 a_602_325.n0 a_602_325.t4 51.386
R24 a_602_325.n4 a_602_325.t2 40.764
R25 a_602_325.n5 a_602_325.n4 39.4
R26 a_602_325.n4 a_602_325.n3 27.703
R27 a_602_325.n0 a_602_325.t1 25.321
R28 a_602_325.n2 a_602_325.n1 11.25
R29 VNB.t4 VNB.t6 6379.46
R30 VNB VNB.t3 5642.92
R31 VNB.t8 VNB.t9 4742.22
R32 VNB.t6 VNB.t5 4522.22
R33 VNB.t12 VNB.t7 3886.67
R34 VNB.t5 VNB.t12 3715.55
R35 VNB.t1 VNB.t8 3264
R36 VNB.t7 VNB.t13 2836.76
R37 VNB.t9 VNB.t4 2688.89
R38 VNB.t13 VNB.t11 2444.44
R39 VNB.t11 VNB.t10 2248.89
R40 VNB.t2 VNB.t1 2030.77
R41 VNB.t0 VNB.t2 2030.77
R42 VNB.t3 VNB.t0 2030.77
R43 VPWR.n1 VPWR.t4 561.841
R44 VPWR.n23 VPWR.t0 556.396
R45 VPWR.n14 VPWR.n13 441.386
R46 VPWR.n2 VPWR.n0 310.839
R47 VPWR.n19 VPWR.n18 308.79
R48 VPWR.n13 VPWR.t6 66.179
R49 VPWR.n0 VPWR.t7 34.475
R50 VPWR.n13 VPWR.t1 29.055
R51 VPWR.n18 VPWR.t2 26.595
R52 VPWR.n18 VPWR.t3 26.595
R53 VPWR.n0 VPWR.t5 26.595
R54 VPWR.n23 VPWR.n22 24.847
R55 VPWR VPWR.n23 14.438
R56 VPWR.n4 VPWR.n3 4.65
R57 VPWR.n6 VPWR.n5 4.65
R58 VPWR.n8 VPWR.n7 4.65
R59 VPWR.n10 VPWR.n9 4.65
R60 VPWR.n12 VPWR.n11 4.65
R61 VPWR.n15 VPWR.n14 4.65
R62 VPWR.n17 VPWR.n16 4.65
R63 VPWR.n20 VPWR.n19 4.65
R64 VPWR.n22 VPWR.n21 4.65
R65 VPWR.n2 VPWR.n1 3.86
R66 VPWR.n4 VPWR.n2 0.142
R67 VPWR.n6 VPWR.n4 0.119
R68 VPWR.n8 VPWR.n6 0.119
R69 VPWR.n10 VPWR.n8 0.119
R70 VPWR.n12 VPWR.n10 0.119
R71 VPWR.n15 VPWR.n12 0.119
R72 VPWR.n17 VPWR.n15 0.119
R73 VPWR.n20 VPWR.n17 0.119
R74 VPWR.n21 VPWR.n20 0.119
R75  VPWR.n21 0.118
R76  VPWR 0.001
R77 a_1031_297.t0 a_1031_297.n3 510.56
R78 a_1031_297.n0 a_1031_297.t3 283.255
R79 a_1031_297.n1 a_1031_297.t2 173.52
R80 a_1031_297.n0 a_1031_297.t4 161.201
R81 a_1031_297.n1 a_1031_297.t5 154.239
R82 a_1031_297.n2 a_1031_297.n1 143.911
R83 a_1031_297.n4 a_1031_297.t0 102.44
R84 a_1031_297.n2 a_1031_297.n0 94.522
R85 a_1031_297.n3 a_1031_297.t1 31.795
R86 a_1031_297.n3 a_1031_297.n2 2.696
R87 VPB.t6 VPB.t9 713.239
R88 VPB.t9 VPB.t7 648.13
R89 VPB.t11 VPB.t12 603.738
R90 VPB.t0 VPB.t8 517.912
R91 VPB.t7 VPB.t0 449.844
R92 VPB.t12 VPB.t6 313.707
R93 VPB.t8 VPB.t1 304.828
R94 VPB.t1 VPB.t13 298.909
R95 VPB.t3 VPB.t11 292.99
R96 VPB.t13 VPB.t10 272.274
R97 VPB.t4 VPB.t3 248.598
R98 VPB.t5 VPB.t4 248.598
R99 VPB.t2 VPB.t5 248.598
R100 VPB VPB.t2 198.286
R101 a_608_49.n1 a_608_49.t5 547.683
R102 a_608_49.n3 a_608_49.n2 489.895
R103 a_608_49.n1 a_608_49.t2 431.354
R104 a_608_49.n2 a_608_49.n0 219.072
R105 a_608_49.n2 a_608_49.n1 117.457
R106 a_608_49.n0 a_608_49.t0 99.375
R107 a_608_49.n3 a_608_49.t3 67.718
R108 a_608_49.t1 a_608_49.n3 34.368
R109 a_608_49.n0 a_608_49.t4 25.312
R110 A.n0 A.t1 239.503
R111 A.n0 A.t0 168.81
R112 A A.n0 87.52
R113 a_1135_365.n5 a_1135_365.t3 483.934
R114 a_1135_365.n9 a_1135_365.n8 349.224
R115 a_1135_365.n1 a_1135_365.t7 241.534
R116 a_1135_365.n1 a_1135_365.t6 170.841
R117 a_1135_365.n8 a_1135_365.n1 76
R118 a_1135_365.n8 a_1135_365.n7 55.794
R119 a_1135_365.n5 a_1135_365.t2 51.982
R120 a_1135_365.n0 a_1135_365.t0 50.422
R121 a_1135_365.n4 a_1135_365.t1 42
R122 a_1135_365.n10 a_1135_365.n9 38.696
R123 a_1135_365.n0 a_1135_365.t4 28.87
R124 a_1135_365.n9 a_1135_365.n0 17.589
R125 a_1135_365.n3 a_1135_365.n2 13.805
R126 a_1135_365.n6 a_1135_365.n4 9.3
R127 a_1135_365.n2 a_1135_365.t5 9.275
R128 a_1135_365.n6 a_1135_365.n5 7.581
R129 a_1135_365.n7 a_1135_365.n6 3.71
R130 a_1135_365.n4 a_1135_365.n3 1
R131 VGND.n25 VGND.t4 197.787
R132 VGND.n15 VGND.t2 165.378
R133 VGND.n1 VGND.n0 125.985
R134 VGND.n2 VGND.t5 113.911
R135 VGND.n21 VGND.n20 107.239
R136 VGND.t2 VGND.t6 51.428
R137 VGND.n0 VGND.t7 32.812
R138 VGND.n0 VGND.t0 25.312
R139 VGND.n20 VGND.t3 24.923
R140 VGND.n20 VGND.t1 24.923
R141 VGND.n3 VGND.n2 15.435
R142 VGND.n16 VGND.n15 9.788
R143 VGND.n26 VGND.n25 6.908
R144 VGND.n4 VGND.n3 4.65
R145 VGND.n6 VGND.n5 4.65
R146 VGND.n8 VGND.n7 4.65
R147 VGND.n10 VGND.n9 4.65
R148 VGND.n12 VGND.n11 4.65
R149 VGND.n14 VGND.n13 4.65
R150 VGND.n17 VGND.n16 4.65
R151 VGND.n19 VGND.n18 4.65
R152 VGND.n22 VGND.n21 4.65
R153 VGND.n24 VGND.n23 4.65
R154 VGND.n4 VGND.n1 0.134
R155 VGND.n6 VGND.n4 0.119
R156 VGND.n8 VGND.n6 0.119
R157 VGND.n10 VGND.n8 0.119
R158 VGND.n12 VGND.n10 0.119
R159 VGND.n14 VGND.n12 0.119
R160 VGND.n17 VGND.n14 0.119
R161 VGND.n19 VGND.n17 0.119
R162 VGND.n22 VGND.n19 0.119
R163 VGND.n24 VGND.n22 0.119
R164  VGND.n24 0.118
R165 VGND.n26 VGND 0.002
R166  VGND.n26 0.001
R167 C.n0 C.t1 229.135
R168 C.n1 C.t0 167.384
R169 C.n0 C.t3 140.989
R170 C.n1 C.t2 102.826
R171 C.n2 C.n1 101.686
R172 C C.n2 31.584
R173 C.n2 C.n0 25.593
R174 a_480_297.t0 a_480_297.n1 410.154
R175 a_480_297.n0 a_480_297.t2 260.815
R176 a_480_297.n1 a_480_297.t1 189.423
R177 a_480_297.n1 a_480_297.n0 183.73
R178 a_480_297.n0 a_480_297.t3 167.627
R179 a_79_21.n9 a_79_21.n8 481.084
R180 a_79_21.n8 a_79_21.n7 252.467
R181 a_79_21.n6 a_79_21.t8 212.079
R182 a_79_21.n4 a_79_21.t9 212.079
R183 a_79_21.n2 a_79_21.t10 212.079
R184 a_79_21.n0 a_79_21.t4 212.079
R185 a_79_21.n0 a_79_21.t11 154.55
R186 a_79_21.n1 a_79_21.t5 139.779
R187 a_79_21.n3 a_79_21.t7 139.779
R188 a_79_21.n5 a_79_21.t6 139.779
R189 a_79_21.n8 a_79_21.n6 86.954
R190 a_79_21.n7 a_79_21.t1 49.687
R191 a_79_21.t0 a_79_21.n9 46.904
R192 a_79_21.n5 a_79_21.n4 46.739
R193 a_79_21.n3 a_79_21.n2 46.739
R194 a_79_21.n1 a_79_21.n0 46.739
R195 a_79_21.n9 a_79_21.t3 42.214
R196 a_79_21.n7 a_79_21.t2 25.312
R197 a_79_21.n6 a_79_21.n5 14.606
R198 a_79_21.n4 a_79_21.n3 14.606
R199 a_79_21.n2 a_79_21.n1 14.606
R200 X.n2 X.n0 120.557
R201 X.n2 X.n1 112.997
R202 X.n4 X.n3 108.047
R203 X X.n5 107.689
R204 X.n5 X.t0 26.595
R205 X.n5 X.t3 26.595
R206 X.n3 X.t2 26.595
R207 X.n3 X.t1 26.595
R208 X.n4 X.n2 26.412
R209 X.n1 X.t6 24.923
R210 X.n1 X.t5 24.923
R211 X.n0 X.t7 24.923
R212 X.n0 X.t4 24.923
R213 X X.n4 2.009
C0 VPWR VGND 0.15fF
C1 VPB VPWR 0.20fF
C2 X VGND 0.20fF
C3 VPWR X 0.32fF
.ends

